C0018935|HCT
C0018935|red blood cell count
C0018935|Hematocrit
C0018935|Hematocrit procedure
C0518014|Hematocrit
C1542366|Hematocrit
C1545323|Hematocrit test status
C1627395|Hematocrit test results
C1627395|Hematocrit test status &or results
C1627395|Hematocrit test status or results
C1254918|Operating Room Misc Labs: Hct
C0018935|Hct
C0018935|Erythrocyte Volumes, Packed
C0018935|Hematocrit
C0018935|Hematocrits
C0018935|Packed Erythrocyte Volume
C0018935|Packed Erythrocyte Volumes
C0018935|Packed Red Cell Volume
C0018935|Packed Red-Cell Volumes
C0018935|Red-Cell Volume, Packed
C0018935|Red-Cell Volumes, Packed
C0018935|Volume, Packed Erythrocyte
C0018935|Volume, Packed Red-Cell
C0018935|Volumes, Packed Erythrocyte
C0018935|Volumes, Packed Red-Cell
C0018935|Haematocrit
C0018935|Hematocrit procedure
C0018935|hematocrit (lab test)
C0018935|Hematocrit Measurement
C0018935|BLOOD COUNT HEMATOCRIT
C0018935|Measurement of hematocrit (Hct)
C0018935|Packed cell volume (observable entity)
C0018935|Haematocrit - PCV - NOS
C0018935|Packed cell volume
C0018935|Haematocrit (observable entity)
C0018935|Haematocrit (procedure)
C0018935|Hematocrit - PCV - NOS
C0018935|Haematocrit - PCV - NOS (procedure)
C0018935|Hematocrit - PCV - NOS (procedure)
C0018935|hematocrit packed cell volume (lab test)
C0018935|hematocrit packed cell volume
C0018935|EVF
C0018935|PCV
C0018935|Erythrocyte Volume Fraction
C0018935|Blood count; hematocrit (Hct)
C0018935|Packed Red-Cell Volume
C0018935|Erythrocyte Volume, Packed
C0018935|Whole Blood Hematocrit Test
C0018935|Hematocrit determination
C0018935|Haematocrit - PCV
C0018935|Hct - Haematocrit
C0018935|Hct - Hematocrit
C0018935|Hematocrit - PCV
C0018935|Haematocrit determination
C0018935|Hematocrit determination (procedure)
C0018935|Packed cell volume measurement (procedure)
C0018935|Packed cell volume measurement
C0373755|Blood count; spun microhematocrit
C0373755|microhematocrit (spun) (lab test)
C0373755|microhematocrit (spun)
C0373755|microhematocrit level
C0373755|BLOOD COUNT SPUN MICROHEMATOCRIT
C0373755|Measurement of spun microhematocrit
C0373755|SPUN MICROHEMATOCRIT
C0518014|Hematocrit
C0518014|Hematocrit level
C0518014|Hematocrit (Hct)
C0518014|Finding of haematocrit
C0518014|Finding of hematocrit
C0518014|hematocrit finding
C0518014|hematocrit finding (lab test)
C0518014|Haematocrit
C0518014|Finding of hematocrit (finding)
C0518014|Haematocrit - finding
C0518014|Hematocrit - finding
C1988891|Hematocrit &#x7C; blood capillary
C1988890|Hematocrit &#x7C; blood arterial
C3478322|Hematocrit &#x7C; Synovial fluid
C1988896|Hematocrit &#124; Dialysis fluid
C1988896|Hematocrit &#x7C; Dialysis fluid
C1988892|Hematocrit &#x7C; blood cord
C1988893|Hematocrit &#x7C; blood mixed venous
C1988899|Hematocrit &#x7C; urine
C1988895|Hematocrit &#x7C; cerebral spinal fluid
C2968636|Hematocrit &#x7C; Stem cell product
C1988897|Hematocrit &#x7C; body fluid
C1988889|Hematocrit &#x7C; bld-ser-plas
C2738043|Hematocrit &#x7C; Bone marrow
C1988894|Hematocrit &#x7C; blood venous
C3478321|Hematocrit &#x7C; Pleural fluid
C2965246|Hematocrit &#x7C; Fetus &#x7C; Bld-Ser-Plas
C3837271|hematocrit packed cell volume finding
C3837271|hematocrit packed cell volume finding (lab test)
C4028949|hematocrit level by automated count
C4028949|hematocrit level by automated count (lab test)
C4028949|hematocrit by automated count
C4064964|hematocrit level by impedance (lab test)
C4064964|hematocrit by impedance
C4064964|hematocrit level by impedance
C0523148|Haematocrit, spun microhaematocrit method
C0523148|Hematocrit, spun microhematocrit method
C0523148|Hematocrit, spun microhematocrit method (procedure)
C1443988|Serial haematocrit determinations
C1443988|Serial hematocrit determinations (procedure)
C1443988|Serial hematocrit determinations
C0580315|Haematocrit - PCV abnormal (finding)
C0580315|Hematocrit - PCV abnormal
C0580315|Haematocrit - PCV abnormal
C0580315|Hematocrit - packed cell volume abnormal (finding)
C0580315|Hematocrit - PCV abnormal (finding)
C0580315|Hematocrit - packed cell volume abnormal
C0580315|Haematocrit - packed cell volume abnormal
C0474548|Haematocrit - PCV - normal
C0474548|Haematocrit - PCV - normal (finding)
C0474548|Hematocrit - PCV - normal
C0474548|Hematocrit - packed cell volume - normal
C0474548|Hematocrit - packed cell volume - normal (finding)
C0474548|Hematocrit - PCV - normal (finding)
C0474548|Haematocrit - packed cell volume - normal
C0474550|Haematocrit - PCV - low (finding)
C0474550|Haematocrit - PCV - low
C0474550|Hematocrit - PCV - low
C0474550|Packed cell volume decreased below normal
C0474550|Hematocrit decreased below normal
C0474550|HCT decreased
C0474550|PCV decreased below normal
C0474550|Hematocrit - packed cell volume - low
C0474550|Hematocrit - PCV - low (finding)
C0474550|Hematocrit - packed cell volume - low (finding)
C0474550|Haematocrit - packed cell volume - low
C0549409|Haematocrit - PCV - high (finding)
C0549409|Haematocrit - PCV - high
C0549409|Hematocrit - PCV - high
C0549409|PCV increased
C0549409|HCT increased
C0549409|Hematocrit increased above normal
C0549409|Hemoconcentration
C0549409|Packed cell volume increased above normal
C0549409|Hematocrit - PCV - high (finding)
C0549409|Hematocrit - packed cell volume - high (finding)
C0549409|Hematocrit - packed cell volume - high
C0549409|Haematocrit - packed cell volume - high
C0549409|Packed cell volume increased
C0474547|Haematocrit - borderline high
C0474547|Haematocrit - borderline high (finding)
C0474547|Hematocrit - borderline high
C0474547|Hematocrit - borderline high (finding)
C0474551|Haematocrit - borderline low (finding)
C0474551|Haematocrit - borderline low
C0474551|Hematocrit - borderline low
C0474551|Hematocrit - borderline low (finding)
C2004297|Finding of hematocrit - packed cell volume level
C2004297|Finding of haematocrit - packed cell volume level
C2004297|Hematocrit - PCV
C2004297|Hematocrit - P.C.V
C2004297|Haematocrit - PCV
C2004297|Haematocrit - P.C.V
C2004297|Haematocrit - PCV level
C2004297|Hematocrit - PCV level
C2004297|Finding of hematocrit - packed cell volume level (finding)
C2004297|Haematocrit - PCV level - finding
C2004297|Hematocrit - PCV level - finding
C1443990|Stable haematocrit
C1443990|Stable hematocrit (finding)
C1443990|Stable hematocrit
C0878707|precipitous drop in hematocrit
C0878707|precipitous drop in hematocrit (diagnosis)
C0878707|Drop, hematocrit, precip
C0878707|Precipitous drop in haematocrit
C0878707|Precipitous drop in hematocrit (finding)
