C0019682|HIV
C0019693|HIV Infections
C0019704|HIV-1
C0019704|human immunodeficiency virus 1
C0019704|AIDS virus
C0019704|HUMAN IMMUNODEFIC VIRUS 1
C0019704|HUMAN IMMUNODEFICIENCY VIRUS 001
C0019704|HUMAN IMMUNODEFIC VIRUS TYPE 1
C0019704|HIV 01
C0019704|IMMUNODEFIC VIRUS TYPE 1 HUMAN
C0019704|HIV 1
C0019704|human T cell leukemia virus III
C0019704|human T lymphotropic virus III
C0019704|Human immunodeficiency virus type I -RETIRED-
C0019704|human immunodeficiency virus 1 HIV-1
C0019704|human immunodeficiency virus HIV-1
C0019704|human immunodeficiency virus type 1 HIV 1
C0019704|human immunodeficiency virus type 1 HIV-1
C0019704|human immunodeficiency virus type 1 HIV1
C0019704|human immunodeficiency virus type 1, HIV-1
C0019704|human immunodeficiency virus type I HIV-1
C0019704|human immunodeficiency virus type-1 HIV-1
C0019704|human immunodeficiency virus-1 HIV-1
C0019704|HTLV-3 - Human T-cell lymphotropic virus type 3
C0019704|Human immunodeficiency virus type I
C0019704|Human immunodeficiency virus type 1
C0019704|Human T-cell lymphotropic virus 3
C0019704|HIV1 - Human immunodeficiency virus type 1
C0019704|Human immunodeficiency virus type I (organism)
C0019704|Human immunodeficiency virus type 1 (organism)
C0019704|LAV-1
C0019704|Human T-cell leukaemia virus III
C0019704|Human T-cell leukemia virus III
C0019704|Immunodeficiency Virus Type 1, Human
C0019704|HIV-I
C0019704|HIV1
C0019704|Human immunodeficiency virus type 1 [Ambiguous]
C0019704|Human Immunodeficiency Virus, Type 1
C0019707|HIV-2
C0019707|human immunodeficiency virus 2
C0019707|IMMUNODEFIC VIRUS TYPE 2 HUMAN
C0019707|LAV AA 02
C0019707|HUMAN IMMUNODEFIC VIRUS 2
C0019707|HUMAN IMMUNODEFIC VIRUS TYPE 2
C0019707|HIV 02
C0019707|HTLV WIV
C0019707|HUMAN LYMPHOTROPIC VIRUS TYPE IV A T
C0019707|HUMAN IMMUNODEFICIENCY VIRUS 002
C0019707|HIV 2
C0019707|Human immunodeficiency virus 2 (HIV-2)
C0019707|Human immunodeficiency virus type 2 -RETIRED-
C0019707|Human immunodeficiency virus-2
C0019707|human immunodeficiency virus type 2 HIV-2
C0019707|human immunodeficiency virus type 2, HIV-2
C0019707|Human immunodeficiency virus type 2
C0019707|Human immunodeficiency virus type 2 (organism)
C0019707|LAV-2
C0019707|HTLV-IV
C0019707|Human T-Lymphotropic Virus Type IV
C0019707|Immunodeficiency Virus Type 2, Human
C0019707|HIV-II
C0019707|Human T Lymphotropic Virus Type IV
C0019707|HIV type 2
C0019707|HIV2 - Human immunodeficiency virus type 2
C0019707|HIV2
C0019707|Human Immunodeficiency Virus, Type 2
C0019682|HIV
C0019682|Lymphadenopathy Associated Virus
C0019682|Lymphadenopathy-Associated Viruses
C0019682|Virus, Lymphadenopathy-Associated
C0019682|Viruses, Lymphadenopathy-Associated
C0019682|human immunodeficiency virus
C0019682|HUMAN IMMUNODEFIC VIRUSES
C0019682|IMMUNODEFIC VIRUSES HUMAN
C0019682|VIRUS HUMAN IMMUNODEFIC
C0019682|HTLV WIII
C0019682|HUMAN LYMPHOTROPIC VIRUS TYPE III A T
C0019682|HUMAN IMMUNODEFIC VIRUS
C0019682|VIRUSES HUMAN IMMUNODEFIC
C0019682|IMMUNODEFIC VIRUS HUMAN
C0019682|HTLV III
C0019682|LAV
C0019682|Human immunodeficiency virus, NOS
C0019682|Human T Cell Leukemia Virus Type III
C0019682|Virus (HIV), Human Immunodeficiency
C0019682|Human Immunodeficiency Virus (HIV)
C0019682|HIV, Human Immunodeficiency Virus
C0019682|Immunodeficiency Viruses, Human
C0019682|Acquired Immune Deficiency Syndrome Virus
C0019682|Human T Cell Lymphotropic Virus Type III
C0019682|Human T-Cell Lymphotropic Virus Type III
C0019682|LAV-HTLV-III
C0019682|Human T-Cell Leukemia Virus Type III
C0019682|Acquired Immunodeficiency Syndrome Virus
C0019682|Human T Lymphotropic Virus Type III
C0019682|Human T-Lymphotropic Virus Type III
C0019682|Immunodeficiency Virus, Human
C0019682|AIDS Virus
C0019682|Human Immunodeficiency Viruses
C0019682|Lymphadenopathy-Associated Virus
C0019682|Virus, Human Immunodeficiency
C0019682|Viruses, Human Immunodeficiency
C0019682|HTLV-III
C0019682|HIV - Human immunodeficiency virus
C0019682|Human immunodeficiency virus (organism)
C0019682|Human T-lymphotropic virus, type III (HTLV-III)
C0019682|Lymphadenopathy-associated virus (LAV)
C0019682|Lymphadenopathy-associated virus, type I (LAV-I)
C0019682|AIDS Viruses
C0019682|Virus, AIDS
C0019682|Viruses, AIDS
C0019682|Virus-HIV
C0497169|HIV/AIDS
C0319089|T-lymphotropic virus
C0319089|T-lymphotropic virus (organism)
C0319089|T-lymphotropic virus, NOS
C1989665|HIV phenotype &#x7C; isolate
C1954120|human immunodeficiency virus genotype:Susceptibility:Point in time:Isolate:Nominal:Genotyping
C1954120|HIV Gentyp Islt
C1954120|HIV genotype:Susc:Pt:Isolate:Nom:Genotyping
C1954120|HIV genotype [Susceptibility]
C0369501|HIV identified
C0369501|human immunodeficiency virus identified
C3534218|HIV 1 integrase gene &#x7C; Isolate
C1440749|HIV reverse transcriptase+protease gene
C1440733|HIV 1+2
C1440733|HIV 1 & 2
C1977331|human immunodeficiency virus genotype:Susceptibility:Point in time:Isolate:Narrative:Genotyping
C1977331|HIV genotype:Susc:Pt:Isolate:Nar:Genotyping
C1977331|HIV genotype [Susceptibility] in Isolate by Genotype method Narrative
C1977331|HIV Gentyp Islt Nar
C3656356|HIV reverse transcriptase+protease+integrase gene
C4038204|HIV proviral DNA &#x7C; Bld-Ser-Plas
C0001175|Acquired Immuno Deficiency Syndrome
C0001175|Acquired Immuno-Deficiency Syndromes
C0001175|Acquired Immunodeficiency Syndrome
C0001175|Acquired Immunodeficiency Syndromes
C0001175|AIDS
C0001175|Immuno-Deficiency Syndrome, Acquired
C0001175|Immuno-Deficiency Syndromes, Acquired
C0001175|Immunodeficiency Syndromes, Acquired
C0001175|Syndrome, Acquired Immuno-Deficiency
C0001175|Syndrome, Acquired Immunodeficiency
C0001175|Syndromes, Acquired Immuno-Deficiency
C0001175|Syndromes, Acquired Immunodeficiency
C0001175|AIDS (disorder)
C0001175|Acquired immune deficiency syndrome (AIDS)
C0001175|IMMUNODEFIC SYNDROME ACQUIRED
C0001175|ACQUIRED IMMUNO DEFIC SYNDROME
C0001175|ACQUIRED IMMUNE DEFIC SYNDROME
C0001175|IMMUNOL DEFIC SYNDROME ACQUIRED
C0001175|ACQUIRED IMMUNODEFIC SYNDROME
C0001175|acquired immunodeficiency syndrome (HIV-1 stage 6)
C0001175|acquired immunodeficiency syndrome (AIDS) (diagnosis)
C0001175|acquired immunodeficiency syndrome (AIDS)
C0001175|Acquired immune deficiency syndr
C0001175|acquired immune deficiency syndrome [AIDS]
C0001175|Acquired Immune Deficiency Syndrome
C0001175|Acquired Immunodeficiency Syndrome [Disease/Finding]
C0001175|Immunodeficiency Syndrome, Acquired
C0001175|Acquired Immuno-Deficiency Syndrome
C0001175|Immunologic Deficiency Syndrome, Acquired
C0001175|Acquired immune deficiency syndrome (disorder)
C0001175|Acquired immune defic. synd.
C0001175|Acquired human immunodeficiency virus infection syndrome NOS
C0001175|Acquired human immunodeficiency virus infection syndrome NOS (disorder)
C0001175|Acquired immune defic. syndr.
C0001175|Acquired immune deficiency syndrome (AIDS) (disorder)
C0001175|Acquired Immunodeficiency Disease
C0001175|AIDS, Acquired Immunodeficiency Syndrome
C0001175|Acquired Immunodeficiency Syndrome, AIDS
C0001175|Acquired immunodeficiency syndrome NOS
C0001175|Acquired immunodeficiency syndrome, unspecified
C0001175|Autoimmune deficiency syndrome
C0001175|AIDS - Acquired immunodeficiency syndrome
C0001175|Immunodeficiency due to human immunodeficiency virus infection
C0001175|acquired; immunodeficiency syndrome
C0001175|AIDS, NOS
C0001175|Acquired immune deficiency syndrome, NOS
C0001175|Acquired immunodeficiency syndrome, NOS
C0001175|Acquired Immune Deficiency
C0001175|Acquired Immun-Deficiency Synd
C0596049|AIDS/HIV neuropathy
C0019693|HIV infection
C0019693|HIV Infections
C0019693|HTLV III Infections
C0019693|HTLV III LAV Infections
C0019693|Infection, HIV
C0019693|Infection, HTLV-III
C0019693|Infection, HTLV-III-LAV
C0019693|Infections, HIV
C0019693|Infections, HTLV-III
C0019693|Infections, HTLV-III-LAV
C0019693|Human immunodeficiency virus [HIV] disease
C0019693|Unspecified human immunodeficiency virus [HIV] disease
C0019693|LYMPHOTROPIC VIRUS TYPE III INFECTIONS HUMAN T
C0019693|HTLV III INFECT
C0019693|HTLV WIII LAV INFECTIONS
C0019693|HTLV WIII INFECTIONS
C0019693|T LYMPHOTROPIC VIRUS TYPE III INFECT HUMAN
C0019693|HIV INFECT
C0019693|HTLV III LAV INFECT
C0019693|HTLV-III/LAV infection, NOS
C0019693|human immunodeficiency virus (HIV) infection
C0019693|human immunodeficiency virus (HIV) infection (diagnosis)
C0019693|HTLV-III/LAV infection -RETIRED-
C0019693|human T-lymphotropic virus 3 (HTLV-III) infection (diagnosis)
C0019693|lymphadenopathy-associated virus (diagnosis)
C0019693|lymphadenopathy-associated virus
C0019693|human T-lymphotropic virus 3 (HTLV-III) infection
C0019693|Human immunodeficiency virus infection, unspecified
C0019693|Human immuno virus dis
C0019693|T-Lymphotropic Virus Type III Infections, Human
C0019693|HIV Infections [Disease/Finding]
C0019693|HTLV-III-LAV Infections
C0019693|HTLV-III Infections
C0019693|Infection;HIV
C0019693|Human immunodeficiency virus [HIV] disease (B20)
C0019693|HTLV-III Infection
C0019693|HTLV-III-LAV Infection
C0019693|T Lymphotropic Virus Type III Infections, Human
C0019693|[X]Human immunodeficiency virus disease (disorder)
C0019693|HTLV-III/LAV infection
C0019693|[X]Unspecified human immunodeficiency virus [HIV] disease
C0019693|Human immunodeficiency virus infection
C0019693|[X]Unspecified human immunodeficiency virus [HIV] disease (disorder)
C0019693|[X]Human immunodeficiency virus disease
C0019693|HTLV-III/LAV infection (disorder)
C0019693|HIV
C0019693|Human immunodeficiency virus syndrome
C0019693|HIV disease
C0019693|HIV infection NOS
C0019693|HIV - Human immunodeficiency virus infection
C0019693|Human immunodeficiency virus infection (disorder)
C0019693|HIV disease; disease (i.e. caused by HIV disease)
C0019693|HIV disease; infection
C0019693|disease (or disorder); HIV disease (resulting from HIV disease)
C0019693|disease (or disorder); resulting from HIV disease
C0019693|human immunodeficiency virus; disease
C0019693|immunodeficiency virus disease; human
C0019693|infection; HIV disease as cause
C0019693|Human immunodeficiency virus infection, NOS
C0019693|Human Immunodeficiency Virus
C0019693|Human immunodeficiency virus disease
C0019693|HUMAN IMMUNODEFICIENCY VIRUS [HIV] INFECTION
C0348209|HIV disease resulting in other infectious and parasitic diseases
C0348209|HIV disease resulting in unspecified infectious or parasitic disease
C0348209|Human immunodeficiency virus [HIV] disease resulting in infectious and parasitic diseases
C0348209|[X]Hiv disease resulting in unspecified infectious and parasitic disease
C0348209|[X]Hiv disease resulting in unspecified infectious and parasitic disease (disorder)
C0348209|[X]Hiv disease resulting in other infectious and parasitic diseases
C0348209|[X]Hiv disease resulting in other infectious and parasitic diseases (disorder)
C0348213|HIV disease resulting in unspecified malignant neoplasm
C0348213|Human immunodeficiency virus [HIV] disease resulting in malignant neoplasms
C0348213|[X]HIV disease resulting in unspecified malignant neoplasm
C0348213|[X]HIV disease resulting in unspecified malignant neoplasm (disorder)
C0348213|HIV disease; neoplasm, malignant
C0494097|Human immunodeficiency virus [HIV] disease resulting in other conditions
C0494096|Human immunodeficiency virus [HIV] disease resulting in other specified diseases
C0152983|Human immunodeficiency virus infection causing other specified conditions
C0152987|Other human immunodeficiency virus infection
C1142553|Primary HIV infection
C0152979|Human immunodeficiency virus infection with specified conditions
C0152988|Human immunodeficiency virus infection causing specified acute infections
C0343752|Acute HIV infection
C0343752|Acute HIV infection syndrome
C0343752|Acute human immunodeficiency virus infection (disorder)
C0343752|Acute HIV infection (disorder)
C0343752|HIV infection acute
C0343752|Acute HIV infection (diagnosis)
C0343752|Acute infection with HIV
C0343752|HIV seroconversion illness
C0343752|Acute human immunodeficiency virus infection
C0343752|Acute human immunodeficiency virus seroconversion illness
C0343751|Asymptomatic HIV infection
C0343751|hiv infection asymptomatic
C0343751|Asymptomatic HIV infection (diagnosis)
C0343751|Asymptomatic infection with HIV
C0343751|Asymptomatic human immunodeficiency virus infection
C0343751|Asymptomatic human immunodeficiency virus infection (disorder)
C0864665|HIV infection, symptomatic
C0864665|symptomatic HIV infection
C0864665|hiv infection symptomatic
C0864665|symptomatic HIV infection (diagnosis)
C0001857|AIDS Related Complex
C0001857|AIDS-Related Complex
C0001857|Complex, AIDS-Related
C0001857|Lymphadenopathy Syndromes
C0001857|Syndrome, Lymphadenopathy
C0001857|Syndromes, Lymphadenopathy
C0001857|AIDS-like syndrome (disorder)
C0001857|AIDS RELAT COMPLEX
C0001857|AIDS-related complex [ARC]
C0001857|Lymphadenopathy Syndrome
C0001857|AIDS-Related Complex [Disease/Finding]
C0001857|ARC
C0001857|Acquired immunodeficiency syndrome (AIDS)-like syndrome (disorder)
C0001857|Acquired immune deficiency syndrome (& [ARC])
C0001857|Acquired immune deficiency syndrome (& [ARC]) (disorder)
C0001857|Aids-related complex (ARC)
C0001857|Acquired immunodeficiency syndrome-like syndrome
C0001857|acquired immunodeficiency syndrome-like syndrome (diagnosis)
C0001857|Acquired immunodeficiency syndrome-related complex, unspecified
C0001857|AIDS-like syndrome
C0001857|Acquired immunodeficiency syndrome (AIDS)-like syndrome
C0001857|Acquired immune deficiency syndrome-related complex (disorder)
C0001857|Acquired immunodeficiency syndrome-like syndrome (disorder)
C0001857|ARC - Acquired immunodeficiency syndrome-related complex
C0001857|Acquired immune deficiency syndrome-related complex
C0019699|AIDS Seroconversions
C0019699|AIDS Seropositivities
C0019699|HIV Seroconversions
C0019699|HIV Seropositivities
C0019699|HIV Seropositivity
C0019699|HTLV III Seroconversion
C0019699|HTLV III Seropositivity
C0019699|HTLV-III Seroconversions
C0019699|HTLV-III Seropositivities
C0019699|Seroconversion, AIDS
C0019699|Seroconversion, HIV
C0019699|Seroconversion, HTLV-III
C0019699|Seroconversions, AIDS
C0019699|Seroconversions, HIV
C0019699|Seroconversions, HTLV-III
C0019699|Seropositivities, AIDS
C0019699|Seropositivities, HIV
C0019699|Seropositivities, HTLV-III
C0019699|Seropositivity, AIDS
C0019699|Seropositivity, HIV
C0019699|Seropositivity, HTLV-III
C0019699|Anti HIV Positivity
C0019699|Anti-HIV Positivities
C0019699|Antibody Positivities, HIV
C0019699|Antibody Positivity, HIV
C0019699|HIV Antibody Positivities
C0019699|Positivities, Anti-HIV
C0019699|Positivities, HIV Antibody
C0019699|Positivity, Anti-HIV
C0019699|Positivity, HIV Antibody
C0019699|HIV positive
C0019699|HIV positive (finding)
C0019699|HIV seropositivity (disorder)
C0019699|Human immunodeficiency virus (HIV) positive
C0019699|HIV ANTIBODY POS
C0019699|HTLV III SEROPOS
C0019699|ANTIHIV POSITIVITY
C0019699|HTLV WIII SEROCONVERSION
C0019699|HIV SEROPOS
C0019699|AIDS SEROPOS
C0019699|HTLV WIII SEROPOSITIVITY
C0019699|ANTI HIV POS
C0019699|seropositive (AIDS test)
C0019699|HIV test positive
C0019699|HIV positve
C0019699|HIV test positve
C0019699|HIV positive NOS
C0019699|AIDS Seroconversion
C0019699|HTLV-III Seroconversion
C0019699|HIV Antibody Positivity
C0019699|HIV Seropositivity [Disease/Finding]
C0019699|Anti-HIV Positivity
C0019699|AIDS Seropositivity
C0019699|HTLV-III Seropositivity
C0019699|HIV Seroconversion
C0019699|antibody positive AIDS test
C0019699|antigen positive AIDS test
C0019699|Human immunodeficiency virus positive (finding)
C0019699|Human immunodeficiency virus (HIV) positive (finding)
C0019699|Human immunodeficiency virus positive
C0019699|Human immunodeficiency virus (HIV) seropositivity (disorder)
C0019699|HIV seropositivity (diagnosis)
C0019699|Human immunodeficiency virus seropositivity (disorder)
C0019699|Human immunodeficiency virus (HIV) seropositivity
C0019699|Human immunodeficiency virus seropositivity
C0019699|Positive test for HIV
C0019699|HTLV III test positive
C0019699|HIV seropositive NOS
C0019699|HTLV-3 antibody positive
C0019699|HIV+
C0019699|HIV-test; positive
C0019699|HIV; positive
C0019699|HIV; test, positive
C0019699|positive; HIV-test
C0019699|positive; HIV
C0019699|test; HIV, positive
C0019699|HIV Positivity
C0001849|AIDS Dementia Complex
C0001849|Complex, AIDS Dementia
C0001849|Dementia, HIV
C0001849|Dementia in human immunodeficiency virus [HIV] disease
C0001849|ADC - Acquired immune deficiency syndrome dementia complex
C0001849|Acquired immune deficiency syndrome dementia complex
C0001849|AIDS - Acquired immune deficiency syndrome dementia complex
C0001849|Acquired immune deficiency syndrome-related dementia
C0001849|Dementia associated with AIDS
C0001849|DEMENTIA COMPLEX AIDS RELAT
C0001849|HIV ASSOC COGNITIVE MOTOR COMPLEX
C0001849|DEMENTIA COMPLEX ACQUIRED IMMUNE DEFIC SYNDROME
C0001849|ACQUIRED IMMUNE DEFIC SYNDROME DEMENTIA COMPLEX
C0001849|AIDS RELAT DEMENTIA COMPLEX
C0001849|acquired immunodeficiency syndrome (AIDS) dementia
C0001849|acquired immunodeficiency syndrome (AIDS) dementia (diagnosis)
C0001849|AIDS dementia
C0001849|Dementia Complex, AIDS
C0001849|AIDS Related Dementia Complex
C0001849|Complex, AIDS-Related Dementia
C0001849|Dementia Complex, AIDS Related
C0001849|Dementias, HIV
C0001849|HIV Dementias
C0001849|Dementia Complex, AIDS-Related
C0001849|Acquired-Immune Deficiency Syndrome Dementia Complex
C0001849|AIDS-Related Dementia Complex
C0001849|Dementia Complex, Acquired Immune Deficiency Syndrome
C0001849|AIDS Dementia Complex [Disease/Finding]
C0001849|HIV Dementia
C0001849|HIV-Associated Cognitive Motor Complex
C0001849|HIV Associated Cognitive Motor Complex
C0001849|HIV associated cognitive and motor complex
C0001849|AIDS with dementia (disorder)
C0001849|Acquired immune deficiency syndrome dementia complex (disorder)
C0001849|AIDS with dementia
C0001849|Dementia associated with AIDS (disorder)
C0001849|Dementia associated with acquired immunodeficiency syndrome
C0001849|Dementia associated with acquired immunodeficiency syndrome (disorder)
C0001849|HIV-related dementia
C0001849|AIDS-dementia complex
C0001849|AIDS-related dementia
C0001849|Dementia due to HIV disease
C0001849|HIV disease; dementia (etiology)
C0001849|HIV disease; dementia (manifestation)
C0001849|HIV disease; resulting in, dementia (etiology)
C0001849|HIV disease; resulting in, dementia (manifestation)
C0001849|dementia; human immunodeficiency virus disease (etiology)
C0001849|dementia; human immunodeficiency virus disease (manifestation)
C0001849|AIDS with dementia, NOS
C0078911|AIDS Associated Nephropathy
C0078911|AIDS Nephropathies
C0078911|AIDS-Associated Nephropathy
C0078911|HIV Associated Nephropathy
C0078911|HIV Related Nephropathy
C0078911|Nephropathies, AIDS
C0078911|Nephropathy, AIDS
C0078911|AIDS Associated Nephropathies
C0078911|HIV Associated Nephropathies
C0078911|HIV Related Nephropathies
C0078911|Nephropathies, AIDS Associated
C0078911|Nephropathies, HIV Associated
C0078911|Nephropathies, HIV Related
C0078911|Nephropathy, AIDS Associated
C0078911|Nephropathy, HIV Associated
C0078911|Nephropathy, HIV Related
C0078911|HIV-Associated Nephropathy
C0078911|AIDS-Related Nephropathy
C0078911|HIV RELAT NEPHROPATHIES
C0078911|HIV RELAT NEPHROPATHY
C0078911|NEPHROPATHY HIV RELAT
C0078911|NEPHROPATHY AIDS ASSOC
C0078911|NEPHROPATHY HIV ASSOC
C0078911|AIDS ASSOC NEPHROPATHIES
C0078911|HIVAN
C0078911|HUMAN IMMUNODEFIC VIRUS ASSOC NEPHROPATHY
C0078911|NEPHROPATHIES AIDS ASSOC
C0078911|NEPHROPATHIES HIV RELAT
C0078911|AIDS ASSOC NEPHROPATHY
C0078911|HIV ASSOC NEPHROPATHIES
C0078911|NEPHROPATHIES HIV ASSOC
C0078911|HIV-associated nephropathy (diagnosis)
C0078911|AIDS-Associated Nephropathies
C0078911|HIV-Related Nephropathies
C0078911|Nephropathies, AIDS-Associated
C0078911|HIV-Associated Nephropathies
C0078911|AIDS Nephropathy
C0078911|Nephropathies, HIV-Associated
C0078911|HIV-Related Nephropathy
C0078911|Nephropathies, HIV-Related
C0078911|Nephropathy, AIDS-Associated
C0078911|Nephropathy, HIV-Associated
C0078911|Nephropathy, HIV-Related
C0078911|AIDS-Associated Nephropathy [Disease/Finding]
C0078911|Human Immunodeficiency Virus-Associated Nephropathy
C0078911|Human Immunodeficiency Virus Associated Nephropathy
C0078911|HIV Nephropathy
C0078911|Human immunodeficiency virus-related nephropathy
C0078911|AIDS - Acquired immune deficiency synd-related nephropathy
C0078911|Acquired immune deficiency syndrome-related nephropathy
C0078911|Acquired immune deficiency syndrome-related nephropathy (disorder)
C0162526|AIDS-Related Opportunistic Infections
C0162526|AIDS Related Opportunistic Infections
C0162526|AIDS-Related Opportunistic Infection
C0162526|Opportunistic Infection, AIDS-Related
C0162526|Opportunistic Infections, AIDS Related
C0162526|HIV Related Opportunistic Infections
C0162526|HIV-Related Opportunistic Infection
C0162526|Infection, HIV-Related Opportunistic
C0162526|Infections, HIV-Related Opportunistic
C0162526|Opportunistic Infection, HIV-Related
C0162526|Opportunistic Infections, HIV Related
C0162526|HIV RELAT OPPORTUNISTIC INFECT
C0162526|OPPORTUNISTIC INFECT AIDS RELAT
C0162526|AIDS RELAT OPPORTUNISTIC INFECT
C0162526|OPPORTUNISTIC INFECT HIV RELAT
C0162526|HIV-Related Opportunistic Infections
C0162526|Opportunistic Infections, HIV-Related
C0162526|AIDS-Related Opportunistic Infections [Disease/Finding]
C0162526|Opportunistic Infections, AIDS-Related
C0162526|Opportunistic Infections in AIDS
C0162526|AIDS Associated Opportunistic Infection
C0162526|AIDS, Opportunistic Infection
C0282616|AIDS Associated Enteropathy
C0282616|AIDS Enteropathies
C0282616|AIDS-Associated Enteropathies
C0282616|Enteropathies, AIDS
C0282616|Enteropathies, AIDS-Associated
C0282616|Enteropathies, HIV
C0282616|Enteropathies, HIV-Associated
C0282616|Enteropathy, AIDS
C0282616|Enteropathy, AIDS Associated
C0282616|Enteropathy, HIV Associated
C0282616|HIV Associated Enteropathy
C0282616|HIV Enteropathies
C0282616|HIV Enteropathy
C0282616|HIV-Associated Enteropathies
C0282616|HIV ASSOC ENTEROPATHY
C0282616|ENTEROPATHY HIV ASSOC
C0282616|ENTEROPATHY AIDS ASSOC
C0282616|AIDS ASSOC ENTEROPATHY
C0282616|infectious diarrhea of HIV patient
C0282616|infectious diarrhea of HIV patient (diagnosis)
C0282616|AIDS Enteropathy
C0282616|AIDS-Associated Enteropathy
C0282616|Enteropathy, HIV
C0282616|Enteropathy, HIV-Associated
C0282616|Idiopathic AIDS Enteropathy
C0282616|Enteropathy, AIDS-Associated
C0282616|HIV Enteropathy [Disease/Finding]
C0282616|HIV-Associated Enteropathy
C0282616|HIV enteropathy (diagnosis)
C0282616|AIDS Enteropathies, Idiopathic
C0282616|AIDS Enteropathy, Idiopathic
C0282616|Enteropathies, Idiopathic AIDS
C0282616|Enteropathy, Idiopathic AIDS
C0282616|Idiopathic AIDS Enteropathies
C0282616|HIV - Human immunodeficiency virus diarrhea
C0282616|HIV - Human immunodeficiency virus diarrhoea
C0282616|HIV - Human immunodeficiency virus enteropathy
C0282616|Human immunodeficiency virus diarrhea
C0282616|Human immunodeficiency virus diarrhoea
C0282616|Human immunodeficiency virus enteropathy
C0282616|Human immunodeficiency virus non-pathogenic diarrhea
C0282616|Human immunodeficiency virus non-pathogenic diarrhoea
C0282616|Human immunodeficiency virus enteropathy (disorder)
C0343755|HIV Wasting Syndrome
C0343755|HIV disease resulting in wasting syndrome
C0343755|Wasting Syndrome, AIDS
C0343755|Human immunodeficiency virus infection wasting syndrome
C0343755|Slim disease
C0343755|HIV - Human immunodeficiency virus infection wasting syndrome
C0343755|Cachexia associated with AIDS
C0343755|HIV WASTING DIS
C0343755|SLIM DIS
C0343755|WASTING DIS HIV
C0343755|AIDS wasting syndrome
C0343755|HIV Wasting Syndrome [Disease/Finding]
C0343755|HIV Wasting Disease
C0343755|Wasting Disease, HIV
C0343755|Wasting Syndrome, HIV
C0343755|Human immunodeficiency virus infection wasting syndrome (disorder)
C0343755|AIDS with cachexia
C0343755|AIDS with cachexia (disorder)
C0343755|Cachexia associated with acquired immunodeficiency syndrome
C0343755|Cachexia associated with acquired immunodeficiency syndrome (finding)
C0343755|Cachexia associated with AIDS (finding)
C0343755|HIV disease; failure to thrive
C0343755|HIV disease; resulting in, failure to thrive
C0343755|HIV disease; resulting in, wasting syndrome
C0343755|disease (or disorder); slim disease (HIV)
C0343755|disease; slim
C0752330|AIDS ARTERITIS CNS
C0752330|CNS AIDS ARTERITIS
C0752330|AIDS Arteritis, Central Nervous System
C0752330|Central Nervous System AIDS Arteritis
C0752330|AIDS Arteritis, Central Nervous System [Disease/Finding]
C1136321|HIV ASSOC LIPODYSTROPHY SYNDROME
C1136321|HIV ASSOC LIPODYSTROPHY
C1136321|HIV Lipodystrophy Syndrome
C1136321|HIV-Associated Lipodystrophy Syndrome
C1136321|HIV-Associated Lipodystrophy
C1136321|HIV-Associated Lipodystrophy Syndrome [Disease/Finding]
C1136321|Lipodystrophy Syndrome, HIV
C1136321|HIV Associated Lipodystrophy
C1136321|HIV Associated Lipodystrophy Syndrome
C1136321|Lipodystrophy Syndrome, HIV-Associated
C1136321|Lipodystrophy, HIV-Associated
C0520783|Congenital HIV infection
C0520783|HIV infection congenital
C0520783|Congenital HIV infection (diagnosis)
C0520783|Congenital human immunodeficiency virus infection
C0520783|Congenital human immunodeficiency virus infection (disorder)
C2319244|HIV infection CDC classification (diagnosis)
C2319244|HIV infection CDC classification
C2046425|HIV infection, stage 0 (diagnosis)
C2046425|HIV infection, stage 0
C2046426|HIV infection, stage 1 (diagnosis)
C2046426|HIV infection, stage 1
C2046427|HIV infection, stage 2 (PGL) (diagnosis)
C2046427|PGL (persistent generalized lymphadenopathy) stage II of HIV infection
C2046427|HIV infection, stage 2 (PGL)
C2240389|HIV infection, stage 3 (PGL) (diagnosis)
C2240389|HIV infection, stage 3 (PGL)
C2240389|PGL (persistent generalized lymphadenopathy) stage III of HIV infection
C2046428|HIV infection, stage 4
C2046428|HIV infection, stage 4 (diagnosis)
C2046429|ARC (AIDS-related complex) stage V of HIV infection
C2046429|HIV infection, stage 5 (ARC)
C2046429|HIV infection, stage 5 (ARC) (diagnosis)
C0276554|AIDS with lymphadenopathy
C0276554|AIDS with lymphadenopathy (disorder)
C0276554|Lymphadenopathy associated with AIDS (disorder)
C0276554|Lymphadenopathy associated with AIDS
C0276554|Lymphadenopathy associated with acquired immunodeficiency syndrome (disorder)
C0276554|Lymphadenopathy associated with acquired immunodeficiency syndrome
C1834751|CORONARY ARTERY DISEASE, DEVELOPMENT OF, IN HIV
C1304455|Oral hairy leukoplakia associated with human immunodeficiency virus disease (disorder)
C1304455|Oral hairy leukoplakia associated with HIV disease (disorder)
C1304455|Oral hairy leukoplakia associated with human immunodeficiency virus disease
C1304455|Oral hairy leucoplakia associated with human immunodeficiency virus disease
C1304455|Oral hairy leucoplakia associated with HIV disease
C1304455|Oral hairy leukoplakia associated with HIV disease
C0276535|AIDS with Kaposi's sarcoma
C0276535|HIV disease resulting in Kaposi's sarcoma
C0276535|Kaposi's sarcoma associated with AIDS
C0276535|AIDS-Related Kaposi Sarcoma
C0276535|AIDS-Related Kaposi's Sarcoma
C0276535|Kaposi's sarcoma AIDS related
C0276535|Kaposi sarcoma associated with AIDS
C0276535|HIV disease resulting in Kaposi's sarcoma (disorder)
C0276535|AIDS with Kaposi's sarcoma (disorder)
C0276535|Kaposi's sarcoma associated with AIDS (disorder)
C0276535|Kaposi's sarcoma associated with acquired immunodeficiency syndrome (disorder)
C0276535|Kaposi's sarcoma associated with acquired immunodeficiency syndrome
C0276535|malignant neoplasm sarcoma kaposi's associated with aids
C0276535|Kaposi's sarcoma associated with AIDS (diagnosis)
C0276535|Kaposi's sarcoma epidemic type
C0276535|Epidemic Kaposi's sarcoma
C0276535|AIDS related Kaposi's sarcoma
C0276535|AIDS related multiple hemorrhagic sarcoma
C0276535|AIDS-associated Kaposi's sarcoma
C0276535|Kaposi's sarcoma, AIDS related
C0276535|Kaposi's sarcoma, epidemic
C0276535|acquired immune deficiency syndrome related Kaposi's sarcoma
C0276535|multiple hemorrhagic sarcoma, AIDS related
C0276535|sarcoma, Kaposi's, AIDS related
C0276535|sarcoma, multiple hemorrhagic, AIDS related
C0276535|HIV disease; Kaposi's sarcoma
C0276535|HIV disease; sarcoma, Kaposi
C0276535|Kaposi; sarcoma, resulting from HIV disease
C0276535|sarcoma; Kaposi, resulting from HIV disease
C0276535|Autoimmune Deficiency Syndrome-Related Kaposi Sarcoma
C0276535|AIDS, Kaposi's Sarcoma
C0348804|HIV disease resulting in Pneumocystis carinii pneumonia
C0348804|HIV disease resulting in Pneumocystis carinii pneumonia (disorder)
C0348804|HIV disease; pneumocystosis
C0348804|HIV disease; resulting in, Pneumocystis carinii pneumonia
C0348804|HIV disease; resulting in, infection, Pneumocystis carinii (pneumonia)
C0348804|Pneumocystis carinii; infection, resulting from HIV disease
C0348804|infection; Pneumocystis carinii, resulting from HIV disease
C0348804|pneumocystosis; pneumonia, resulting from HIV disease
C0348804|pneumocystosis; resulting from HIV disease
C0348804|pneumonia; pneumocystosis, resulting from HIV disease
C0452192|HIV disease resulting in other types of non-Hodgkin's lymphoma
C0452192|HIV disease resulting in other types of non-Hodgkin's lymphoma (disorder)
C0452192|Human immunodeficiency virus (HIV) disease resulting in other types of non-Hodgkin's lymphoma (disorder)
C0452192|Human immunodeficiency virus (HIV) disease resulting in other types of non-Hodgkin's lymphoma
C0348983|Human immunodef virus resulting in other disease (disorder)
C0348983|Human immunodef virus resulting in other disease
C0343749|Human immunodeficiency virus with other clinical findings
C0343749|Human immunodeficiency virus with other clinical findings (disorder)
C0343757|HIV neuropathy
C0343757|Human immunodeficiency virus neuropathy (disorder)
C0343757|HIV - Human immunodeficiency virus neuropathy
C0343757|Human immunodeficiency virus neuropathy
C0343757|Neuropathy due to human immunodeficiency virus
C0343757|neuropathy due to human immunodeficiency virus (diagnosis)
C0343757|Neuropathy due to human immunodeficiency virus (disorder)
C0343757|Neuropathy caused by human immunodeficiency virus (disorder)
C0343757|Neuropathy caused by human immunodeficiency virus
C0343757|Neuropathy caused by HIV - human immunodeficiency virus
C0343757|Neuropathy due to HIV - human immunodeficiency virus
C3648901|HIV infection complicating pregnancy, childbirth, and puerperium
C3648901|HIV infection complicating pregnancy, childbirth, and puerperium (diagnosis)
C3648903|HIV infection complicating childbirth
C3648903|hiv infection complicating childbirth (diagnosis)
C3648900|HIV infection complicating puerperium
C3648900|HIV infection complicating puerperium (diagnosis)
C3661937|Symptomatic human immunodeficiency virus infection (disorder)
C3661937|Symptomatic human immunodeficiency virus infection
C0343748|HIV infection with secondary cancers
C0343748|HIV infection with secondary cancers (diagnosis)
C0343748|Human immunodeficiency virus with secondary cancers
C0343748|Human immunodeficiency virus with secondary cancers (disorder)
C0343754|HIV infection constitutional disease (diagnosis)
C0343754|HIV infection constitutional disease
C0343754|HIV infection with constitutional disease
C0343754|HIV - Human immunodeficiency virus infection constitutional disease
C0343754|Human immunodeficiency virus infection constitutional disease
C0343754|Human immunodeficiency virus infection constitutional disease (disorder)
C1274337|HIV seroconversion exanthem (disorder)
C1274337|Human immunodeficiency virus (HIV) seroconversion exanthem (disorder)
C1274337|HIV seroconversion exanthem
C1274337|HIV seroconversion exanthem (diagnosis)
C1274337|Human immunodeficiency virus seroconversion exanthem
C1274337|Human immunodeficiency virus (HIV) seroconversion exanthem
C1274337|Human immunodeficiency virus seroconversion exanthem (disorder)
C0276600|HIV infection with aseptic meningitis (disorder)
C0276600|Human immunodeficiency virus (HIV) infection with aseptic meningitis
C0276600|Human immunodeficiency virus infection with aseptic meningitis
C0276600|Human immunodeficiency virus infection with aseptic meningitis (disorder)
C0276600|Human immunodeficiency virus (HIV) infection with aseptic meningitis (disorder)
C0276600|AIDS virus with aseptic meningitis (disorder)
C0276600|AIDS virus with aseptic meningitis
C0276600|HIV infection with aseptic meningitis
C0276600|HIV infection with aseptic meningitis (diagnosis)
C0276600|HIV infection with aseptic meningitis (disorder) [Ambiguous]
C0206019|HIV disease resulting in encephalopathy
C0206019|ENCEPH HIV
C0206019|ENCEPH AIDS
C0206019|HIV ENCEPH
C0206019|AIDS ENCEPH
C0206019|HIV encephalopathy
C0206019|acquired immunodeficiency syndrome (AIDS) encephalopathy
C0206019|acquired immunodeficiency syndrome (AIDS) encephalopathy (diagnosis)
C0206019|AIDS encephalopathy
C0206019|AIDS Encephalopathies
C0206019|Encephalopathies, AIDS
C0206019|Encephalopathies, HIV
C0206019|HIV Encephalopathies
C0206019|AIDS with encephalopathy
C0206019|Human immunodefiency virus encephalopathy
C0206019|AIDS with encephalopathy (disorder)
C0206019|HIV encephalopathy (diagnosis)
C0206019|Human immunodeficiency virus encephalopathy
C0206019|Human immunodeficiency virus encephalopathy (disorder)
C0206019|Human immunodefiency virus encephalopathy (disorder)
C0206019|Encephalopathy, HIV
C0206019|Encephalopathy, AIDS
C0206019|HIV disease; encephalopathy
C0206019|HIV disease; resulting in, encephalopathy
C0206019|encephalopathy; resulting from HIV disease
C0399449|HIV associated peridontitis
C0399449|HIV associated peridontitis (diagnosis)
C0399449|Human immunodeficiency virus-associated periodontitis
C0399449|Human immunodeficiency virus-associated periodontitis (disorder)
C0348990|HIV disease resulting in candidiasis
C0348990|HIV disease resulting in candidiasis (disorder)
C0348990|Human immunodeficiency virus (HIV) disease resulting in candidiasis (disorder)
C0348990|HIV infection resulting in candidiasis (diagnosis)
C0348990|HIV infection resulting in candidiasis
C0348990|Human immunodeficiency virus disease resulting in candidiasis (disorder)
C0348990|Human immunodeficiency virus (HIV) disease resulting in candidiasis
C0348990|Human immunodeficiency virus disease resulting in candidiasis
C0348990|HIV disease; candidiasis
C0348990|HIV disease; resulting in, candidiasis
C0348990|HIV disease; resulting in, infection, Candida
C0348990|candida; infection, resulting from HIV disease
C0348990|candidiasis; resulting from HIV disease
C0348990|infection; Candida, resulting from HIV disease
C0343747|Human immunodeficiency virus infection with neurological disease (disorder)
C0343747|Human immunodeficiency virus with neurological disease
C0343747|Human immunodeficiency virus infection with neurological disease
C0343747|Human immunodeficiency virus with neurological disease (disorder)
C0343747|HIV infection with neurological disease (diagnosis)
C0343747|HIV infection with neurological disease
C0348969|HIV disease resulting in mycobacterial infection
C0348969|HIV disease resulting in mycobacterial infection (disorder)
C0348969|Human immunodeficiency virus (HIV) disease resulting in mycobacterial infection (disorder)
C0348969|HIV infection resulting in mycobacterial infection (diagnosis)
C0348969|HIV infection resulting in mycobacterial infection
C0348969|Human immunodeficiency virus (HIV) disease resulting in mycobacterial infection
C0348969|Human immunodeficiency virus disease resulting in mycobacterial infection (disorder)
C0348969|Human immunodeficiency virus disease resulting in mycobacterial infection
C0348969|HIV disease; Mycobacterium
C0348969|HIV disease; resulting in, infection, mycobacterial
C0348969|HIV disease; resulting in, mycobacterial infection
C0348969|Mycobacterium; infection, resulting from HIV disease
C0348969|Mycobacterium; resulting from HIV disease
C0348969|infection; Mycobacterium, mycobacterial, resulting from HIV disease
C0348969|infection; tuberculous, resulting from HIV disease
C0348982|HIV disease resulting in cytomegaloviral disease
C0348982|HIV disease resulting in cytomegaloviral disease (disorder)
C0348982|Human immunodeficiency virus (HIV) disease resulting in cytomegaloviral disease (disorder)
C0348982|HIV infection resulting in cytomegaloviral infection
C0348982|HIV infection resulting in cytomegaloviral infection (diagnosis)
C0348982|Human immunodeficiency virus disease resulting in cytomegaloviral disease
C0348982|Human immunodeficiency virus disease resulting in cytomegaloviral disease (disorder)
C0348982|Human immunodeficiency virus (HIV) disease resulting in cytomegaloviral disease
C0348982|HIV disease; cytomegaloviral disease
C0348982|HIV disease; resulting in, cytomegaloviral disease
C0348982|HIV disease; resulting in, infection, cytomegaloviral
C0348982|cytomegaloviral disease; resulting from HIV disease
C0348821|HIV disease resulting in lymphoid interstitial pneumonitis
C0348821|HIV disease resulting in lymphoid interstitial pneumonitis (disorder)
C0348821|Human immunodeficiency virus (HIV) disease resulting in lymphoid interstitial pneumonitis (disorder)
C0348821|HIV infection resulting in lymphoid interstitial pneumonitis (diagnosis)
C0348821|HIV infection resulting in lymphoid interstitial pneumonitis
C0348821|Human immunodeficiency virus disease resulting in lymphoid interstitial pneumonitis
C0348821|Human immunodeficiency virus (HIV) disease resulting in lymphoid interstitial pneumonitis
C0348821|Human immunodeficiency virus disease resulting in lymphoid interstitial pneumonitis (disorder)
C0348821|HIV disease; resulting in, lymphoid interstitial pneumonitis
C0348821|HIV disease; resulting in, pneumonitis, interstitial, lymphatic
C0348207|HIV disease resulting in multiple infections
C0348207|HIV disease resulting in multiple infections (disorder)
C0348207|Human immunodeficiency virus (HIV) disease resulting in multiple infections (disorder)
C0348207|HIV infection resulting in multiple infections (diagnosis)
C0348207|HIV infection resulting in multiple infections
C0348207|Human immunodeficiency virus (HIV) disease resulting in multiple infections
C0348207|Human immunodeficiency virus disease resulting in multiple infections
C0348207|Human immunodeficiency virus disease resulting in multiple infections (disorder)
C0348207|HIV disease; resulting in multiple infections
C0348207|HIV disease; resulting in, infection, multiple
C0349036|HIV disease resulting in multiple malignant neoplasms
C0349036|HIV disease resulting in multiple malignant neoplasms (disorder)
C0349036|Human immunodeficiency virus (HIV) disease resulting in multiple malignant neoplasms
C0349036|Human immunodeficiency virus (HIV) disease resulting in multiple malignant neoplasms (disorder)
C0349036|HIV infection resulting in multiple malignant neoplasms
C0349036|HIV infection resulting in multiple malignant neoplasms (diagnosis)
C0349036|Human immunodeficiency virus disease resulting in multiple malignant neoplasms (disorder)
C0349036|Human immunodeficiency virus disease resulting in multiple malignant neoplasms
C0349036|HIV disease; resulting in, neoplasm, malignant, multiple
C0410223|HIV-associated myopathy
C0410223|HIV-associated myopathy (diagnosis)
C0410223|HIV associated myopathy
C0410223|HIV associated myopathy (diagnosis)
C0410223|HIV - Human immunodeficiency virus myopathy
C0410223|Human immunodeficiency virus myopathy
C0410223|Human immunodeficiency virus myopathy (disorder)
C0276500|HIV I infection
C0276500|HIV I infection (diagnosis)
C0276500|Human immunodeficiency virus I infection
C0276500|Human immunodeficiency virus I infection (disorder)
C0338422|HIV leukoencephalopathy (diagnosis)
C0338422|HIV leukoencephalopathy
C0338422|Human immunodeficiency virus leucoencephalopathy
C0338422|Human immunodeficiency virus leukoencephalopathy (disorder)
C0338422|Human immunodefiency virus leucoencephalopathy
C0338422|HIV - Human immunodeficiency virus leucoencephalopathy
C0338422|HIV - Human immunodeficiency virus leukoencephalopathy
C0338422|HIV - Human immunodefiency virus leukoencephalopathy
C0338422|HIV - Human immunodefiency virus leucoencephalopathy
C0338422|Human immunodefiency virus leukoencephalopathy
C0338422|Human immunodefiency virus leukoencephalopathy (disorder)
C0338422|Human immunodeficiency virus leukoencephalopathy
C0276501|HIV II infection
C0276501|HIV II infection (diagnosis)
C0276501|HIV 2 infection
C0276501|Human immunodeficiency virus II infection
C0276501|Human immunodeficiency virus II infection (disorder)
C0276548|HIV encephalitis
C0276548|AIDS with encephalitis
C0276548|AIDS with encephalitis (disorder)
C0276548|HIV - Human immunodefiency virus encephalitis
C0276548|Human immunodefiency virus subacute encephalitis
C0276548|Human immunodefiency virus encephalitis
C0276548|HIV encephalitis (diagnosis)
C0276548|HIV - Human immunodeficiency virus encephalitis
C0276548|Human immunodefiency virus encephalitis (disorder)
C0276548|Human immunodeficiency virus encephalitis
C0276548|Human immunodeficiency virus encephalitis (disorder)
C0452189|HIV disease resulting in Burkitt's lymphoma
C0452189|HIV disease resulting in Burkitt's lymphoma (disorder)
C0452189|Human immunodeficiency virus (HIV) disease resulting in Burkitt's lymphoma (disorder)
C0452189|HIV infection resulting in Burkitt's lymphoma
C0452189|HIV infection resulting in Burkitt's lymphoma (diagnosis)
C0452189|Human immunodeficiency virus disease resulting in Burkitt's lymphoma (disorder)
C0452189|Human immunodeficiency virus disease resulting in Burkitt's lymphoma
C0452189|Human immunodeficiency virus (HIV) disease resulting in Burkitt's lymphoma
C0452189|Human immunodeficiency virus (HIV) disease resulting in Burkitt lymphoma
C0452189|HIV disease; Burkitt
C0452189|HIV disease; lymphoma, Burkitt
C0452189|Burkitt; lymphoma, resulting from HIV disease
C0452189|lymphoma; Burkitt, resulting from HIV disease
C0276601|HIV infection with infection by another virus (disorder)
C0276601|Human immunodeficiency virus (HIV) infection with infection by another virus (disorder)
C0276601|HIV infection with infection by another virus
C0276601|HIV infection with infection by another virus (diagnosis)
C0276601|Human immunodeficiency virus infection with infection caused by another virus
C0276601|Human immunodeficiency virus (HIV) infection with infection by another virus
C0276601|Human immunodeficiency virus infection with infection caused by another virus (disorder)
C0276601|Human immunodeficiency virus (HIV) infection with infection caused by another virus
C0276601|Human immunodeficiency virus infection with infection by another virus (disorder)
C0276601|Human immunodeficiency virus infection with infection by another virus
C0276601|HIV infection with infection caused by another virus
C0276601|AIDS virus with viral infection
C0343756|Human immunodeficiency viral myelitis
C0343756|HIV myelitis
C0343756|HIV myelitis (diagnosis)
C0343756|HIV - Human immunodeficiency virus myelitis
C0343756|Human immunodeficiency virus myelitis
C0343756|Human immunodeficiency virus myelitis (disorder)
C0456101|hiv congenital positive status syndrome
C0456101|congenital HIV positive status syndrome (diagnosis)
C0456101|congenital HIV positive status syndrome
C0456101|Congenital human immunodeficiency virus positive status syndrome
C0456101|HIV - Congenital human immunodeficiency virus positive status syndrome
C0456101|Congenital human immunodeficiency virus positive status syndrome (disorder)
C0276599|HIV infection with acute lymphadenitis (disorder)
C0276599|Human immunodeficiency virus (HIV) infection with acute lymphadenitis
C0276599|Human immunodeficiency virus infection with acute lymphadenitis (disorder)
C0276599|Human immunodeficiency virus infection with acute lymphadenitis
C0276599|Human immunodeficiency virus (HIV) infection with acute lymphadenitis (disorder)
C0276599|AIDS virus with acute lymphadenitis (disorder)
C0276599|HIV infection with acute lymphadenitis
C0276599|AIDS virus with acute lymphadenitis
C0276599|hiv infection with acute lymphadenitis (diagnosis)
C0276602|HIV infection with infectious mononucleosis-like syndrome (disorder)
C0276602|Human immunodeficiency virus (HIV) infection with infectious mononucleosis-like syndrome
C0276602|Human immunodeficiency virus infection with infectious mononucleosis-like syndrome
C0276602|Human immunodeficiency virus (HIV) infection with infectious mononucleosis-like syndrome (disorder)
C0276602|Human immunodeficiency virus infection with infectious mononucleosis-like syndrome (disorder)
C0276602|HIV infection with infectious mononucleosis-like syndrome
C0276602|HIV infection with infectious mononucleosis-like syndrome (diagnosis)
C0276602|AIDS virus with "infectious mononucleosis-like syndrome"
C0343746|HIV infection with secondary clinically infectious disease
C0343746|HIV infection with secondary clinically infectious disease (diagnosis)
C0343746|Human immunodeficiency virus infection with secondary clinical infectious disease
C0343746|Human immunodeficiency virus infection with secondary clinical infectious disease (disorder)
C1319296|pediatric HIV infection
C1319296|hiv infection pediatric
C1319296|pediatric HIV infection (diagnosis)
C1319296|HIV infection, paediatric
C1319296|HIV infection, pediatric
C1319296|Paediatric human immunodeficiency virus infection
C1319296|Pediatric human immunodeficiency virus infection (disorder)
C1319296|Pediatric human immunodeficiency virus infection
C3840061|Human immunodeficiency virus in mother complicating childbirth (disorder)
C3840061|Human immunodeficiency virus in mother complicating childbirth
C3840061|HIV (human immunodeficiency virus) in childbirth
C3874345|Human immunodeficiency virus (HIV) infection category B2 (disorder)
C3874345|Human immunodeficiency virus (HIV) infection category B2
C3874330|Human immunodeficiency virus (HIV) infection category B1 (disorder)
C3874330|Human immunodeficiency virus (HIV) infection category B1
C3874341|Human immunodeficiency virus (HIV) II infection category B2
C3874341|Human immunodeficiency virus (HIV) II infection category B2 (disorder)
C4076110|Disorder of respiratory system co-occurrent with human immunodeficiency virus infection
C4076110|Disorder of respiratory system co-occurrent with human immunodeficiency virus infection (disorder)
C4076215|Infection caused by Salmonella co-occurrent with human immunodeficiency virus infection (disorder)
C4076215|Salmonellosis co-occurrent with human immunodeficiency virus infection
C4076215|Infection caused by Salmonella co-occurrent with human immunodeficiency virus infection
C4075735|Fever of unknown origin co-occurrent with human immunodeficiency virus infection
C4075735|Pyrexia of unknown origin co-occurrent with human immunodeficiency virus infection
C4075735|Pyrexia of unknown origin co-occurrent with human immunodeficiency virus infection (disorder)
C4075750|Infection caused by Aspergillus co-occurrent with human immunodeficiency virus infection
C4075750|Aspergillosis co-occurrent with human immunodeficiency virus infection
C4075750|Infection caused by Aspergillus co-occurrent with human immunodeficiency virus infection (disorder)
C4076090|Neuritis co-occurrent with human immunodeficiency virus infection
C4076090|Neuritis co-occurrent with human immunodeficiency virus infection (disorder)
C4075393|Immune reconstitution inflammatory syndrome caused by human immunodeficiency virus infection
C4075393|Immune reconstitution inflammatory syndrome caused by human immunodeficiency virus infection (disorder)
C4075812|Infection caused by herpes zoster virus co-occurrent with human immunodeficiency virus infection
C4075812|Herpes zoster infection co-occurrent with human immunodeficiency virus infection
C4075812|Infection caused by herpes zoster virus co-occurrent with human immunodeficiency virus infection (disorder)
C4075921|Disorder of central nervous system co-occurrent with human immunodeficiency virus infection (disorder)
C4075921|Disorder of central nervous system co-occurrent with human immunodeficiency virus infection
C4074813|Coccidiosis co-occurrent with human immunodeficiency virus infection
C4074813|Infection caused by Coccidia co-occurrent with human immunodeficiency virus infection (disorder)
C4074813|Infection caused by Coccidia co-occurrent with human immunodeficiency virus infection
C4076083|Hepatomegaly co-occurrent with human immunodeficiency virus infection
C4076083|Enlargement of liver co-occurrent with human immunodeficiency virus infection
C4076083|Enlargement of liver co-occurrent with human immunodeficiency virus infection (disorder)
C4076083|Large liver co-occurrent with human immunodeficiency virus infection
C4076016|Disorder of peripheral nervous system co-occurrent with human immunodeficiency virus infection (disorder)
C4076016|Disorder of peripheral nervous system co-occurrent with human immunodeficiency virus infection
C4075583|Disseminated atypical infection caused by Mycobacterium co-occurrent with human immunodeficiency virus infection
C4075583|Disseminated atypical infection caused by Mycobacterium co-occurrent with human immunodeficiency virus infection (disorder)
C4076290|Splenomegaly co-occurrent with human immunodeficiency virus infection (disorder)
C4076290|Splenomegaly co-occurrent with human immunodeficiency virus infection
C4076117|Infection caused by Pneumocystis co-occurrent with human immunodeficiency virus infection
C4076117|Infection caused by Pneumocystis co-occurrent with human immunodeficiency virus infection (disorder)
C4076117|Pneumocystosis co-occurrent with human immunodeficiency virus infection
C4076026|Infective arthritis co-occurrent with human immunodeficiency virus infection (disorder)
C4076026|Infective arthritis co-occurrent with human immunodeficiency virus infection
C4075796|Infection caused by herpes simplex virus co-occurrent with human immunodeficiency virus infection (disorder)
C4075796|Herpes simplex virus infection co-occurrent with human immunodeficiency virus infection
C4075796|Infection caused by herpes simplex virus co-occurrent with human immunodeficiency virus infection
C4075629|Microsporidiosis co-occurrent with human immunodeficiency virus infection
C4075629|Infection caused by Microsporidia co-occurrent with human immunodeficiency virus infection (disorder)
C4075629|Infection caused by Microsporidia co-occurrent with human immunodeficiency virus infection
C4075653|Opportunistic mycosis co-occurrent with human immunodeficiency virus infection
C4075653|Opportunistic mycosis co-occurrent with human immunodeficiency virus infection (disorder)
C4076086|Candidiasis of mouth co-occurrent with human immunodeficiency virus infection (disorder)
C4076086|Candidiasis of mouth co-occurrent with human immunodeficiency virus infection
C4076155|Hemophagocytic syndrome co-occurrent with human immunodeficiency virus infection
C4076155|Hemophagocytic syndrome co-occurrent with human immunodeficiency virus infection (disorder)
C4075982|Nocardiosis co-occurrent with human immunodeficiency virus infection
C4075982|Infection caused by Nocardia co-occurrent with human immunodeficiency virus infection (disorder)
C4075982|Infection caused by Nocardia co-occurrent with human immunodeficiency virus infection
C4076042|Visual impairment co-occurrent with human immunodeficiency virus infection (disorder)
C4076042|Visual impairment co-occurrent with human immunodeficiency virus infection
C4075766|Infection caused by Cytomegalovirus co-occurrent with human immunodeficiency virus infection
C4075766|Infection caused by Cytomegalovirus co-occurrent with human immunodeficiency virus infection (disorder)
C4075766|Cytomegalovirus infection co-occurrent with human immunodeficiency virus infection
C4075814|Dermatophytosis co-occurrent with human immunodeficiency virus infection
C4075814|Infection caused by Dermatophyte co-occurrent with human immunodeficiency virus infection
C4075814|Infection caused by Dermatophyte co-occurrent with human immunodeficiency virus infection (disorder)
C4076115|Polyneuropathy co-occurrent with human immunodeficiency virus infection
C4076115|Polyneuropathy co-occurrent with human immunodeficiency virus infection (disorder)
C4076275|Disorder of eye proper co-occurrent with human immunodeficiency virus infection
C4076275|Disorder of eye proper co-occurrent with human immunodeficiency virus infection (disorder)
C4076275|Disorder of eye co-occurrent with human immunodeficiency virus infection
C4076216|Anaemia co-occurrent with human immunodeficiency virus infection
C4076216|Anemia co-occurrent with human immunodeficiency virus infection (disorder)
C4076216|Anemia co-occurrent with human immunodeficiency virus infection
C4076274|Heart disease co-occurrent with human immunodeficiency virus infection (disorder)
C4076274|Heart disease co-occurrent with human immunodeficiency virus infection
C4075781|Infection caused by Strongyloides co-occurrent with human immunodeficiency virus infection (disorder)
C4075781|Infection caused by Strongyloides co-occurrent with human immunodeficiency virus infection
C4075781|Strongyloidiasis co-occurrent with human immunodeficiency virus infection
C4076265|Disorder of gastrointestinal tract co-occurrent with human immunodeficiency virus infection
C4076265|Disorder of gastrointestinal tract co-occurrent with human immunodeficiency virus infection (disorder)
C4076101|Lymphadenopathy co-occurrent with human immunodeficiency virus infection
C4076101|Lymphadenopathy co-occurrent with human immunodeficiency virus infection (disorder)
C4075933|Malignant neoplastic disease co-occurrent with human immunodeficiency virus infection (disorder)
C4075933|Malignant neoplastic disease co-occurrent with human immunodeficiency virus infection
C4076103|Nephropathy co-occurrent with human immunodeficiency virus infection
C4076103|Disorder of kidney co-occurrent with human immunodeficiency virus infection
C4076103|Disorder of kidney co-occurrent with human immunodeficiency virus infection (disorder)
C4076222|Disorder of skin co-occurrent with human immunodeficiency virus infection (disorder)
C4076222|Disorder of skin co-occurrent with human immunodeficiency virus infection
C4076020|Agranulocytosis co-occurrent with human immunodeficiency virus infection (disorder)
C4076020|Agranulocytosis co-occurrent with human immunodeficiency virus infection
C0856916|Persistent generalised lymphadenopathy
C0856916|Persistant generalized lymphadenopathy
C0856916|Persistant generalised lymphadenopathy
C0856916|PLG
C0856916|lymphadenopathy persistent generalized (diagnosis)
C0856916|lymphadenopathy persistent generalized
C0856916|Persistent generalized lymphadenopathy
C0856916|Human immunodeficiency virus infection with persistent generalised lymphadenopathy
C0856916|Human immunodeficiency virus infection with persistent generalized lymphadenopathy
C0856916|PGL - Persistent generalised lymphadenopathy
C0856916|PGL - Persistent generalized lymphadenopathy
C0856916|Persistent generalized lymphadenopathy (disorder)
C0686714|AIDS virus infection associated with pregnancy (disorder)
C0686714|Acquired immunodeficiency syndrome (AIDS) virus infection associated with pregnancy
C0686714|Acquired immunodeficiency syndrome virus infection associated with pregnancy (disorder)
C0686714|Acquired immunodeficiency syndrome (AIDS) virus infection associated with pregnancy (disorder)
C0686714|Acquired immunodeficiency syndrome virus infection associated with pregnancy
C0686714|AIDS virus infection associated with pregnancy
C0559284|HIV-related gut disease - cause unknown (disorder)
C0559284|Human immunodeficiency virus HIV-related gut disease - cause unknown (disorder)
C0559284|Human immunodeficiency virus-related gut disease - cause unknown (disorder)
C0559284|HIV-related gut disease - cause unknown
C0559284|Human immunodeficiency virus HIV-related gut disease - cause unknown
C0559284|Human immunodeficiency virus-related gut disease - cause unknown
C0559283|HIV-related sclerosing cholangitis (disorder)
C0559283|Human immunodeficiency virus HIV-related sclerosing cholangitis
C0559283|Human immunodeficiency virus-related sclerosing cholangitis (disorder)
C0559283|Human immunodeficiency virus-related sclerosing cholangitis
C0559283|Human immunodeficiency virus HIV-related sclerosing cholangitis (disorder)
C0559283|sclerosing cholangitis human immunodeficiency virus-realted
C0559283|Human immunodeficiency virus-related sclerosing cholangitis (diagnosis)
C0559283|HIV-related sclerosing cholangitis
C0276605|Positive serological or viral culture findings for human ummunodeficiency virus
C0276605|Positive serological AND/OR viral culture findings for human immunodeficiency virus (disorder)
C0276605|Positive serological AND/OR viral culture findings for human immunodeficiency virus
C0276605|Positive serological or viral culture findings for human immunodeficiency virus
C0348204|HIV disease resulting in other bacterial infections
C0348204|[X]HIV disease resulting in other bacterial infections
C0348204|[X]HIV disease resulting in other bacterial infections (disorder)
C0348204|bacterial; infection, resulting from HIV disease
C0348204|infection; bacterial, resulting from HIV disease
C0348212|HIV disease resulting in other malignant neoplasms
C0348212|[X]HIV disease resulting in other malignant neoplasms
C0348212|[X]HIV disease resulting in other malignant neoplasms (disorder)
C0348206|HIV disease resulting in other mycoses
C0348206|[X]HIV disease resulting in other mycoses (disorder)
C0348206|[X]HIV disease resulting in other mycoses
C0348206|HIV disease; mycosis
C0348206|HIV disease; resulting in, infection, fungus
C0348206|HIV disease; resulting in, infection, mycotic
C0348206|HIV disease; resulting in, mycosis
C0348206|fungus; infection, resulting from HIV disease
C0348206|infection; fungus, resulting from HIV disease
C0348206|infection; mycotic, resulting from HIV disease
C0348206|mycosis; resulting from HIV disease
C0348206|mycotic; infection, resulting from HIV disease
C0348210|[X]HIV disease resulting in other non-Hodgkin's lymphoma
C0348210|[X]HIV disease resulting in other non-Hodgkin's lymphoma (disorder)
C0276555|HIV disease resulting in other specified conditions
C0276555|AIDS with other specified conditions -RETIRED-
C0276555|AIDS with other specified conditions
C0276555|[X]HIV disease resulting in other specified conditions (disorder)
C0276555|AIDS with other specified conditions (disorder)
C0276555|[X]HIV disease resulting in other specified conditions
C0348205|HIV disease resulting in other viral infections
C0348205|[X]HIV disease resulting in other viral infections
C0348205|[X]HIV disease resulting in other viral infections (disorder)
C0348215|[X]Hiv disease resulting in hematological and immunological abnormalities, not elsewhere classified
C0348215|[X]Hiv disease resulting in haematological and immunological abnormalities, not elsewhere classified
C0348215|[X]Hiv disease resulting in haematological and immunological abnormalities, not elsewhere classified (disorder)
C0348215|[X]Hiv disease resulting in hematological and immunological abnormalities, not elsewhere classified (disorder)
C0348215|[X]Hiv disease resulting in haematological and immunological abnormalities, NEC (disorder) in SNOMEDCT_US_2016_03_01
C0348211|HIV disease resulting in other malignant neoplasms of lymphoid, haematopoietic and related tissue
C0348211|HIV disease resulting in other malignant neoplasms of lymphoid, hematopoietic and related tissue
C0348211|[X]Hiv disease resulting in other malignant neoplasms of lymphoid, hematopoietic and related tissue
C0348211|[X]Hiv disease resulting in other malignant neoplasms of lymphoid, hematopoietic and related tissue (disorder)
C0348211|[X]Hiv disease resulting in other malignant neoplasms of lymphoid, haematopoietic and related tissue (disorder)
C0348211|[X]Hiv disease resulting in other malignant neoplasms of lymphoid, haematopoietic and related tissue
C0348214|HIV disease resulting in multiple diseases classified elsewhere
C0348214|[X]HIV disease resulting in multiple diseases classified elsewhere (disorder)
C0348214|[X]HIV disease resulting in multiple diseases classified elsewhere
C0348214|HIV disease; resulting in, multiple, diseases classified elsewhere
C0393489|Vacuolar myelopathy
C0393489|Vacuolar myelopathy (disorder)
C0456100|AIDS - Congenital acquired immune deficiency syndrome
C0456100|Congenital acquired immune deficiency syndrome
C0456100|Congenital acquired immune deficiency syndrome (disorder)
C1562915|uveitis immune recovery
C1562915|Immune recovery uveitis
C1562915|Immune recovery uveitis (diagnosis)
C1562915|Immune recovery uveitis (disorder)
C0276528|AIDS with viral pneumonia (disorder)
C0276528|Viral pneumonia associated with AIDS
C0276528|Acquired immunodeficiency syndrome (AIDS) with viral pneumonia
C0276528|AIDS with viral pneumonia
C0276528|Acquired immunodeficiency syndrome (AIDS) with viral pneumonia (disorder)
C0276528|Viral pneumonia associated with AIDS (diagnosis)
C0276528|pneumonia viral associated with aids
C0276528|Viral pneumonia associated with acquired immunodeficiency syndrome
C0276528|Viral pneumonia associated with acquired immunodeficiency syndrome (disorder)
C0276528|Viral pneumonia associated with AIDS (disorder)
C0276528|AIDS with viral pneumonia, NOS
C1720105|AIDS-associated disorder
C1720105|Complication of AIDS
C1720105|AIDS complication
C1720105|Acquired immunodeficiency syndrome-associated disorder (disorder)
C1720105|AIDS-associated disorder (disorder)
C1720105|Acquired immunodeficiency syndrome-associated disorder
