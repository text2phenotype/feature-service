1|%
2|10*12/l
3|10*3
4|10*3 iu/24 h
5|10*3 iu/l
6|10*3/mm3
7|10*3/ul
8|10*6
9|10*6 eq/ml
10|10*6/d
11|10*6/l
12|10*6/ml
13|10*6/ul
14|10*9/l
15|10*9/ul
16|10-9 mol/l
17|acu/ml
18|akat
19|angstrom
20|aru
21|attct repeats
22|au/ml
23|beats/min
24|bp
25|breaths/min
26|cells/ul
27|cfu/g
28|cgg repeats
29|cgy
30|ch 100 units/ml
31|ch 50 u/ml
32|clock time
33|cm
34|cm h2o
35|cm/cm
36|cm/s
37|cm2
38|cm3
39|coefficient of variation
40|copies
41|copies/l
42|copies/ml
43|copies/ul
44|cp
45|cpm
46|ctcs/7.5 ml
47|ctg repeats
48|d
49|dapa
50|days
51|days/12 mo
52|days/3 mo
53|days/30 days
54|days/5 days
55|days/7 days
56|days/mo
57|days/week
58|deg
59|deg c
60|deg f
61|dils
62|diopter
63|dye units
64|dyn.s/cm5
65|ehrlich units/100 g
66|ehrlich units/24 h
67|ehrlich units/dl
68|eia index
69|eia units
70|elisa index
71|elisa units
72|eq/ml
73|ery/ul
74|eu
75|eu/ml
76|eus
77|feet/day
78|feet/week
79|fl
80|fl/nl
81|fmol
82|fmol/l
83|fmol/mg
84|fmol/mg protein
85|fraction
86|ft
87|ft-in
88|ft/ft
89|g
90|g/10 h
91|g/100 g
92|g/12 h
93|g/18 h
94|g/2 h
95|g/24 h
96|g/4 h
97|g/48 h
98|g/5 h
99|g/6 h
100|g/72 h
101|g/8 h
102|g/cm2
103|g/d
104|g/dl
105|g/g creatinine
106|g/kg
107|g/l
108|g/ml
109|g/mmol
110|g/mmol creatinine
111|gaa repeats
112|gf/cm2
113|gm
114|gm/l
115|gm/mmol_cre
116|gpl u
117|gps u
118|grams
119|h
120|hhmm
121|hhmm/night
122|hours
123|hours/5 days
124|hours/days
125|hours/night
126|hours/session
127|hours/week
128|hr
129|hz
130|ifa titer
131|in
132|index
133|index value
#134|inr
135|isr
136|iu/24 h
137|iu/24h
138|iu/dl
139|iu/g creatinine
140|iu/l
141|iu/ml
142|kcal
143|kcal/24 h
144|kcal/24h
145|kcal/day
146|kcal/week
147|kd/s
148|keu/l
149|kg
150|kg/m2
151|kilometers
152|kiu/l
153|kiu/ml
154|km
155|km/24 h
156|km/24h
157|km/h
158|km/wk
159|kpa
160|ku/l
161|ku/ml
162|l
163|l/24 h
164|l/24h
165|l/l
166|l/min
167|l/s
168|lb
169|lb-oz
170|lb/d
171|lbf
172|leu/ul
173|liley unit
174|liters
175|liv
176|log copies/ml
177|log iu/ml
178|log reduction
179|lu
180|m
181|m-cm
182|m.o.m
183|m/6 min
184|m/s
185|m2
186|mcg/100mg
187|mcg/dl
188|mcg/g creatinine
189|mcg/gm
190|mcg/gm cr
191|mcg/l
192|mcg/mg cr
193|mcg/ml
194|mcmol/dl
195|mcmol/l
196|mcu/ml
197|meq/12h
198|meq/24 h
199|meq/d
200|meq/g
201|meq/g creatinine
202|meq/kg
203|meq/kg liq stl
204|meq/l
205|mg
206|mg/100 g
207|mg/100g
208|mg/12 h
209|mg/12h
210|mg/18 h
211|mg/18h
212|mg/2 h
213|mg/2h
214|mg/24 h
215|mg/24h
216|mg/24h
217|mg/4 h
218|mg/4h
219|mg/48 h
220|mg/48h
221|mg/6 h
222|mg/6h
223|mg/72 h
224|mg/72h
225|mg/d
226|mg/dl
227|mg/g
228|mg/h
229|mg/kg
230|mg/l
231|mg/m3
232|mg/ml
233|mg2/dl2
234|mi
235|mi/24 h
236|mi/24h
237|mi/h
238|mi/wk
239|miles
240|min
241|min/d
242|minutes
243|miu/24 h
244|miu/24h
245|miu/l
246|miu/ml
247|mj
248|mkat/l
249|ml/24 h
250|ml/24h
251|ml/7 d
252|ml/7d
253|ml/72 h
254|ml/72h
255|ml/beat
256|ml/dl
257|ml/kg
258|ml/lb
259|ml/min
260|ml/s
261|ml/sec
262|mm
263|mm/15 min
264|mm/15min
265|mm/2 h
266|mm/2h
267|mm/h
268|mm/mm
269|mm2
270|mm3
271|mmddyy
272|mmol
273|mmol/100 g
274|mmol/100g
275|mmol/12 h
276|mmol/12h
277|mmol/18 h
278|mmol/18h
279|mmol/2 h
280|mmol/2h
281|mmol/24 h
282|mmol/24h
283|mmol/4 h
284|mmol/4h
285|mmol/5 h
286|mmol/5h
287|mmol/6 h
288|mmol/6h
289|mmol/72 h
290|mmol/72h
291|mmol/cp
292|mmol/d
293|mmol/dl
294|mmol/g
295|mmol/h
296|mmol/kg
297|mmol/l
298|mmol/ml
299|mmol/mmol
300|mmol/mol
301|mmol2/l2
302|mmyyyy
303|mo
304|mo/year
305|mol/24 h
306|mol/24h
307|mol/kg
308|mol/l
309|mol/mol
310|mosm/kg
311|mosm/kg water
312|mosm/l
313|mosmol/kg
314|mph
315|mpl u
316|mps u
317|ms
318|mu/g hb
319|mu/l
320|mu/ml
321|mu/mmol creatinine
322|mv
323|mv/s
324|mw
325|ng ab n/ml
326|ng/24 h
327|ng/dl
328|ng/g
329|ng/g creatinine
330|ng/l
331|ng/l
332|pg/ml
333|pmol/l
334|ng/l
335|pmol/l
336|ng/mg creatinine
337|ng/ml
338|ng/mol creatinine
339|ng/ng
340|ng/ng creatinine
341|nm
342|nmol bce/l
343|nmol/10*7
344|nmol/10*9
345|nmol/24 h
346|nmol/d
347|nmol/dl
348|nmol/g
349|nmol/g creatinine
350|nmol/g hb
351|nmol/kg faeces
352|nmol/l
353|nmol/mg
354|nmol/mg creatinine
355|nmol/mg protein
356|nmol/min
357|nmol/ml
358|nmol/ml rbc
359|nmol/mmo
360|nmol/mmol
361|nmol/mmol creat
362|nmol/mmol creatinine
363|nmol/mol creatinine
364|nmol/nmol
365|nmole/mmole_cr
366|nmoles/ml
367|od ratio
368|od units
369|osm/kg
370|oz
371|oz/wk
372|peiu/ml
373|pg
374|pg/dl
375|pg/g creatinine
376|pg/mg creatinine
377|pg/ml
378|pg/ml slt
379|pg/pg
380|ph
381|pmol/24 h
382|pmol/24h
383|pmol/8x10*8 rbc
384|pmol/g
385|pmol/l
386|pmol/ml
387|pmol/mol
388|pmol/mol creatinine
389|ppb
390|ppg
391|ppm
392|pru
393|psi
394|ratio
395|rbc/min
396|rbcs/ul
397|rev
398|rfu
399|risk
400|ru
401|ru/ml
402|score
403|sd
404|si
405|thous miu/ml
406|titer
407|tmstp
408|todd units
409|tscore
410|u/10*10 cells
411|u/10*12
412|u/12 h
413|u/12h
414|u/18 h
415|u/18h
416|u/2 h
417|u/2h
418|u/24 h
419|u/24h
420|u/d
421|u/dl
422|u/g
423|u/g creatinine
424|u/g hb
425|u/g protein
426|u/gm
427|u/h
428|u/kg
429|u/kg bw
430|u/kg hb
431|u/kg hgb
432|u/l
433|u/mg protein
434|u/ml
435|u/ml rbc
436|u/u
437|ug
438|ug eq/ml
439|ug/100g dry wt
440|ug/12 h
441|ug/24 h
442|ug/72 h
443|ug/8 h
444|ug/dl
445|ug/dl
446|nmol/l
447|ug/g
448|ug/g cre
449|ug/g creatinine
450|ug/g hb
451|ug/kg
452|ug/l
453|ug/l ddu
454|ug/l feu
455|ug/m3
456|ug/mg creatinine
457|ug/min
458|ug/ml
459|ug/ml equivalents
460|ug/ml feu
461|ug/mmol creatinine
462|ug/ug
463|ug/ul
464|ui/l
465|uiu/l
466|uiu/ml
467|ukat/l
468|um
469|um/gcr
470|um/s
471|umol/2 h
472|umol/2h
473|umol/24 h
474|umol/24h
475|umol/d
476|umol/dl
477|umol/ejaculate
478|umol/g
479|umol/g creatinine
480|umol/kg
481|umol/l
482|umol/ml
483|umol/mmol
484|umol/mmol creatinine
485|umol/mol
486|umol/mol cr
487|umol/mol crea
488|umol/mol creat
489|umol/mol creatinine
490|umol/mol hb
491|umol/umol
492|umole/l
493|units/l
494|units/ml
495|uu/ml
496|wbc/min
497|wbcs/ul
498|mgAlb/gCre
499|uug
500|um3
501|k/ul
502|m/ul
503|inches
504|pounds
505|pound
