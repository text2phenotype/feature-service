C2910651|Unknown Route of HCV Transmission
C2910651|Unknown Route of HCV Infection 
C2910651|Contact with and (suspected) exposure to viral hepatitis
C2910651|Contact with viral hepatitis
C2910651|Contact with hepatitis C virus  
C2910651|Contact with viral hepatitis
C2910651|Contact with HCV
C2919618|Exposure to HCV
C2919618|Exposure to Hepatitis C
C2919618|Exposure to Hepatitis C virus
C2910651|Contact with and (suspected) exposure to viral hepatitis
C1096517|exposure to hepatitis C (history)
C1096517|exposure to hepatitis C
C1096517|Hepatitis C exposure
