C0011570|Mental Depression
C0011581|Depressive disorder
C0344315|Depressed mood
C0460137|Depression motion
C0812393|Cancer patients and suicide and depression
C1579931|Depressed - symptom
C1999266|Depression Adverse Event
C4049644|Depression Scale (BASC-2)
C4084909|Depression Subordinate Domain
C4085311|Depression - recess
C0743072|psychotic depression
C0743072|depressive psychosis
C0743072|Depression;psychotic
C0743072|Psychosis;depressive
C0743072|Depressive psychoses
C0743072|Depression, psychotic
C0743072|Depression psychotic
C0743072|Psychosis depressive
C0743072|depression; psychotic
C0743072|depressive; psychosis
C0743072|psychosis; depressive
C0743072|psychotic; depression
C0541868|Depression functional
C0541869|Depression worsened
C0221074|Postpartum depression
C0221074|Depression, Post-Natal
C0221074|Depression, Post-Partum
C0221074|Depression, Postnatal
C0221074|Depression, Postpartum
C0221074|Post Natal Depression
C0221074|Post Partum Depression
C0221074|postpartum depression (diagnosis)
C0221074|Depression, Postpartum [Disease/Finding]
C0221074|Post-Natal Depression
C0221074|Post-Partum Depression
C0221074|Postnatal Depression
C0221074|Depression;postnatal
C0221074|Depression;puerperal
C0221074|Depression postpartum (excl psychosis)
C0221074|[X]Postnatal depression NOS
C0221074|[X]Postpartum depression NOS
C0221074|Depression - postnatal
C0221074|Postnatal depressive disorder (disorder)
C0221074|Postnatal depressive disorder
C0221074|Depressive Episode with Postpartum Onset
C0221074|Major Depressive Episode with Peripartum Onset
C0221074|Postnatal blues
C0221074|Postnatal depression (excl psychosis)
C0221074|Depression puerperal
C0221074|Puerperal depression
C0221074|Postnatal depression (excluding psychosis)
C0221074|Postpartum depression (disorder)
C0221074|depression; postnatal
C0221074|depression; postpartum
C0221074|postnatal; depression
C0221074|postpartum; depression
C0221074|Depression postpartum (excluding psychosis)
C0494397|Mild depressive episode
C0494397|[X]Mild depressive episode (disorder)
C0494397|[X]Mild depressive episode
C0494397|episode; depressive, mild
C0494398|Moderate depressive episode
C0494398|[X]Moderate depressive episode (disorder)
C0494398|[X]Moderate depressive episode
C0494398|episode; depressive, moderate
C0154411|Major depressive disorder, recurrent episode, moderate degree
C0154411|Recurrent depressive disorder, current episode moderate
C0154411|moderate recurrent major depression (diagnosis)
C0154411|moderate recurrent major depression
C0154411|Recurr depr psychos-mod
C0154411|Major depressive disorder, recurrent, moderate
C0154411|Major depressive affective disorder, recurrent episode, moderate
C0154411|[X]Recurrent depressive disorder, current episode moderate (disorder)
C0154411|[X]Recurrent depressive disorder, current episode moderate
C0154411|Moderate recurrent major depression (disorder)
C0235876|Depression aggravated
C0236764|recurrent major depression in partial remission
C0236764|recurrent major depression in partial remission (diagnosis)
C0236764|Major depressive disorder, recurrent, in partial remission
C0236764|Recurrent major depression in partial remission (disorder)
C0041696|Depressions, Unipolar
C0041696|Unipolar Depressions
C0041696|Unipolar Depression
C0041696|Major Depressive Disorder
C0041696|Major Depression
C0041696|Unipolar depressive illness
C0041696|Depression, Unipolar
C0154403|Major depressive disorder, single episode, mild degree
C0154403|mild single episode major depression (diagnosis)
C0154403|mild single episode major depression
C0154403|Depress psychosis-mild
C0154403|Major depressive disorder, single episode, mild
C0154403|Major depressive affective disorder, single episode, mild
C0154403|Mild major depression, single episode
C0154403|Single major depressive episode, mild
C0154403|Mild major depression, single episode (disorder)
C0154403|Single major depressive episode, mild (disorder)
C0154403|disorder; depressive, major, single episode, mild
C0154404|Major depressive disorder, single episode, moderate degree
C0154404|moderate single episode major depression (diagnosis)
C0154404|moderate single episode major depression
C0154404|Depressive psychosis-mod
C0154404|Major depressive disorder, single episode, moderate
C0154404|Major depressive affective disorder, single episode, moderate
C0154404|Moderate major depression, single episode
C0154404|Single major depressive episode, moderate
C0154404|Moderate major depression, single episode (disorder)
C0154404|Single major depressive episode, moderate (disorder)
C0154404|disorder; depressive, major, single episode, moderate
C3665435|Major depressive disorder, recurrent episode, mild degree
C3665435|Recurr depr psychos-mild
C3665435|Major depressive affective disorder, recurrent episode, mild
C3665435|major depression, recurrent, mild episode
C3665435|recurrent major depressive episode, mild (diagnosis)
C3665435|recurrent major depressive episode, mild
C3665435|Recurrent major depressive episodes, mild
C3665435|Recurrent major depressive episodes, mild (disorder)
C0154412|Major depressive disorder, recurrent episode, severe degree, without mention of psychotic behavior
C0154412|Recurrent depressive disorder, current episode severe without psychotic symptoms
C0154412|severe recurrent major depression without psychotic features
C0154412|severe recurrent major depression without psychotic features (diagnosis)
C0154412|Recur depr psych-severe
C0154412|Major depressive disorder, recurrent severe without psychotic features
C0154412|Major depressv disorder, recurrent severe w/o psych features
C0154412|Major depressive affective disorder, recurrent episode, severe, without mention of psychotic behavior
C0154412|[X]Major depression, recurrent without psychotic symptoms
C0154412|[X]Recurrent depressive disorder, current episode severe without psychotic symptoms
C0154412|[X]Recurrent depressive disorder, current episode severe without psychotic symptoms (disorder)
C0154412|Severe recurrent major depression without psychotic features (disorder)
C0270455|Mild major depression
C0270455|major depression mild
C0270455|Mild major depression (diagnosis)
C0270455|Mild major depression (disorder)
C0235136|Agitated depression
C0235136|Agitated depression (disorder)
C0235136|Agitated depression (diagnosis)
C0235136|depression agitated
C0235136|depression; agitated
C0235136|agitated; depression
C0011570|Depressions
C0011570|Depression
C0011570|Mental Depression
C0011570|Depression psychic
C0011570|Monopolar depression NOS
C0011570|Depression NOS
C0011570|[X] Depression NOS
C0011570|Depression NOS (disorder)
C0011570|Depression (finding)
C0011570|[X]Depression NOS
C0011570|Depression, Mental
C0011570|Depressed Mood
C0011570|Depression mental
C0011570|Depressive state
C0011570|Depressed state
C0011570|depression; mental
C0011570|depression; monopolar
C0011570|depressive; state
C0011570|mental; depression
C0011570|monopolar; depression
C0011570|state; depressive
C0011570|Depression, NOS
C0011570|Depression (Emotion)
C0011570|Depressive state NOS
C0011570|Disorder;depression
C1269683|MAJOR DEPRESSIVE DISORDER
C1269683|major depression
C1269683|Disorder, Major Depressive
C1269683|Disorders, Major Depressive
C1269683|Major Depressive Disorders
C1269683|MDD
C1269683|DEPRESSIVE DIS MAJOR
C1269683|MAJOR DEPRESSIVE DIS
C1269683|Major depression NOS
C1269683|Depressive Disorder, Major [Disease/Finding]
C1269683|Depressive Disorder, Major
C1269683|Major depressive disorder (diagnosis)
C1269683|Major depressive disorder NOS
C1269683|Major depressive illness
C1269683|Major depressive disorder (disorder)
C1269683|Major depression, NOS
C1269683|Major depressive disorder, NOS
C1269683|Depressive Disorders, Major
C0086132|Depression, Emotional
C0086132|Depressions, Emotional
C0086132|Depressive Symptom
C0086132|Emotional Depressions
C0086132|Symptom, Depressive
C0086132|Symptoms, Depressive
C0086132|Symptoms of depression
C0086132|Symptoms of depression (finding)
C0086132|Depressive symptoms
C0086132|Emotional Depression
C2700639|[X] (Depression: [episode, unspecified] or [NOS (& reactive)] or [depressive disorder NOS] (disorder)
C2700639|[X] (Depression: [episode, unspecified] or [NOS (& reactive)] or [depressive disorder NOS]
C2363919|Childhood depression
C0270458|severe major depressive disorder with psychotic features
C0270458|major depression severe with psychotic features
C0270458|severe major depressive disorder with psychotic features (diagnosis)
C0270458|Severe major depression with psychotic features
C0270458|Psychotic depression
C0270458|Severe major depression with psychotic features (disorder)
C0270458|Severe major depression with psychotic features, NOS
C0270458|Psychotic depression, NOS
C0011579|Depressions, Reactive
C0011579|Reactive Depressions
C0011579|Neurotic Depressive Reaction
C0011579|Reactive Depression
C0011579|Reactive depression (situational) (finding)
C0011579|Reactive depression (situational) (disorder)
C0011579|Depression;reactive
C0011579|reactive depression (diagnosis)
C0011579|Reactive (neurotic) depression
C0011579|[X] Reactive depression NOS
C0011579|[X]Prolonged single episode of reactive depression
C0011579|Neurotic depression reactive type
C0011579|Depressive reaction
C0011579|Depression reactive
C0011579|Reactive depression (situational)
C0011579|depression; reactive
C0011579|depressive; reaction
C0011579|reaction; depressive
C0011579|reactive; depression
C0011579|Depressive Reaction (Neurotic)
C0011579|Depression, Reactive
C2362914|clinical depression
C0013415|Dysthymia
C0013415|Dysthymic Disorder
C0013415|Dysthymic Disorders
C0013415|Disorder, Dysthymic
C0013415|DYSTHYMIC DIS
C0013415|dysthymia (diagnosis)
C0013415|Dysthymic Disorder [Disease/Finding]
C0013415|Dysthymia (disorder)
C0013415|persistent depressive disorder (dysthymia) (diagnosis)
C0013415|persistent depressive disorder (dysthymia)
C0013415|disorder; dysthymic
C0013415|dysthymic; disorder
C0013415|Dysthymia, NOS
C0344315|Depressed mood
C0344315|depressed mood (physical finding)
C0344315|mood depressed
C0344315|Low mood
C0344315|Depressed mood (finding)
C0344315|Feeling low
C0344315|Morose mood
C0344315|Morose mood (finding)
C0344315|Miserable
C0344315|Depressed
C0344315|Morosity
C0344315|Melancholic
C0344315|Decreased Mood
C0344315|Feeling blue
C0344315|Feeling down
C0344315|Mood depressions
C0344315|Mood depression
C0344315|Melancholy
C0344315|Feeling;down
C1868594|PERRY SYNDROME
C1868594|Parkinsonism with Alveolar Hypoventilation and Mental Depression
C1868594|Perry syndrome (disorder)
C0455770|Loss (of);feeling
C0455770|Feeling of loss of feeling
C0455770|Feeling of loss of feeling (finding)
C0455770|loss of feeling
C0349217|Depressive episode, unspecified
C0349217|Depressive episode
C0349217|[X]Depressive episode, unspecified
C0349217|[X]Depressive episode, unspecified (disorder)
C0349217|depressive; episode
C0349217|episode; depressive
C0812393|Cancer patients and suicide and depression
C0812393|depression
C0812393|suicide
C0812393|cancer patients and depression and suicide
C0812393|depression and suicide
C0812393|suicide and depression
C0494399|Severe depressive episode without psychotic symptoms
C0494399|[X]Severe depressive episode without psychotic symptoms
C0494399|[X]Severe depressive episode without psychotic symptoms (disorder)
C0494399|depressive; disorder, major, single episode, major (without psychotic symptoms)
C0494399|depressive; episode, severe (without psychotic symptoms)
C0494399|disorder; depressive, major, single episode, major (without psychotic symptoms)
C0494399|episode; depressive, severe (without psychotic symptoms)
C0494400|Severe depressive episode with psychotic symptoms
C0494400|[X]Severe depressive episode with psychotic symptoms
C0494400|[X]Severe depressive episode with psychotic symptoms (disorder)
C0494400|depressive; disorder, major, single episode, major, with psychotic symptoms
C0494400|depressive; episode, severe, with psychotic symptoms
C0494400|disorder; depressive, major, single episode, major, with psychotic symptoms
C0494400|episode; depressive, severe, with psychotic symptoms
C0439020|Complaining of feeling depressed
C0439020|C/O - feeling depressed
C0439020|C/O - feeling depressed (context-dependent category)
C0439020|Complaining of feeling depressed (finding)
C0005587|Bipolar Depression
C0005587|bipolar affective disorder, current episode depressed (diagnosis)
C0005587|bipolar affective disorder, current episode depressed
C0005587|bipolar disorder affective, current episode depressed
C0005587|Bipolar affective disorder, depressed
C0005587|Bipolar affective disorder, current episode depression
C0005587|Manic-depressive - now depressed
C0005587|Bipolar affective disorder, current episode depression (disorder)
C0005587|Depression, Bipolar
C0025193|Melancholia
C0025193|Melancholias
C0025193|Melancholic Depression
C0025193|Depression with Melancholic Features
C0025193|Melancholia, NOS
C0025193|Melancholia NOS
C0282126|Depressions, Neurotic
C0282126|Neurotic Depressions
C0282126|Neurotic depression
C0282126|Depression, Neurotic
C0282126|Depression neurotic
C0282126|depression; neurotic
C0282126|depressive; state, neurotic
C0282126|neurotic; depression
C0282126|state; depressive, neurotic
C0282126|Neurotic depressive state
C0011573|Depressions, Endogenous
C0011573|Endogenous Depressions
C0011573|Endogenous Depression
C0011573|Depression;endogenous
C0011573|Endogenous depression (disorder)
C0011573|depression endogenous
C0011573|Endogenous depression (diagnosis)
C0011573|depression; endogenous
C0011573|endogenous; depression
C0011573|Endogenous depression [Ambiguous]
C0011573|Depression, Endogenous
C0520669|single episode major depression with atypical features (diagnosis)
C0520669|single episode major depression with atypical features
C0520669|Major depressive disorder, single episode with atypical features
C0520669|Major depressive disorder, single episode with atypical features (disorder)
C0154413|Major depressive disorder, recurrent episode, severe degree, specified as with psychotic behavior
C0154413|Recurrent depressive disorder, current episode severe with psychotic symptoms
C0154413|severe recurrent major depression with psychotic features (diagnosis)
C0154413|recurrent major depression with psychotic features (diagnosis)
C0154413|recurrent major depression with psychotic features
C0154413|severe recurrent major depression with psychotic features
C0154413|Major depressive disorder, recurrent episode, severe degree, specified as with psychotic behaviour
C0154413|Rec depr psych-psychotic
C0154413|Major depressive affective disorder, recurrent episode, severe, specified as with psychotic behavior
C0154413|[X]Recurrent severe episodes of psychotic depression
C0154413|[X]Recurrent depressive disorder, current episode severe with psychotic symptoms
C0154413|[X]Recurrent depressive disorder, current episode severe with psychotic symptoms (disorder)
C0154413|[X]Recurrent severe episodes of psychogenic depressive psychosis
C0154413|[X]Recurrent severe episodes of major depression with psychotic symptoms
C0154413|severe recurrent major depression with psychosis
C0154413|severe recurrent major depression with psychosis (diagnosis)
C0154413|major depression recurrent severe with psychosis
C0154413|Severe recurrent major depression with psychotic features (disorder)
C0024517|Major depressive disorder, single episode, unspecified degree
C0024517|single episode major depression (diagnosis)
C0024517|single episode major depression
C0024517|Depress psychosis-unspec
C0024517|Major depressive disorder, single episode, unspecified
C0024517|Major depressive disorder, single episode
C0024517|single episode of major depression
C0024517|Major depressive affective disorder, single episode, unspecified
C0024517|Single major depressive episode
C0024517|Single major depressive episode, unspecified
C0024517|Single major depressive episode NOS (disorder)
C0024517|Single major depressive episode (disorder)
C0024517|Single major depressive episode NOS
C0024517|Single major depressive episode, unspecified (disorder)
C0024517|Major depression, single episode (disorder)
C0024517|Major depression, single episode
C0024517|depressive; episode, major
C0024517|Major depression, single episode, NOS
C0024517|Single Episode of Major Depressive Disorder
C0024517|Major depressive disorder; single episode
C0302874|Depressive personality disorder
C0302874|Personality;depressive
C0302874|Depressive personality
C0302874|depressive; personality disorder
C0302874|personality disorder; depressive
C0154405|Major depressive disorder, single episode, severe degree, without mention of psychotic behavior
C0154405|severe single episode major depression without psychotic features (diagnosis)
C0154405|severe single episode major depression without psychotic features
C0154405|Depress psychosis-severe
C0154405|Major depressive disorder, single episode, severe without psychotic features
C0154405|Major depressv disord, single epsd, sev w/o psych features
C0154405|Major depressive affective disorder, single episode, severe, without mention of psychotic behavior
C0154405|Severe major depression, single episode, without psychotic features
C0154405|Severe major depression, single episode, without psychotic features (disorder)
C0154406|Major depressive disorder, single episode, severe degree, specified as with psychotic behavior
C0154406|Severe major depression, single episode, with psychotic features (disorder)
C0154406|Severe major depression, single episode, with psychotic features
C0154406|Major depressive disorder, single episode, severe with psychotic features
C0154406|severe single episode major depression with psychotic features
C0154406|severe single episode major depression with psychotic features (diagnosis)
C0154406|Depr psychos-sev w psych
C0154406|Major depressv disord, single epsd, severe w psych features
C0154406|Major depressive affective disorder, single episode, severe, specified as with psychotic behavior
C0154409|Major depressive disorder, recurrent episode, unspecified degree
C0154409|recurrent major depression
C0154409|recurrent major depression (diagnosis)
C0154409|Recurr depr psychos-unsp
C0154409|Major depressive disorder, recurrent, unspecified
C0154409|Major depressive disorder, recurrent
C0154409|recurrent episodes of major depression
C0154409|Major depressive affective disorder, recurrent episode, unspecified
C0154409|Recurrent major depressive episode NOS (disorder)
C0154409|Recurrent major depressive episodes, unspecified (disorder)
C0154409|Recurrent major depressive episodes, unspecified
C0154409|Recurrent major depressive episode
C0154409|Recurrent major depressive episode NOS
C0154409|Recurrent major depressive episodes
C0154409|Recurrent major depressive episodes (diagnosis)
C0154409|major depression recurrent episodes
C0154409|Major depressive disorder, recurrent episode
C0154409|Recurrent major depression (disorder)
C0154409|Recurrent major depressive disorder
C0154409|Recurrent major depressive episodes (disorder)
C0154409|Recurrent major depression, NOS
C0154409|Recurrent major depressive disorder, NOS
C0154409|Major depressive disorder; recurrent episode
C0154437|atypical depressive disorder (diagnosis)
C0154437|atypical depressive disorder
C0154437|Atypical depressive dis
C0154437|Atypical depression
C0154437|Atypical depressive disorder (disorder)
C0154437|[X]Atypical depression
C0154437|atypical; depression
C0154437|depression; atypical
C0338893|Major depressive disorder, recurrent episode, in partial or unspecified remission
C0338893|Recur depr psyc-part rem
C0338893|Major depressive affective disorder, recurrent episode, in partial or unspecified remission
C0338893|Recurrent major depressive episodes, in partial or unspecified remission
C0338893|Recurrent major depressive episodes, in partial or unspecified remission (disorder)
C0085159|Affective Disorder, Seasonal
C0085159|Affective Disorders, Seasonal
C0085159|Disorder, Seasonal Affective
C0085159|Disorder, Seasonal Mood
C0085159|Disorders, Seasonal Affective
C0085159|Disorders, Seasonal Mood
C0085159|Mood Disorder, Seasonal
C0085159|Mood Disorders, Seasonal
C0085159|Seasonal Affective Disorder
C0085159|Seasonal Mood Disorders
C0085159|SAD
C0085159|SEASONAL AFFECTIVE DIS
C0085159|seasonal depression
C0085159|depression in a seasonal pattern
C0085159|seasonal depression (symptom)
C0085159|depression seasonal pattern (diagnosis)
C0085159|depression seasonal pattern
C0085159|seasonal pattern depression
C0085159|Seasonal Affective Disorders
C0085159|Seasonal Mood Disorder
C0085159|Seasonal Affective Disorder [Disease/Finding]
C0085159|[X]Seasonal depressive disorder
C0085159|Seasonal affective disorder (disorder)
C0085159|[X] Seasonal depressive disorder
C0085159|[X]SAD - Seasonal affective disorder
C0085159|seasonal affective disorder (diagnosis)
C0085159|SAD - Seasonal affective disorder
C0085159|depression; seasonal
C0085159|seasonal; depression
C0011581|Depressive neurosis
C0011581|Depressive Disorders
C0011581|Depressive Disorder
C0011581|Depressive Neuroses
C0011581|Disorder, Depressive
C0011581|Disorders, Depressive
C0011581|Neuroses, Depressive
C0011581|DEPRESSIVE DIS
C0011581|depression
C0011581|depression (diagnosis)
C0011581|Depressive disorder NOS
C0011581|Depressive Disorder [Disease/Finding]
C0011581|Neurosis, Depressive
C0011581|Mood disorder of depressed type
C0011581|[X]Depressive disorder NOS
C0011581|Mood disorder of depressed type (disorder)
C0011581|Mood disorder with depressive feature
C0011581|-- Depression
C0011581|Depressive illness
C0011581|Depressive disorder (disorder)
C0011581|depression; behavioral disorder
C0011581|depressive; disorder
C0011581|depressive; neurosis
C0011581|disorder; depressive
C0011581|neurosis; depressive
C0011581|Depressive disorder, NOS
C0011581|Disorder;depressive
C0362037|Depression postoperative
C0362037|[D]Postoperative depression
C0362037|Postoperative depression (diagnosis)
C0362037|Postoperative depression
C0362037|Postoperative depression (disorder)
C0362037|Postoperative depression, NOS
C0221745|Depression suicidal
C0221745|Suicidal depression
C0520665|Menopausal depression
C0520665|depression menopausal
C0520665|depression menopausal (diagnosis)
C0520665|Postmenopausal depression
C0520665|Depression postmenopausal
C0520665|Menopausal depression (disorder)
C0520665|depression; menopausal
C0520665|menopausal; depression
C0520665|Menopausal depression, NOS
C0520665|Postmenopausal depression, NOS
C3665457|chronic depressive personality disorder (diagnosis)
C3665457|chronic depressive personality disorder
C3665457|Chronic depressive personality disorder (disorder)
C3665457|Chr depressive person
C3665457|Chronic depressive disorder
C0871610|winter depression
C0871610|depression more in winter (symptom)
C0871610|depression more in winter
C2165514|summer depression
C2165514|depression more in summer (symptom)
C2165514|depression more in summer
C2165515|depression preceded by high activity level
C2165515|depression preceded by high activity level (symptom)
C2165509|depression accompanied by eating more
C2165509|depression accompanied by eating more (symptom)
C2165508|depression accompanied by eating less
C2165508|depression accompanied by eating less (symptom)
C2165511|depression accompanied by sleeping more (symptom)
C2165511|depression accompanied by sleeping more
C2165510|depression accompanied by sleeping less (symptom)
C2165510|depression accompanied by sleeping less
C2165507|depression accompanied by persistent worry (symptom)
C2165507|depression accompanied by persistent worry
C2165518|depression relieved by good news
C2165518|depression relieved by good news (symptom)
C2165519|depression relieved by medication (symptom)
C2165519|depression relieved by medication
C2165517|depression relieved by counseling (symptom)
C2165517|depression relieved by counseling
C2165520|depression seasonal pattern with few nonseasonal occurrences
C2165520|depression seasonal pattern w/ few nonseasonal occurrences
C2165520|depression seasonal pattern with few nonseasonal occurrences (symptom)
C2165520|seasonal depression with few nonseasonal occurrences
C0338908|Mixed anxiety and depressive disorder
C0338908|depression with anxiety
C0338908|depression with anxiety (diagnosis)
C0338908|Anxiety/depression
C0338908|Anxiety with depression
C0338908|Mixed anxiety and depressive disorder (disorder)
C0338908|[X]Mixed anxiety and depressive disorder
C0338908|Anxiety depression
C0338908|Anxious depression
C0338908|Mixed anxiety & depressive
C0338908|depression; anxiety
C0338908|disorder; mixed, anxiety and depressive
C0338908|mixed; disorder, anxiety and depressive
C0338908|anxiety; depression
C2063289|chronic major depression (diagnosis)
C2063289|chronic major depression
C2063866|Resistant Depression, Treatment
C2063866|Treatment-Resistant Depressive Disorders
C2063866|Therapy-Resistant Depressions
C2063866|Depressions, Refractory
C2063866|Therapy Resistant Depression
C2063866|Depression, Refractory
C2063866|Depressive Disorder, Treatment-Resistant
C2063866|Disorders, Treatment-Resistant Depressive
C2063866|Depression, Treatment Resistant
C2063866|Depressions, Treatment Resistant
C2063866|Treatment Resistant Depressions
C2063866|Depressive Disorder, Treatment Resistant
C2063866|Depressive Disorders, Treatment-Resistant
C2063866|Disorder, Treatment-Resistant Depressive
C2063866|Treatment-Resistant Depressive Disorder
C2063866|Depression, Therapy-Resistant
C2063866|Depressions, Therapy-Resistant
C2063866|Resistant Depressions, Treatment
C2063866|Refractory Depressions
C2063866|Refractory Depression
C2063866|Therapy-Resistant Depression
C2063866|Treatment Resistant Depression
C2063866|Depressive Disorder, Treatment-Resistant [Disease/Finding]
C2063866|treatment-refractory depression (diagnosis)
C2063866|treatment-refractory depression
C2938940|Post stroke depression
C3203510|Postictal depression
C0086133|Depressive Syndromes
C0086133|Syndrome, Depressive
C0086133|Syndromes, Depressive
C0086133|Depressive Syndrome
C0349712|[X]Recurrent brief depressive episodes
C0349712|[X] Recurrent brief depressive episodes
C0349712|depression recurrent brief
C0349712|Recurrent brief depressive disorder (diagnosis)
C0349712|Recurrent brief depressive disorder
C0349712|Recurrent brief depressive disorder (disorder)
C0349712|disorder; recurrent brief depressive
C0349712|recurrent brief depressive; disorder
C0270461|Major depressive disorder, in remission (MDD)
C0270461|MDD IN REMISSION
C0270461|MAJOR DEPRESSIVE DISORDER REMISSION
C0270461|Major depression, in remission
C0270461|major depression - in remission
C0270461|major depressive disorder - in remission
C0270461|major depressive disorder, in remission (diagnosis)
C0270461|major depressive disorder, in remission
C0270461|Major depression in remission (disorder)
C0270461|Major depression in remission
C0270461|Major depression in remission, NOS
C0270457|major depression severe without psychotic features
C0270457|severe major depressive disorder without psychotic features (diagnosis)
C0270457|severe major depressive disorder without psychotic features
C0270457|Severe major depression without psychotic features
C0270457|Severe major depression without psychotic features (disorder)
C0270456|major depression moderate
C0270456|Moderate major depression (diagnosis)
C0270456|Moderate major depression
C0270456|Moderate major depression (disorder)
C1282644|Major depression, melancholic type (disorder)
C1282644|Major depression, melancholic type
C1282644|major depression melancholic type
C1282644|Major depression, melancholic type (diagnosis)
C1282644|Major depression, melancholic type (disorder) [Ambiguous]
C0349218|Recurrent depressive disorder
C0349218|Recurrent depressive disorder, unspecified
C0349218|[X]Recurrent depressive disorder, unspecified
C0349218|[X]Recurrent depressive disorder
C0349218|[X] Recurrent episodes of reactive depression
C0349218|[X] Recurrent episodes of depressive reaction
C0349218|[X]Recurrent depressive disorder, unspecified (disorder)
C0349218|[X]Recurrent depressive disorder (disorder)
C0349218|[X]Recurrent episodes of reactive depression
C0349218|[X]Recurrent episodes of depressive reaction
C0349218|[X]Recurrent depressive disorder (finding)
C0701819|recurrent major depression with melancholia
C0701819|recurrent major depression with melancholia (diagnosis)
C0701819|Recurrent major depressive disorder with melancholic features
C0701819|Recurrent major depressive disorder with melancholic features (disorder)
C0012706|Depressive disorder NEC in SNOMEDCT
C0012706|Depressive disorder NEC
C0012706|Depressive disorder NEC (disorder)
C0588006|Mild depression
C0588006|Mild depression (disorder)
C0588006|depression mild
C0588006|Mild depression (diagnosis)
C0588006|Mild depression -RETIRED-
C0338808|Post-schizophrenic depression
C0338808|Post-schizophrenic depression (disorder)
C0338808|Post-schizophrenic depression (diagnosis)
C0338808|depression post-schizophrenic
C0338808|depression; post-schizophrenic
C0338808|post-schizophrenic; depression
C0338808|postpsychotic depression; schizophrenic
C0338808|postschizophrenic depression
C0338808|schizophrenia; postpsychotic depression
C0588007|Moderate depression (disorder)
C0588007|Moderate depression
C0588007|Moderate depression (diagnosis)
C0588007|depression moderate
C0270488|depression stuporous
C0270488|Stuporous depression
C0270488|Stuporous depression (diagnosis)
C0270488|Stuporous depression (disorder)
C0581390|Postviral depression
C0581390|Postviral depression (diagnosis)
C0581390|depression postviral
C0581390|Postviral depression (disorder)
C0588008|Severe depression
C0588008|Severe depression (disorder)
C0588008|Severe depression (diagnosis)
C0588008|depression severe
C0588008|depression; severe
C0588008|severe; depression
C0581391|depression chronic
C0581391|chronic depression
C0581391|chronic depression (symptom)
C0581391|chronic depression (diagnosis)
C0581391|Chronic depression (disorder)
C0520675|Minor depressive disorder (diagnosis)
C0520675|Minor depressive disorder
C0520675|depression minor
C0520675|Minor depressive disorder (disorder)
C0338897|Masked depression
C0338897|Masked depression (disorder)
C0338897|depression masked
C0338897|Masked depression (diagnosis)
C0338897|depression; masked
C0338897|masked; depression
C0221480|depression recurrent
C0221480|recurrent depression
C0221480|recurrent depression (symptom)
C0221480|Recurrent depression (disorder)
C0221480|recurrent depression (diagnosis)
C3697979|Depressive disorder in remission
C3697979|Depressive disorder in remission (disorder)
C3838728|Depressive disorder in mother complicating childbirth (disorder)
C3838728|Depressive disorder in mother complicating childbirth
C3838728|Depression in childbirth
C0520676|premenstrual dysphoric disorder
C0520676|PMDD
C0520676|premenstrual dysphoric disorder (diagnosis)
C0520676|premenstrual disorder
C0520676|Dysphoric Disorder, Premenstrual
C0520676|Syndrome, Premenstrual Dysphoric
C0520676|Disorder, Premenstrual Dysphoric
C0520676|Premenstrual Dysphoric Disorder [Disease/Finding]
C0520676|Premenstrual Dysphoric Syndrome
C0520676|Premenstrual dysphoric disorder (disorder)
C3825465|Depression in infants
C3825452|Depression in old age
C0005586|Bipolar Disorders
C0005586|MANIC DEPRESSIVE ILLNESS
C0005586|Bipolar Affective Psychosis
C0005586|Bipolar Disorder
C0005586|Manic Depressive Psychosis
C0005586|Manic-Depressive Psychoses
C0005586|Psychoses, Bipolar Affective
C0005586|Psychoses, Manic Depressive
C0005586|Psychosis, Bipolar Affective
C0005586|Psychosis, Manic Depressive
C0005586|Bipolar affective disorder
C0005586|Disorder, Bipolar
C0005586|Manic-depressive psychosis
C0005586|Bipolar affective disorder, unspecified
C0005586|BIPOLAR DIS
C0005586|Manic-Depression
C0005586|manic depressive disorder
C0005586|BPAD
C0005586|unspecified bipolar disorder
C0005586|unspecified bipolar disorder (diagnosis)
C0005586|bipolar disorder not otherwise specified
C0005586|Manic depressive
C0005586|Bipolar disorder NOS
C0005586|manic-depressive reaction
C0005586|manic-depressive illness
C0005586|Bipolar disorder, unspecified
C0005586|Affective Psychosis, Bipolar
C0005586|Bipolar Disorder [Disease/Finding]
C0005586|Psychoses, Manic-Depressive
C0005586|Psychosis, Manic-Depressive
C0005586|Disorder;bipolar
C0005586|Depression;manic
C0005586|Psychosis;manic depressive
C0005586|Bi-polar Disorder
C0005586|Bipolar disorder (disorder)
C0005586|Unspecified bipolar affective disorder
C0005586|Depressive-manic psych.
C0005586|Unspecified bipolar affective disorder (disorder)
C0005586|Unspecified bipolar affective disorder, unspecified
C0005586|[X]Bipolar affective disorder, unspecified
C0005586|[X]Bipolar affective disorder, unspecified (disorder)
C0005586|Unspecified bipolar affective disorder, unspecified (disorder)
C0005586|Unspecified bipolar affective disorder, NOS
C0005586|Manic-depress.psychoses
C0005586|Unspecified bipolar affective disorder, NOS (disorder)
C0005586|Manic depression
C0005586|Manic depressive reaction
C0005586|Reaction manic-depressive
C0005586|Psychosis manic-depressive
C0005586|MDI - Manic-depressive illness
C0005586|bipolar; disorder, affective
C0005586|bipolar; disorder
C0005586|disorder; bipolar, affective
C0005586|disorder; bipolar
C0005586|manic-depressive; disorder
C0005586|manic-depressive; psychosis
C0005586|manic-depressive; syndrome
C0005586|psychosis; manic-depressive
C0005586|syndrome; manic-depressive
C0005586|Bipolar disorder, NOS
C0005586|Bipolar Mood Disorder
C0005586|Manic-depressive reaction NOS
C0005586|Manic-depressive syndrome NOS
C4065471|disruptive mood dysregulation disorder (diagnosis)
C4065471|depression disruptive mood dysregulation disorder
C4065471|disruptive mood dysregulation disorder
C1386135|Acute depression
C1386135|Acute depression (disorder)
C1386135|depression; acute
C1386135|acute; depression
C4074822|Depressive disorder in mother complicating pregnancy
C4074822|Depressive disorder in mother complicating pregnancy (disorder)
C1282921|Cotard's syndrome
C1282921|Cotard syndrome
C1282921|Cotard syndrome (disorder)
C1282921|Cotard's syndrome (diagnosis)
C1282921|Cotard's syndrome (disorder)
C1282921|Cotard
C0011580|reactive psychotic depression
C0011580|reactive depressive psychosis
C0011580|reactive depressive psychosis (diagnosis)
C0011580|depressive type psychosis (mdd) reactive
C0011580|Psychotic reactive depression
C0011580|Reactive depressive psychosis (disorder)
C0011580|depression; reactive, psychotic
C0011580|depressive; reaction, psychotic
C0011580|psychosis; depressive, reactive
C0011580|psychosis; reactive, depressive
C0011580|reaction; depressive, psychotic
C0011580|reactive; depression, psychotic
C0011580|Psychotic Depressive Reaction
C0011580|Depression, Reactive, Psychotic
C0270497|Schizoaffective disorder, depressive type
C0270497|Schizoaffective disorder depressive type
C0270497|Schizophreniform psychosis, depressive type
C0270497|Schizoaffective disorder, depressive type (disorder)
C0270497|disorder; schizoaffective, depressive type
C0270497|psychosis; schizophreniform, depressive type
C0339017|Depressive conduct disorder
C0339017|Depressive conduct disorder (disorder)
C0339017|depressive conduct disorder (diagnosis)
C0339017|behavioral disorder; depressive
C0339017|depressive; behavioral disorder
C0349216|Other depressive episodes
C0349216|[X]Other depressive episodes (disorder)
C0349216|[X]Other depressive episodes
C0556016|[X]Single episode agitated depression without psychotic symptoms
C0556016|[X] Single episode agitated depression without psychotic symptoms (disorder)
C0556016|[X] Single episode agitated depression without psychotic symptoms
C0556018|[X] Manic-depressive psychosis, depressed type without psychotic symptoms
C0556018|[X]Manic-depressive psychosis, depressed type without psychotic symptoms
C0556018|[X] Manic-depressive psychosis, depressed type without psychotic symptoms (disorder)
C0556018|psychosis; manic-depressive, depressed type (without psychotic symptoms)
C0556017|[X]Single episode vital depression without psychotic symptoms
C0556017|[X] Single episode major depression without psychotic symptoms
C0556017|[X]Single episode major depression without psychotic symptoms
C0556017|[X] Single episode major depression without psychotic symptoms (disorder)
C0436599|On examination - depressed
C0436599|O/E - depressed
C0436599|O/E - depressed (finding)
C0436599|On examination - depressed (context-dependent category)
C0436599|On examination - depressed (disorder)
C0338715|Drug-induced depressive state
C0338715|Drug-induced organic affective syndrome
C0338715|Drug-induced depressive state (disorder)
C0338715|Depressive state induced by drugs
C0338715|Drug-induced depression
C2712011|Decreased Depressed Mood
C1579931|Depressed - symptom
C1579931|depression (symptom)
C1579931|depression
C1579931|Miserable
C3874774|Depressed mood with postpartum onset (finding)
C3874774|Depressed mood with postpartum onset
C3874774|Depressed mood in postpartum period
C3874774|Depressed Mood During Post Partum Period
C3698286|Depressed mood in Alzheimer disease
C3698286|Depressed mood in Alzheimer's disease (disorder)
C3698286|Alzheimers dementia with depressed mood
C3698286|Depressed mood in Alzheimer's disease
C2165504|depressed, but unlike previous grieving for a death or loss
C2165504|depressed, but unlike previous grieving for a death or loss (physical finding)
C3836786|mood depressed postpartum (physical finding)
C3836786|mood depressed postpartum
C0150041|Hopelessness
C0150041|feelings of hopelessness (symptom)
C0150041|feelings of hopelessness
C0150041|Feeling of Hopelessness
C0150041|Hopeless
C0150041|rndx hopelessness (diagnosis)
C0150041|rndx hopelessness
C0150041|Feeling;hopeless
C0150041|Loss of hope for the future
C0150041|Feeling of hopelessness (finding)
C0150041|Loss of hope for the future (finding)
C0150041|Feels there is no future
C0150041|No hope for the future
C0150041|Negative about the future
C0150041|Cannot see a future
C0150041|Feeling hopeless
C0150041|Feeling hopeless (finding)
C2219873|feels pessimistic about future or brooding about past
C2219873|feels pessimistic about future or brooding about past (symptom)
C2219873|feel pessimistic about future, or brooding about past
C2219873|pessimistic about the future, or brooding about the past
C2165505|depression 1-3 days prior to menstruation
C2165505|depression 1-3 days prior to menstruation (symptom)
C2165506|depression accompanied by (symptom)
C2165506|depression accompanied by
C2165506|depression accompanied
C2165516|depression is relieved
C2165516|factors relieving depression
C2165516|factors relieving depression (symptom)
C2051715|depression occurring
C2051715|pattern of depression (symptom)
C2051715|pattern of depression
C2169543|depression recently
C2169543|recent depression
C2169543|recent depression (symptom)
C1561368|CTCAE Grade 3 Depression
C1561368|Grade 3 Depression
C1561366|CTCAE Grade 1 Depression
C1561366|Grade 1 Depression
C1561367|CTCAE Grade 2 Depression
C1561367|Grade 2 Depression
C1561369|CTCAE Grade 4 Depression
C1561369|Grade 4 Depression
C1561370|CTCAE Grade 5 Depression
C1561370|Grade 5 Depression
