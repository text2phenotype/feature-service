C3160090|HCV NS3/4A Protease Inhibitors [MoA]
C2605855|simeprevir
C3696072|simeprevir sodium
C3696747|simeprevir Pill
C3696511|simeprevir 150 MG [Olysio]
C3696563|simeprevir Oral Capsule [Olysio]
C3696697|simeprevir 150 MG
C3696720|simeprevir Oral Capsule
C3696748|simeprevir Oral Product
C3695381|simeprevir 150 MG Oral Capsule [Olysio]
C3695403|simeprevir 150 MG Oral Capsule
C1738934|boceprevir
C3209784|boceprevir Pill
C3655064|Boceprevir:Susc:Pt:Isolate:OrdQn:Genotyping
C3154647|boceprevir 200 MG
C3154648|boceprevir Oral Capsule
C3154649|boceprevir 200 MG Oral Capsule
C3154651|boceprevir 200 MG [Victrelis]
C3154652|boceprevir Oral Capsule [Victrelis]
C3209783|boceprevir Oral Product
C3655750| Isolate
C3154653|boceprevir 200 MG Oral Capsule [Victrelis]
C1876229|telaprevir
C3215243|telaprevir Pill
C3655063|Telaprevir:Susc:Pt:Isolate:OrdQn:Genotyping
C3154700|telaprevir 375 MG
C3154702|telaprevir 375 MG [Incivek]
C3154710|telaprevir Oral Tablet
C3154711|telaprevir 375 MG Oral Tablet
C3154712|telaprevir Oral Tablet [Incivek]
C3215242|telaprevir Oral Product
C3655696|Telaprevir Isolate
C3154713|telaprevir 375 MG Oral Tablet [Incivek]
C0717864|Ribavirin+interferon alpha-2b
C0789390|Ribavirin 200 MG Oral Tablet
C0789393|Ribavirin 40 MG/ML Oral Solution
C0979999|Ribavirin 20 MG/ML Inhalant Solution
C1128545|Ribavirin 200 MG
C1131183|Ribavirin 40 MG/ML
C0035525|Ribavirin
C0073221|ribavirin amidine
C0571293|Tribavirin allergy
C0627880|tributylribavirin
C0935908|palivizumab/ribavirin
C1875630|PEGINTERFERON/RIBAVIRIN
C3189667|Ribavirin Powder
C3219702|Ribavirin Pill
C3547186|response to ribavirin
C0979998|Ribavirin 200 MG Oral Capsule
C0361571|Ribavirin 100 MG Oral Capsule
C0413496|Tribavirin adverse reaction
C0717864|Ribavirin+interferon alpha-2b
C0789390|Ribavirin 200 MG Oral Tablet
C0789393|Ribavirin 40 MG/ML Oral Solution
C0979999|Ribavirin 20 MG/ML Inhalant Solution
C1128545|Ribavirin 200 MG
C1131183|Ribavirin 40 MG/ML
C1140523|Ribavirin 20 MG/ML
C1186936|Ribavirin 100 MG
C1240752|Ribavirin Oral Capsule [Rebetol]
C1242547|Ribavirin Oral Tablet [Copegus]
C1247842|Ribavirin Oral Capsule
C1247843|Ribavirin Oral Solution
C1247844|Ribavirin Oral Tablet
C1253016|Ribavirin Inhalant Solution
C1382829|Ribavirin 400 MG
C1454123|5-nor carbocyclic ribavirin
C1589272|Ribavirin Oral Solution [Rebetol]
C1593466|Ribavirin 200 MG [Rebetol]
C1593727|Ribavirin 200 MG [Copegus]
C1601182|Ribavirin 200 MG [Ribasphere]
C1601183|Ribavirin Oral Capsule [Ribasphere]
C1621221|Ribavirin Inhalant Solution [Virazole]
C1626919|Ribavirin 400 MG Oral Tablet
C1641488|Ribavirin:MCnc:Pt:Ser/Plas:Qn
C1676705|Ribavirin 600 MG Oral Tablet
C1677789|Ribavirin 600 MG
C1694682|Ribavirin Oral Tablet [RibaTab]
C1702720|Ribavirin 400 MG [Ribasphere]
C1703270|Ribavirin 600 MG [Ribasphere]
C1704170|Ribavirin Oral Tablet [Ribasphere]
C1878904|Ribavirin 400 MG [RibaTab]
C1589271|Ribavirin 40 MG/ML [Rebetol]
C1616510|Ribavirin 20 MG/ML [Virazole]
C0021747|Interferons
C0733470|human leukocyte interferon
C3652465|Interferon
C3653501|DIRECT ACTING ANTIVIRALS
C3541967|Thiosemicarbazones, direct acting antivirals
C3653501|DIRECT ACTING ANTIVIRALS
C3540755|Protease inhibitors, direct acting antivirals
C3541969|Neuraminidase inhibitors, direct acting antivirals
C3653443|Cyclic amines, direct acting antivirals
C3653392|Phosphonic acid derivatives, direct acting antivirals
C0330845|Astragalus Plant
C1095897|Astragalus preparation
C3864824|paritaprevir
C3864824|paritaprevir
C3883274|paritaprevir dihydrate
C3864967|ombitasvir / paritaprevir / Ritonavir
C3865150|paritaprevir 75 MG
C3865210|ombitasvir / paritaprevir / Ritonavir Pill
C3882783|dasabuvir / ombitasvir / paritaprevir / Ritonavir
C4075296|Paritaprevir in oral dosage form
C4276327|paritaprevir 50 MG
C4298645|Paritaprevir:Susc:Pt:Isolate:Ord:Genotyping
C3865188|ombitasvir / paritaprevir / Ritonavir Oral Tablet
C3865211|ombitasvir / paritaprevir / Ritonavir Oral Product
C4276383|dasabuvir / ombitasvir / paritaprevir / Ritonavir Pill
C3864964|{2 (dasabuvir 250 MG Oral Tablet) / 2 (ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet) } Pack
C3871501|Dasabuvir;Ombitasvir, Paritaprevir, Ritonavir Oral tablet
C3871617|Dasabuvir;Ombitasvir/Paritaprevir/Ritonavir NA Oral Tablet
C3882779|dasabuvir/ombitasvir/paritaprevir/ritonavir oral kit
C4047040|ombitasvir / paritaprevir / Ritonavir Oral Tablet [Technivie]
C4276384|dasabuvir / ombitasvir / paritaprevir / Ritonavir Oral Product
C3854281|{2 (dasabuvir 250 MG Oral Tablet) / 2 (ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet) } Pack [Viekira Pak]
C3865125|ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet
C4046961|ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG [Technivie]
C4276118|dasabuvir 200 MG / ombitasvir 8.33 MG / paritaprevir 50 MG / Ritonavir 33.33 MG Extended Release Oral Tablet (3) 24HR Pack
C4276368|dasabuvir / ombitasvir / paritaprevir / Ritonavir Extended Release Oral Tablet
C4046169|ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet [Technivie]
C4275375|24 HR dasabuvir 200 MG / ombitasvir 8.33 MG / paritaprevir 50 MG / Ritonavir 33.33 MG Extended Release Oral Tablet
C3696409|Olysio
C3696630|Olysio Pill
C3695381|simeprevir 150 MG Oral Capsule [Olysio]
C3696511|simeprevir 150 MG [Olysio]
C3696563|simeprevir Oral Capsule [Olysio]
C3696631|Olysio Oral Product
C4080053|grazoprevir
C4080453|elbasvir / grazoprevir
C4255551|Grazoprevir anhydrous
C4080449|grazoprevir 100 MG
C4080450|elbasvir / grazoprevir Oral Product
C4080451|elbasvir / grazoprevir Pill
C4080452|elbasvir / grazoprevir Oral Tablet
C4298643|Grazoprevir:Susc:Pt:Isolate:Ord:Genotyping
C4307658|elbasvir-grazoprevir drug combination
C4080454|elbasvir 50 MG / grazoprevir 100 MG Oral Tablet
C4080457|elbasvir / grazoprevir Oral Tablet [Zepatier]
C4080456|elbasvir 50 MG / grazoprevir 100 MG [Zepatier]
C4080460|elbasvir 50 MG / grazoprevir 100 MG Oral Tablet [Zepatier]
C3854280|Viekira Pak
C2976303|sofosbuvir
C3857383|ledipasvir
C3858025|Harvoni
C3858199|Harvoni Pill
C3858200|Harvoni Oral Product
C3852670|ombitasvir
C3854280|Viekira Pak  
C4080455|Zepatier
C4080052|elbasvir
C4299883|Elbasvir
C4080453|elbasvir grazoprevir
C4080453|grazoprevir  
C3252090|daclatasvir
C3892852|daclatasvir dihydrochloride
C4047229|daclatasvir Pill
C4298749|Daclatasvir
C4299898|Daclatasvir  
C3851350|ledipasvir
C3858051|ledipasvir / sofosbuvir
C3858262|ledipasvir 90 MG
C3858300|ledipasvir / sofosbuvir Oral Tablet
C3858321|ledipasvir / sofosbuvir Pill
C3858322|ledipasvir / sofosbuvir Oral Product
C4075037|Ledipasvir in oral dosage form
C4298751|Ledipasvir:Susc:Pt:Isolate:Ord:Genotyping
C4299632| Isolate
C3858080|ledipasvir 90 MG / sofosbuvir 400 MG Oral Tablet
C3858162|ledipasvir / sofosbuvir Oral Tablet [Harvoni]
C3858113|ledipasvir 90 MG / sofosbuvir 400 MG [Harvoni]
C3857383|ledipasvir 90 MG / sofosbuvir 400 MG Oral Tablet [Harvoni]  
C2605856|435350, TMC
C2605856|TMC435350
C2605856|TMC-435350
C2605856|TMC 435350
C2745868|435, TMC
C2745868|TMC435
C2745868|TMC-435
C2745868|TMC 435
C3696409|Olysio
C2605855|simeprevir
C2605855|simeprevir (medication)
C2605855|antiviral simeprevir
C2605855|Simeprevir (substance)
C2605855|N-(17-(2-(4-isopropylthiazole-2-yl)-7-methoxy-8-methylquinolin-4-yloxy)-13-methyl-2,14-dioxo-3,13-diazatricyclo(13.3.0.04,6)octadec-7-ene-4-carbonyl)(cyclopropyl)sulfonamide
C2605855|Simeprevir [Chemical/Ingredient]
C2605855|Simeprevir (product)
C3696072|simeprevir sodium
C3696072|simeprevir (as sodium)
C3696748|simeprevir Oral Product
C3696748|Oral form simeprevir (product)
C3696748|Oral form simeprevir
C4075528|Simeprevir + sofosbuvir (product)
C4075528|Simeprevir + sofosbuvir
C3696720|simeprevir Oral Capsule
C3696630|Olysio Pill
C3695403|Simeprevir 150 MG Oral Capsule
C3695403|Simeprevir 150mg Oral capsule
C3695403|Simeprevir Sodium Cap 150 MG (Base Equivalent)
C3695403|SIMEPREVIR 150MG CAP
C3695403|SIMEPREVIR 150MG CAP [VA Product]
C3695381|simeprevir 150 MG Oral Capsule [Olysio]
C3695381|Olysio 150 MG Oral Capsule
C3695381|OLYSIO 150mg Capsule
C3695381|simeprevir 150 MG (as simeprevir sodium 154.4 mg ) Oral Capsule [Olysio]
C3695381|Olysio, 150 mg oral capsule
C3696511|simeprevir 150 MG [Olysio]
C3696563|simeprevir Oral Capsule [Olysio]
C3696631|Olysio Oral Product
C3154650|Victrelis
C3154650|vicrtelis
C1738934|N-(3-amino-1-(cyclobutylmethyl)-2,3-dioxopropyl)-3-(2-((((1,1-dimethylethyl)amino)carbonyl)amino)-3,3-dimethyl-1-oxobutyl)-6,6-dimethyl-3-azabicyclo(3.1.0)hexan-2-carboxamide
C1738934|boceprevir
C1738934|antivirals boceprevir
C1738934|antivirals boceprevir (medication)
C1738934|Boceprevir (substance)
C1738934|Boceprevir (product)
C1738934|3-Azabicyclo(3.1.0)hexane-2-carboxamide, N-(3-amino-1-(cyclobutylmethyl)-2,3-dioxopropyl)-3-((2S)-2-((((1,1- dimethylethyl)amino)carbonyl)amino)-3,3-dimethyl-1-oxobutyl)-6,6- dimethyl-, (1R,2S,5S)-
C3154649|Boceprevir Cap 200 MG
C3154649|BOCEPREVIR 200MG CAP
C3154649|boceprevir 200 mg oral capsule
C3154649|BOCEPREVIR 200MG CAP [VA Product]
C3154649|Boceprevir 200mg Oral capsule
C3154649|Boceprevir 200mg capsule (product)
C3154649|Boceprevir 200mg capsule
C1741239|Sch-503034
C1741239|Sch 503034
C1741239|Sch503034
C3896865|EBP 520
C3240332|Victrelis Pill
C3154648|boceprevir Oral Capsule
C3655064|Boceprevir:Susc:Pt:Isolate:OrdQn:Genotyping
C3655064|Boceprevir [Susceptibility] by Genotype method
C3655064|Boceprevir Islt Genotyp
C3655064|Boceprevir:Susceptibility:Point in time:Isolate:Quantitative or Ordinal:Genotyping
C3154651|boceprevir 200 MG [Victrelis]
C3154652|boceprevir Oral Capsule [Victrelis]
C3154653|BOCEPREVIR 200 mg ORAL CAPSULE [VICTRELIS]
C3154653|Victrelis 200 MG Oral Capsule
C3154653|VICTRELIS 200mg Capsule
C3154653|Victrelis, 200 mg oral capsule
C3240331|Victrelis Oral Product
C3154701|Incivek
C1876229|telaprevir
C1876229|antiviral telaprevir
C1876229|antiviral telaprevir (medication)
C1876229|Telaprevir (substance)
C1876229|Telaprevir (product)
C3281323|VRT-111950
C3281324|MP-424
C3281325|LY-570310
C1956374|VX-950
C1956374|VX 950
C1956374|VX950 cpd
C3154711|telaprevir 375 MG Oral Tablet
C3154711|Telaprevir Tab 375 MG
C3154711|TELAPREVIR 375MG TAB
C3154711|TELAPREVIR 375MG TAB,28 [VA Product]
C3154711|TELAPREVIR 375MG TAB,28
C3154711|TELAPREVIR 375MG TAB [VA Product]
C3154711|Telaprevir 375mg Oral tablet
C3154711|TELAPREVIR 375MG TAB,UD
C3154711|TELAPREVIR 375MG UD TAB
C3154711|TELAPREVIR 375MG TAB,UD [VA Product]
C3154711|Telaprevir 375mg tablet
C3154711|Telaprevir 375mg tablet (product)
C3226078|Incivek Pill
C3154710|telaprevir Oral Tablet
C3655063|Telaprevir Islt Genotyp
C3655063|Telaprevir [Susceptibility] by Genotype method
C3655063|Telaprevir:Susc:Pt:Isolate:OrdQn:Genotyping
C3655063|Telaprevir:Susceptibility:Point in time:Isolate:Quantitative or Ordinal:Genotyping
C3154702|telaprevir 375 MG [Incivek]
C3154712|telaprevir Oral Tablet [Incivek]
C3154713|telaprevir 375 MG Oral Tablet [Incivek]
C3154713|Incivek 375 MG Oral Tablet
C3154713|INCIVEK 375mg Tablet
C3154713|Incivek, 375 mg oral tablet
C3154713|INCIVEK 375 MG Oral Tablet, Twice Daily
C3226077|Incivek Oral Product
C0979954|Rebetron, single dose 1000 mg/day oral and injectable kit
C0979954|REBETRON 1000/PAK 3 PKT (1241-02)
C0979954|Rebetron Combination Package for Patients < = 75 KG, Intron A 6,000,000 UNT/ML Single Dose Vials / 70 Rebetol Capsules
C0979954|REBETRON 1000/PAK 3 PKT (1241-02) [VA Product]
C0979954|{6 (0.5 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution [Intron A]) / 70 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Patients < = 75 KG, Intron A 6,000,000 UNT/ML Single Dose Vials / 70 Rebetol Capsules]
C0979953|Rebetron Combination Package for Patients < = 75 KG, Intron A 6,000,000 UNT/ML Multi-Dose Vial / 70 Rebetol Capsules
C0979953|REBETRON 1000/MDV PKT (1236-02)
C0979953|REBETRON 1000/MDV PKT (1236-02) [VA Product]
C0979953|{1 (3 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution [Intron A]) / 70 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Patients < = 75 KG, Intron A 6,000,000 UNT/ML Multi-Dose Vial / 70 Rebetol Capsules]
C0979955|REBETRON 1000/PEN PKT (1258-02)
C0979955|Rebetron Combination Package for Patients < = 75 KG, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 70 Rebetol Capsules
C0979955|REBETRON 1000/PEN PKT (1258-02) [VA Product]
C0979955|{1 (1.2 ML) (Interferon Alfa-2b 15000000 UNT/ML Injectable Solution [Intron A]) / 70 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Patients < = 75 KG, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 70 Rebetol Capsules]
C0979955|Interferon Alfa-2b;Ribavirin 3MILLION IU/0.2ML-200MG Multiple Routes Kit [REBETRON 1000]
C0979957|Rebetron, single dose 1200 mg/day oral and injectable kit
C0979957|Rebetron Combination Package for Patients > = 75 KG, Intron A 6,000,000 UNT/ML Single Dose Vials / 84 Rebetol Capsules
C0979957|REBETRON 1200/PAK 3 PKT (1241-01)
C0979957|REBETRON 1200/PAK 3 PKT (1241-01) [VA Product]
C0979957|{6 (0.5 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution [Intron A]) / 84 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Patients > = 75 KG, Intron A 6,000,000 UNT/ML Single Dose Vials / 84 Rebetol Capsules]
C2342666|REBETRON 1200/PEN PKT (1258-01)
C2342666|Rebetron Combination Package for Patients > = 75 KG, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 84 Rebetol Capsules
C2342666|{1 (1.2 ML Interferon Alfa-2b 15000000 UNT/ML Injectable Solution [Intron A]) / 84 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Patients > = 75 KG, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 84 Rebetol Capsules]
C2342666|REBETRON 1200/PEN PKT (1258-01) [VA Product]
C2342666|{1 (1.2 ML) (Interferon Alfa-2b 15000000 UNT/ML Injectable Solution [Intron A]) / 84 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Patients > = 75 KG, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 84 Rebetol Capsules]
C2342666|Interferon Alfa-2b;Ribavirin 3MILLION IU/0.2ML-200MG Multiple Routes Kit [REBETRON 1200]
C0979959|Rebetron, multiple dose 600 mg/day oral and injectable kit
C0979959|Rebetron Combination Package for Rebetol Dose Reduction, Intron A 6,000,000 UNT/ML Multi-Dose Vial / 42 Rebetol Capsules
C0979959|REBETRON 600/MDV PKT (1236-03)
C0979959|REBETRON 600/MDV PKT (1236-03) [VA Product]
C0979959|{1 (3 ML Interferon Alfa-2b 6000000 UNT/ML Injectable Solution [Intron A]) / 42 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Rebetol Dose Reduction, Intron A 6,000,000 UNT/ML Multi-Dose Vial / 42 Rebetol Capsules]
C0979959|{1 (3 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution [Intron A]) / 42 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Rebetol Dose Reduction, Intron A 6,000,000 UNT/ML Multi-Dose Vial / 42 Rebetol Capsules]
C0979959|Interferon Alfa-2b;Ribavirin 3MILLION IU/0.2ML-200MG Multiple Routes Kit [REBETRON 600]
C2342670|Rebetron Combination Package for Rebetol Dose Reduction, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 42 Rebetol Capsules
C2342670|REBETRON 600/PEN PKT (1258-03)
C2342670|REBETRON 600/PEN PKT (1258-03) [VA Product]
C2342670|{1 (1.2 ML Interferon Alfa-2b 15000000 UNT/ML Injectable Solution [Intron A]) / 42 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Rebetol Dose Reduction, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 42 Rebetol Capsules]
C2342670|{1 (1.2 ML) (Interferon Alfa-2b 15000000 UNT/ML Injectable Solution [Intron A]) / 42 (Ribavirin 200 MG Oral Capsule [Rebetol]) } Pack [Rebetron Combination Package for Rebetol Dose Reduction, Intron A 15,000,000 UNT/ML Multi-Dose Pen / 42 Rebetol Capsules]
C1444872|Ribavirin 200mg capsule+interferon alpha-2b 3million iu/vial injection solution (product)
C1444872|Ribavirin 200mg capsule+interferon alpha-2b 3million iu/vial injection solution
C0705810|interferon alfa-2b-ribavirin single dose 1000 mg/day oral and injectable kit
C0705812|interferon alfa-2b-ribavirin single dose 600 mg/day oral and injectable kit
C0705811|interferon alfa-2b-ribavirin single dose 1200 mg/day oral and injectable kit
C0789390|Ribavirin 200 MG Oral Tablet
C0789390|Ribavirin 200mg Oral tablet
C0789390|RIBAVIRIN 200MG TAB
C0789390|Ribavirin Tab 200 MG
C0789390|RIBAVIRIN 200 mg ORAL TABLET, FILM COATED
C0789390|RIBAVIRIN 200MG TAB [VA Product]
C0789390|RIBAVIRIN 200 mg ORAL TABLET, FILM COATED [Ribavirin]
C0789390|Ribavirin 200mg tablet (product)
C0789390|Ribavirin 200mg tablet
C0789390|Ribavirin, 200 mg oral tablet
C3473212|Ribavirin 200mg Oral tablet, Ribavirin 400mg Oral tablet
C3473212|RIBASPHERE RibaPak KIT
C3473212|Ribavirin Tab 200 MG & Ribavirin Tab 400 MG Dose Pack
C3473212|{7 (Ribavirin 200 MG Oral Tablet) / 7 (Ribavirin 400 MG Oral Tablet) } Pack
C3473212|RibaPak 600, 200 mg-400 mg oral tablet
C3473212|RIBAVIRIN 200MGX7/400MGX7 TAB DOSEPK 14
C3473212|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14 [VA Product]
C3473212|RIBAVIRIN 200MG X 7/400MG X 7 TAB DOSEPACK,14
C3473212|ribavirin 200 MG (7) Oral Tablet / ribavirin 400 MG (7) Oral Tablet Pack
C3473212|Ribavirin;Ribavirin 200 MG; 400 MG Oral Tablet [RIBASPHERE RIBAPAK]
C3473212|Ribasphere RibaPak 600mg/day Dose Pack Tablet
C3700547|RIBAVIRIN 200 mg ORAL TABLET, FILM COATED [Moderiba]
C3700547|Moderiba 200 MG Oral Tablet
C3700547|Ribavirin 200 MG Oral Tablet [Moderiba]
C3700547|Moderiba, 200 mg oral tablet
C3700547|Moderiba 200mg Tablet
C1169961|Copegus 200 MG Oral Tablet
C1169961|Ribavirin 200 MG Oral Tablet [Copegus]
C1169961|Copegus 200mg Tablet
C1169961|Ribavirin 200 mg ORAL TABLET, FILM COATED [Copegus]
C1169961|Copegus, 200 mg oral tablet
C1694693|Ribasphere, 200 mg oral tablet
C1694693|Ribasphere 200 MG Oral Tablet
C1694693|Ribavirin 200 MG Oral Tablet [Ribasphere]
C1694693|RIBAVIRIN 200 mg ORAL TABLET, FILM COATED [RIBASPHERE]
C1694693|Ribasphere 200mg Tablet
C0789393|Ribavirin 40 MG/ML Oral Solution
C0789393|Ribavirin Soln 40 MG/ML
C0789393|RIBAVIRIN 200MG/5ML SOLN,ORAL
C0789393|RIBAVIRIN 200MG/5ML ORAL SOLN
C0789393|RIBAVIRIN 200MG/5ML SOLN,ORAL [VA Product]
C0789393|Ribavirin 40mg Oral solution
C0789393|Ribavirin 40mg/mL oral solution (product)
C0789393|Ribavirin 40mg/mL oral solution
C1586219|Rebetol 40 MG/ML Oral Solution
C1586219|Ribavirin 40 MG/ML Oral Solution [Rebetol]
C1586219|Rebetol 40mg/ml Solution
C1586219|ribavirin 40 mg in 1 mL ORAL LIQUID [REBETOL]
C1586219|Rebetol, 40 mg/mL oral solution
C0350923|Ribavirin 20 MG/ML Inhalant Solution [Virazid]
C0350923|Virazid 20 MG/ML Inhalant Solution
C0979999|Ribavirin 20 MG/ML Inhalant Solution
C0979999|RIBAVIRIN 6GM/VI INHL SOLN
C0979999|RIBAVIRIN 6GM/VIL INHL [VA Product]
C0979999|RIBAVIRIN 6GM/VIL INHL
C0979999|Ribavirin 6g Powder for nebulizer solution
C0979999|Ribavirin 6 GM Inhalation Powder for Solution
C0979999|Ribavirin 6g/vial powder (product)
C0979999|Ribavirin 6g/vial powder
C0979999|ribavirin 6 GM Powder for Inhalant Solution
C0979999|Ribavirin For Inhal Soln 6 GM
C0979999|Tribavirin 6g inhalation (pdr for recon)
C0979999|Tribavirin 6g inhalation (pdr for recon) (product)
C0979999|Tribavirin 6g inhalation (pdr for recon) (substance)
C0979999|ribavirin 6 g inhalation powder for reconstitution
C0708742|Ribavirin 20 MG/ML Inhalant Solution [Virazole]
C0708742|Virazole 20 MG/ML Inhalant Solution
C0708742|Virazole 6g Powder for Inhalation Solution
C0708742|Ribavirin 6 GM Inhalation Powder for Solution [VIRAZOLE]
C0708742|Ribavirin 6 g RESPIRATORY (INHALATION) POWDER, FOR SOLUTION [Virazole]
C0708742|Virazole, 6 g inhalation powder for reconstitution
C3701057|Ribavirin 200 MG [Moderiba]
C1601182|Ribavirin 200 MG [Ribasphere]
C1593466|Ribavirin 200 MG [Rebetol]
C1593727|Ribavirin 200 MG [Copegus]
C1589271|Ribavirin 40 MG/ML [Rebetol]
C1622085|Virazole
C1622085|Vilona
C1622085|ICN Brand of Ribavirin
C0702025|ICN-1229
C0702025|ICN 1229
C0702025|ICN1229
C0702024|Ribamide
C0702024|Ribamidyl
C0702024|Ribamidil
C0035525|Ribavirin
C0035525|1H-1,2,4-Triazole-3-carboxamide, 1-beta-D-ribofuranosyl-
C0035525|1-Beta-D-ribofuranosyl-1,2,4-triazolo-3-carboxamide
C0035525|1-Beta-D-ribofuranosyl-1H-1,2,4-triazole-3-carboxamide
C0035525|RTCA
C0035525|RIBA
C0035525|ribavirin (medication)
C0035525|Tribavirin
C0035525|Ribavirin [Chemical/Ingredient]
C0035525|Ribovirin
C0035525|Tribavirin (product)
C0035525|1-.beta.-D-Ribofuranosyl-1H-1,2, 4-triazole-3-carboxamide
C0035525|Ribavirin (product)
C0035525|Ribavirin (substance)
C2317046|Respiratory form ribavirin
C2317046|Respiratory form ribavirin (product)
C2315948|Oral form ribavirin (product)
C2315948|Oral form ribavirin
C2148525|ribavirin 200mg capsules given with interferon alfa-2b (medication)
C2148525|ribavirin 200mg capsules given with interferon alfa-2b
C1626919|ribavirin 400 mg oral tablet
C1626919|Ribavirin Tab 400 MG
C1626919|Ribavirin 400mg Oral tablet
C1626919|RIBAVIRIN 400MG TAB
C1626919|Ribavirin, 400 mg oral tablet
C1626919|RIBAVIRIN 400MG TAB [VA Product]
C1626919|RIBAVIRIN 400 mg ORAL TABLET, FILM COATED
C1626919|Ribavirin 400mg tablet (product)
C1626919|Ribavirin 400mg tablet
C1676705|ribavirin 600 mg oral tablet
C1676705|Ribavirin Tab 600 MG
C1676705|Ribavirin 600mg tablet (product)
C1676705|Ribavirin 600mg tablet
C1676705|Ribavirin, 600 mg oral tablet
C1676705|Ribavirin 600mg Oral tablet
C1676705|RIBAVIRIN 600MG TAB
C1676705|RIBAVIRIN 600MG TAB [VA Product]
C1676705|RIBAVIRIN 600 mg ORAL TABLET, FILM COATED
C1170183|Copegus
C1870873|2-(3-amino-3-deoxyxylofuranosyl)thiazole-4-carboxamide
C3700973|Moderiba
C0637676|methyl 1-ribofuranosyl-1,2,4-triazole-3-carboxamidate
C0637676|MRTC
C0627880|TB-ribavirin
C0627880|tributylribavirin
C0640066|3-ribofuranosyl-1,2,4-triazole-5-carboxamide
C0076656|2-ribofuranosylthiazole-4-carboxamide
C0076656|riboxamide
C0076656|tiazofurin
C0076656|TCAR
C0639452|1-(5'-O-sulfamoyl-beta-D-ribofuranosyl)(1,2,4)triazole-3-carbonitrile
C0639452|SRTCN
C1454123|5'-nor carbocyclic ribavirin
C0073218|ribavirin 5'-diphosphate
C0073218|ribavirin-DP
C0637674|ethyl 1-ribofuranosyl-1,2,4-triazole-3-carboximidate
C0637674|ERTC
C0764977|4-fluoro-1-ribofuranosyl-1H-pyrazole-3-carboxamide
C0764977|4-FRPC
C0605624|1-(4-thio-beta-D-ribofuranosyl)-1,2,4-triazole-3-carboxamide
C0632093|5'-O-beta-D-glucopyranosyl ribavirin
C0632093|5'-O-glucopyranosyl ribavirin
C0647853|2-(2',3'-dideoxyglyceropent-2-enofuranosyl)thiazole-4-carboxamide
C0647853|2',3'-didehydro-2',3'-dideoxytiazofurin
C0640069|2-ribofuranosyl-1,2,3-triazole-4,5-dicarboxamide
C1957632|tiazofurin monophosphate
C0632095|5'-O-beta-D-galactopyranosyl ribavirin
C0632095|5'-O-galactopyranosyl ribavirin
C0073219|1H-1,2,4-Triazole-3-carboxamide, 1-(5-O-(aminosulfonyl)-beta-D-ribofuranosyl)-
C0073219|5'-O-sulfamoyl-1-ribofuranosyl-1,2,4-triazole-3-carboxamide
C0073219|ribavirin 5'-sulfamate
C0073219|1-(5'-O-sulfamoyl-beta-ribofuranosyl)-(1,2,4)triazole-3-carboxamide
C0140479|ribavirin 2',3',5'-triacetate
C0073221|1-beta-D-ribofuranosyl-1,2,4-triazole-3-carboxamidine
C0073221|ribamidine
C0073221|ribavirin amidine
C0073221|TCNR
C0073221|Taribavirin
C0073221|viramidine
C0639450|1-(5'-O-sulfamoyl-beta-ribofuranosyl)(1,2,4)triazole-3-thiocarboxamide
C0639450|SRTC
C0647851|2-(2',3'-dideoxyglyceropentafuranosyl)thiazole-4-carboxamide
C0647851|2',3'-dideoxytiazofurin
C0050823|adenylyl-(3'-5')-virazole
C0050823|adenylyl-(3'-5')ribavirin
C0050823|3'-Adenylic acid, 3'-5'-ester with 1-beta-D-ribofuranosyl-1H-1,2,4-triazole-3-carboxamide
C2240463|{7 (Ribavirin 400 MG Oral Tablet) / 7 (Ribavirin 600 MG Oral Tablet) } Pack
C2240463|Ribavirin 400mg Oral tablet, Ribavirin 600mg Oral tablet
C2240463|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14 [VA Product]
C2240463|RIBAVIRIN 600MG X 7/400MG X 7 TAB DOSEPACK,14
C2240463|RIBAVIRIN 600MGX7/400MGX7 TAB DOSEPK 14
C4075513|Ribavirin Injectable Product
C4075513|Parenteral form ribavirin (product)
C4075513|Parenteral form ribavirin
C0361571|Ribavirin 100 MG Oral Capsule
C0361571|Ribavirin 100mg capsule
C0361571|Ribavirin 100mg capsule (product)
C0361571|Ribavirin 100mg capsule (substance)
C0979998|Ribavirin 200 MG Oral Capsule
C0979998|Ribavirin 200mg Oral capsule
C0979998|RIBAVIRIN 200MG CAP
C0979998|Ribavirin Cap 200 MG
C0979998|RIBAVIRIN 200MG CAP [VA Product]
C0979998|RIBAVIRIN 200 mg ORAL CAPSULE [Ribavirin]
C0979998|Ribavirin 200mg capsule
C0979998|Ribavirin 200mg capsule (product)
C0979998|Ribavirin 200mg capsule (substance)
C0979998|Ribavirin, 200 mg oral capsule
C0717864|INTERFERON ALFA-2B/RIBAVIRIN
C0717864|interferon alfa-2b-ribavirin
C0717864|Ribavirin+interferon alpha-2b (product)
C0717864|Ribavirin+interferon alpha-2b
C0702029|Viramide
C0731013|Virazid
C1170576|Rebetol
C1170576|Ribavirin Merck Brand
C1170576|Merck Brand of Ribavirin
C1170576|Pfizer Brand of Ribavirin
C1170576|Essex Brand of Ribavirin
C1564036|Grossman Brand of Ribavirin
C1564036|Virazide
C1564036|Dermatech Brand of Ribavirin
C1564336|Ribasphere
C1564336|Three Rivers Pharmaceuticals Brand of Ribavirin
C0722990|Rebetron
C1878903|RibaTab
C0935908|palivizumab/ribavirin
C0935908|PALI/RIBA
C1339084|Ribavirin 400 MG Oral Capsule
C2341626|Ribavirin 500mg Oral tablet
C2341626|Ribavirin 500 MG Oral Tablet
C2341626|RIBAVIRIN 500 mg ORAL TABLET, FILM COATED
C2341626|Ribavirin, 500 mg oral tablet
C3222959|Copegus Pill
C3232238|Rebetol Pill
C3237959|RibaTab Pill
C3237961|Ribasphere Pill
C1247842|Ribavirin Oral Capsule
C1247844|Ribavirin Oral Tablet
C3701173|Moderiba Pill
C1169620|Rebetol 200 MG Oral Capsule
C1169620|Ribavirin 200 MG Oral Capsule [Rebetol]
C1169620|Rebetol 200mg Capsule
C1169620|Rebetol, 200 mg oral capsule
C1584733|Ribasphere 200 MG Oral Capsule
C1584733|Ribavirin 200 MG Oral Capsule [Ribasphere]
C1584733|Ribasphere 200mg Capsule
C1584733|Ribasphere, 200 mg oral capsule
C2342580|{6 (0.5 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution) / 70 (Ribavirin 200 MG Oral Capsule) } Pack
C2342658|{1 (3 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution) / 70 (Ribavirin 200 MG Oral Capsule) } Pack
C2342661|{1 (1.2 ML) (Interferon Alfa-2b 15000000 UNT/ML Injectable Solution) / 70 (Ribavirin 200 MG Oral Capsule) } Pack
C2342663|{1 (3 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution) / 84 (Ribavirin 200 MG Oral Capsule) } Pack
C2342664|{6 (0.5 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution) / 84 (Ribavirin 200 MG Oral Capsule) } Pack
C2342665|{1 (1.2 ML) (Interferon Alfa-2b 15000000 UNT/ML Injectable Solution) / 84 (Ribavirin 200 MG Oral Capsule) } Pack
C2342667|{1 (3 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution) / 42 (Ribavirin 200 MG Oral Capsule) } Pack
C2342668|{6 (0.5 ML) (Interferon Alfa-2b 6000000 UNT/ML Injectable Solution) / 42 (Ribavirin 200 MG Oral Capsule) } Pack
C2342669|{1 (1.2 ML) (Interferon Alfa-2b 15000000 UNT/ML Injectable Solution) / 42 (Ribavirin 200 MG Oral Capsule) } Pack
C0413496|Adverse reaction to tribavirin
C0413496|Adverse reaction to tribavirin (finding)
C0413496|Tribavirin adverse reaction
C0413496|Tribavirin adverse reaction (disorder)
C0413496|Ribavirin adverse reaction
C1595591|Ribavirin 20 MG/ML [Virazid]
C1616510|Ribavirin 20 MG/ML [Virazole]
C1240752|Ribavirin Oral Capsule [Rebetol]
C1601183|Ribavirin Oral Capsule [Ribasphere]
C0789392|Ribavirin 20 MG/ML Oral Solution
C1589272|Ribavirin Oral Solution [Rebetol]
C3701110|Ribavirin Oral Tablet [Moderiba]
C1242547|Ribavirin Oral Tablet [Copegus]
C1704170|Ribavirin Oral Tablet [Ribasphere]
C1694682|Ribavirin Oral Tablet [RibaTab]
C1621221|Ribavirin Inhalant Solution [Virazole]
C1235816|Ribavirin Inhalant Solution [Virazid]
C3701058|Ribavirin 400 MG [Moderiba]
C1702720|Ribavirin 400 MG [Ribasphere]
C1878904|Ribavirin 400 MG [RibaTab]
C3668937|Moderiba 400 MG Oral Tablet
C3668937|Ribavirin 400 MG Oral Tablet [Moderiba]
C3668937|RIBAVIRIN 400 mg ORAL TABLET, FILM COATED [Moderiba]
C1694134|Ribasphere, 400 mg oral tablet
C1694134|Ribasphere 400 MG Oral Tablet
C1694134|Ribavirin 400 MG Oral Tablet [Ribasphere]
C1694134|RIBAVIRIN 400 mg ORAL TABLET, FILM COATED [RIBASPHERE]
C1694134|Ribasphere 400mg Tablet
C1878399|RibaTab 400mg Tablet
C1878399|Ribavirin 400 MG Oral Tablet [RibaTab]
C1878399|RibaTab 400 MG Oral Tablet
C1878399|RibaTab, 400 mg oral tablet
C2240739|{14 (Ribavirin 400 MG Oral Tablet) } Pack
C2240739|RIBAVIRIN 400MG TAB DOSEPACK 14
C2240739|RIBAVIRIN 400MG TAB DOSEPACK,14 [VA Product]
C2240739|RIBAVIRIN 400MG TAB DOSEPACK,14
C1641488|Ribavirin:MCnc:Pt:Ser/Plas:Qn
C1641488|Ribavirin [Mass/volume] in Serum or Plasma
C1641488|Ribavirin SerPl-mCnc
C1641488|Ribavirin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C3668939|Ribavirin 600 MG Oral Tablet [Moderiba]
C3668939|Moderiba 600 MG Oral Tablet
C3668939|RIBAVIRIN 600 mg ORAL TABLET, FILM COATED [Moderiba]
C1694694|Ribasphere, 600 mg oral tablet
C1694694|Ribasphere 600 MG Oral Tablet
C1694694|Ribavirin 600 MG Oral Tablet [Ribasphere]
C1694694|RIBAVIRIN 600 mg ORAL TABLET, FILM COATED [RIBASPHERE]
C1694694|Ribasphere 600mg Tablet
C1878400|Ribavirin 600 MG Oral Tablet [RibaTab]
C1878400|RibaTab 600mg Tablet
C1878400|RibaTab 600 MG Oral Tablet
C2240738|{14 (Ribavirin 600 MG Oral Tablet) } Pack
C2240738|Ribavirin 600 MG Oral Tablet 7 Day Pack
C2240738|RIBAVIRIN 600MG X 14 TAB DOSEPACK 14
C2240738|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14 [VA Product]
C2240738|RIBAVIRIN 600MG X 14 TAB DOSEPACK,14
C2240738|Ribavirin 600 MG Oral Tablet 14 Count 7 Day Pack
C3701056|Ribavirin 600 MG [Moderiba]
C1703270|Ribavirin 600 MG [Ribasphere]
C1878905|Ribavirin 600 MG [RibaTab]
C0002199|alpha Interferon
C0002199|Interferon alpha
C0002199|Interferon-alpha
C0002199|Leukocyte Interferon
C0002199|Lymphoblast Interferon
C0002199|Lymphoblastoid Interferon
C0002199|interferon alfa
C0002199|alpha-interferon
C0002199|Interferon, Leukocyte
C0002199|Interferon, Lymphoblastoid
C0002199|Interferon, alpha
C0002199|Interferon, Lymphoblast
C0002199|Interferon-alpha [Chemical/Ingredient]
C0002199|Interferon.alpha
C0002199|IFNa
C0002199|Interferon alfa (substance)
C0002199|Interferon alfa (product)
C0002199|Alpha interferon (substance)
C0002199|interferon A
C0002199|IFN-A
C0021745|Immune Interferon
C0021745|Interferon, Type II
C0021745|interferon gamma
C0021745|Interferon gamma (human lymphocyte protein moiety reduced)
C0021745|Interferon Type II
C0021745|Interferon gamma (substance)
C0021745|gamma interferon
C0021745|gamma-interferon
C0021745|Interferon-gamma
C0021745|Interferon, Immune
C0021745|Interferon, gamma
C0021745|Interferon-gamma [Chemical/Ingredient]
C0021745|Type II Interferon
C0021745|Interferon.gamma
C0021745|IFNg
C0021745|Gamma interferon (substance)
C0021745|Interferon gamma (product)
C0021745|IFN-G
C0021745|lFN-Gamma
C0015980|beta Interferon
C0015980|Fibroblast Interferon
C0015980|Interferon beta
C0015980|Interferon-beta
C0015980|Interferon beta (substance)
C0015980|Interferon, Fibroblast
C0015980|Interferon, beta
C0015980|Interferon-beta [Chemical/Ingredient]
C0015980|beta-Interferon
C0015980|Interferon.beta
C0015980|IFNb
C0015980|Interferon beta (product)
C0015980|Beta interferon (substance)
C0015980|IFN-B
C0015980|Endogenous Interferon Beta
C0015980|IFN-Beta
C0015980|Interferon Beta, Natural
C0015980|Natural human interferon beta
C2352835|locteron
C0021743|Interferon Type I
C0021743|Interferon, Type I
C0021743|Interferons, Type I
C0021743|Interferons Type I
C0021743|Type I Interferons
C0021743|Interferon Type I [Chemical/Ingredient]
C0021743|Type I Interferon
C0021747|Interferons
C0021747|interferon
C0021747|interferons (medication)
C0021747|Interferons [Chemical/Ingredient]
C0021747|IFN
C0021747|Interferons (product)
C0021747|Interferon (substance)
C2743274|IFNphi1 protein, zebrafish
C2743274|interferon phi1, zebrafish
C2743275|inteferon phi2, zebrafish
C2743275|IFNphi2 protein, zebrafish
C0164613|IFN-alpha Con 1
C0164613|consensus IFN-alpha
C0164613|rIFN-con-1
C0164613|recombinant consensus interferon alpha
C0164613|interferon-alpha Con(1)
C0164613|interferon alfacon-1
C0164613|methionyl-interferon-consensus
C0164613|methionyl interferon consensus
C0164613|interferon consensus, methionyl
C0164613|Recombinant methionyl human consensus interferon
C0164613|IFN Alfacon-1
C0164613|Recombinant Consensus Interferon
C0164613|r-metHuIFN-Con1
C0164613|CIFN
C0164613|Interferon alfacon-1 agent
C0164613|CIFN (interferon)
C0164613|interferon alfacon-1 (medication)
C0164613|interferon alfacon-1 [Chemical/Ingredient]
C0164613|Interferon alfacon-1 agent (substance)
C0164613|Interferon alfacon-1 preparation
C0164613|consensus interferon
C0164613|Interferon alfacon-1 preparation (substance)
C0021741|Interferon gamma-1b
C0021741|Interferon gamma-1b preparation
C0021741|interferon gamma-2a
C0021741|interferon gamma-1b [Chemical/Ingredient]
C0021741|Recombinant Interferon Gamma-1b
C0021741|N(Sup 2)-L-Methionyl-1-139-Interferon G
C0021741|interferon gamma-1b (medication)
C0021741|Interferon gamma-1b (substance)
C0021741|Interferon gamma-1b preparation (product)
C0021741|Interferon gamma-1b preparation (substance)
C0021734|Interferon Alfa-2a
C0021734|recombinant interferon alpha-2a
C0021734|Recombinant Interferon Alfa-2a
C0021734|Alpha 2 Interferon
C0021734|IFN alpha-2A
C0021734|rHuIFN-a 2a
C0021734|IFN-Alpha 2
C0021734|Interferon alfa 2a
C0021734|Interferon Alfa
C0021734|Interferon alpha-2a preparation
C0021734|INTERFERON ALFA-2A,RECOMBINANT
C0021734|interferon alfa-2a [Chemical/Ingredient]
C0021734|interferon alfa-2a (medication)
C0021734|Interferon alpha-2a (substance)
C0021734|Interferon alpha-2a preparation (product)
C0021734|Interferon alpha-2a
C0021734|Interferon alpha-2a preparation (substance)
C0021735|Interferon Alfa-2b
C0021735|IFN alpha-2B
C0021735|recombinant interferon alfa-2b
C0021735|interferon alpha-2b
C0021735|Interferon alpha-2b preparation
C0021735|INTERFERON ALFA 2-B
C0021735|INTERFERON ALFA-2B,RECOMBINANT
C0021735|recombinant interferon alpha-2b
C0021735|interferon alfa-2b [Chemical/Ingredient]
C0021735|Interferon alpha-2b, recombinant
C0021735|IFNalpha-2b, recombinant
C0021735|interferon alfa-2b (medication)
C0021735|Interferon alpha-2b (substance)
C0021735|Interferon alpha-2b preparation (product)
C0021735|Interferon alpha-2b preparation (substance)
C0021735|Interferon alfa 2b
C0982233|INTERFERON ALFA-3N,HUMAN LEUKOCYTE DERIVED
C0982234|interferon beta-1a
C0982234|interferon beta-1a (medication)
C0982234|INTERFERON BETA-1A,RECOMBINANT
C0982234|Recombinant interferon beta-1a
C0796545|peginterferon alfa-2b
C0796545|PEG interferon alfa-2b
C0796545|pegylated interferon alfa-2b
C0796545|PEG-IFN-a 2b
C0796545|PEG-IFNA2b
C0796545|PEG-Interferon Alfa-2b
C0796545|PEG-IFNalpha-2b
C0796545|PEG-IFN alfa-2b
C0796545|pegylated interferon alpha-2b
C0796545|PEG INF alpha-2b
C0796545|PEG-interferon alpha-2b
C0796545|peginterferon alpha-2b
C0796545|polyethylene glycol-interferon alfa-2b
C0796545|peginterferon alfa-2b [Chemical/Ingredient]
C0796545|polyethylene glycol-interferon alpha-2b
C0796545|PEG INF alfa-2b
C0796545|PEG-IFN alpha-2b
C0796545|Peginterferon alfa-2b (substance)
C0796545|PEG-Intron
C0796545|peginterferon alfa-2b (medication)
C0796545|Peginterferon alfa-2b (product)
C0796545|polyethylene glycol interferon alfa-2b
C0796545|polyethylene glycol IFN-A2b
C0391001|PEG-IFN alfa-2A
C0391001|PEG-IFN alpha-2A
C0391001|PEG-interferon alfa-2A
C0391001|peginterferon alfa-2a
C0391001|Peginterferon alpha-2a (substance)
C0391001|Peginterferon alpha-2a
C0391001|pegylated interferon alfa-2a
C0391001|polyethylene glycol-interferon alfa-2a
C0391001|PEG-interferon alpha-2a
C0391001|pegylated interferon alpha-2a
C0391001|polyethylene glycol-interferon alpha-2a
C0391001|peginterferon alfa-2a [Chemical/Ingredient]
C0391001|peginterferon alfa-2a (medication)
C0391001|Peginterferon alfa-2a (product)
C0391001|PEG-IFNA2a
C3161968|antiviral alpha interferons
C3161968|antiviral alpha interferons (medication)
C0301340|Injectable interferon (substance)
C0301340|Injectable interferon
C0301340|Injectable interferon (product)
C2969476|Interferon drug &#x7C; patient
C1990798|Interferon &#x7C; bld-ser-plas
C1990803|Interferon omega &#x7C; bld-ser-plas
C3657894|INF-epsilon
C3657894|interferon-epsilon, mouse
C4077145|IFN-lambda3, mouse
C4077145|interferon-lambda3, mouse
C0733469|human fibroblast interferon
C0733470|Human Leukocyte Interferon
C0733470|Human Lymphoblastoid Interferon
C0733470|Human Fibroblast Interferon
C0733470|Interferon
C0733470|IFN
C0063697|interferon eicosapeptide
C0063697|interferon eicosapeptide (human lymphoblastoid)
C0063697|ITF-ECP
C0063697|L-Glutamine, L-seryl-L-alpha-aspartyl-L-leucyl-L-prolyl-L-glutaminyl-L-threonyl-L-histidyl-L-seryl-L-leucylglycyl-L-asparaginyl-L-arginyl-L-arginyl-L-alanyl-L-leucyl-L-isoleucyl-L-leucyl-L-leucyl-L-alanyl-
C0965287|(2-sulfo-9-fluorenylmethoxycarbonyl)7-interferon-alpha2
C0965287|hepta-FMS-interferon-alpha2
C1522537|recombinant interferon
C1522537|Human lymphoblastoid interferon
C1522537|Interferons
C1522537|IFN
C1522537|Human Leukocyte Interferon
C1621234|Interferon Alfa-n3
C1621234|INTERFERON ALFA-3N
C1621234|Interferon alpha-n3 agent
C1621234|Interferon alfa-n3 agent
C1621234|interferon alfa-n3 (medication)
C1621234|Interferon alpha-n3 agent (substance)
C1621234|Interferon alpha-n3 preparation
C1621234|Interferon alpha-n3 preparation (substance)
C1621234|Alfa-N3 Interferon
C0876233|Interferon alfa-n1 lymphoblastoid
C0876233|interferon alfa-n1, lymphoblastoid
C0876233|Interferon alfa-n1 lymphoblastoid (substance)
C2000620|IFN-epsilon, human
C2000620|interferon-epsilon, human
C1610033|Ginterferon
C1610033|Human leukocyte interferon
C1610033|alpha interferon
C1610033|leukocyte interferon
C1610033|G-interferon
C1610033|IFN Alpha
C1610033|Interferon Alfa-N3
C1610033|Interferon Alpha
C1610033|alfa-n3 interferon
C1610033|lymphoblast interferon
C1610033|lymphoblastoid interferon
C1610033|Interferon Alpha, Human
C0083028|interferon omega 1
C0083028|interferon omega1
C0083028|interferon omega
C0083028|Interferon.omega
C0083028|Interferon Omega-1
C0083028|IFNW1 protein, human
C0083028|IFN-Alpha-Like
C0083028|IFN-Omega 1
C0083028|IFNW1 Protein
C0083028|IFNW1
C0083028|Interferon Alpha-II-1
C0949830|Astragalus gummifer
C0949830|Astragalus gummifers
C0949830|gummifer, Astragalus
C0949830|gummifers, Astragalus
C0949830|Astragalus gummifer Labill.
C0330845|Astragalus
C0330845|Astragalus Plants
C0330845|Plant, Astragalus
C0330845|Plants, Astragalus
C0330845|Astragalus Plant
C0330845|Astragalus L., 1753
C0330845|Astragalus (Plants)
C0330845|Astragalus species
C0330845|Astragalus species (organism)
C0330845|Locoweeds
C0330845|Astragalus (organism)
C0330845|Astragalus, NOS
C0330845|Locoweeds, NOS
C0949831|membranaceus, Astragalus
C0949831|Astragalus membranaceus
C0949831|Astragalus membranaceus Moench
C1135771|Locoweeds, Wooly
C1135771|Wooly Locoweeds
C1135771|Wooly Locoweed
C1135771|Locoweed, Wooly
C0949829|Milk Vetch
C0949829|MILKVETCH
C0949829|Milk Vetchs
C0949829|Vetchs, Milk
C0949829|Vetch, Milk
C2613731|Astragalus acantherioceras
C2613731|Astragalus acantherioceras Rech.f. & Koie
C2613732|Astragalus aegobromus
C2613732|Astragalus aegobromus Boiss. & Hohen.
C2613733|Astragalus alyssoides
C2613733|Astragalus alyssoides Lam.
C2613734|Astragalus anacamptus
C2613734|Astragalus anacamptus Bunge
C2613735|Astragalus annularis
C2613735|Astragalus annularis Forssk.
C2613736|Astragalus arpilobus
C2613736|Astragalus arpilobus Kar. & Kir.
C2613737|Astragalus asciocalyx
C2613737|Astragalus asciocalyx Bunge
C2613738|Astragalus bakaliensis
C2613738|Astragalus bakaliensis Bunge
C2613739|Astragalus basineri
C2613739|Astragalus basineri Trautv.
C2613740|Astragalus biserrula
C2613740|Astragalus biserrula Bunge
C2613741|Astragalus bombycinus
C2613741|Astragalus bombycinus Boiss.
C2613742|Astragalus brachycalyx
C2613742|Astragalus brachycalyx Fisch. ex Boiss.
C2613743|Astragalus brachypetalus
C2613743|Astragalus brachypetalus Trautv.
C2613744|Astragalus camptoceras
C2613744|Astragalus camptoceras Bunge
C2613745|Astragalus campylanthus
C2613745|Astragalus campylanthus Boiss.
C2613746|Astragalus campylorrhynchus
C2613746|Astragalus campylorhynchus Fisch. & C.A.Mey.
C2613747|Astragalus campylosema
C2613747|Astragalus campylosema Boiss.
C2613748|Astragalus cancellatus
C2613748|Astragalus cancellatus Bunge
C2613749|Astragalus capito
C2613749|Astragalus capito Boiss. & Hohen.
C2613750|Astragalus caraganae
C2613750|Astragalus caraganae Fisch. & C.A.Mey.
C2613751|Astragalus caspicus
C2613751|Astracantha caspica (M.Bieb.) Podlech
C2613751|Astragalus caspicus M.Bieb.
C2613752|Astragalus cephalanthus
C2613752|Astragalus cephalanthus DC.
C2613753|Astragalus chiwensis
C2613753|Astragalus chivensis
C2613753|Astragalus chiwensis Bunge
C2613754|Astragalus chrysostachys
C2613754|Astragalus chrysostachys Boiss.
C2613755|Astragalus citrinus
C2613755|Astragalus citrinus Bunge
C2613756|Astragalus coelicolor
C2613756|Astragalus coelicolor Sirj. & Rech.f.
C2613757|Astragalus commixtus
C2613757|Astragalus commixtus Bunge
C2613758|Astragalus coronilla
C2613758|Astragalus coronilla Bunge
C2613759|Astragalus crenatus
C2613759|Astragalus crenatus Schult.
C2613760|Astragalus curviflorus
C2613760|Astragalus curviflorus Boiss.
C2613761|Astragalus curvipes
C2613761|Astragalus curvipes Trautv.
C2613762|Astragalus dactylocarpus
C2613762|Astragalus dactylocarpus Boiss.
C2613763|Astragalus daenensis
C2613763|Astragalus daenensis Boiss.
C2613764|Astragalus deickianus
C2613764|Astragalus deickianus Bornm.
C2613765|Astragalus dictyolobus
C2613765|Astragalus dictyolobus C.A.Mey. ex Bung
C2613766|Astragalus dieterlei
C2613766|Astragalus dieterlei Podl.
C2613767|Astragalus dipelta
C2613767|Astragalus dipelta Bunge
C2613768|Astragalus dolichophyllus
C2613768|Astragalus dolichophyllus Pall.
C2613769|Astragalus duplostrigosus
C2613769|Astragalus duplostrigosus Post & Beauverd
C2613770|Astragalus eremophilus
C2613770|Astragalus eremophilus Boiss.
C2613771|Astragalus eriostomus
C2613772|Astragalus fasciculifolius
C2613772|Astragalus fasciculifolius Boiss.
C2613773|Astragalus filicaulis
C2613773|Astragalus filicaulis Kar. & Kir.
C2613774|Astragalus fragrans
C2613774|Astragalus fragrans Willd.
C2613775|Astragalus gigantirostratus
C2613775|Astragalus gigantirostratus Maassoumi, Ghahr. & Ghahrem.
C2613776|Astragalus glaucacanthos
C2613776|Astragalus glaucacanthos Fischer & Mey.
C2613777|Astragalus grammocalyx
C2613777|Astragalus grammocalyx Boiss. & Hohen.
C2613778|Astragalus guttatus
C2613778|Astragalus guttatus Banks & Sol.
C2613779|Astragalus hemsleyi
C2613779|Astragalus hemsleyi Aitch. & Baker ex Aitch.
C2613780|Astragalus heterodoxus
C2613780|Astragalus heterodoxus Bunge
C2613781|Astragalus holopsilus
C2613781|Astragalus holopsilus Bunge
C2613782|Astragalus horridus
C2613782|Astragalus horridus Boiss.
C2613783|Astragalus hystrix
C2613783|Astragalus hystrix Fisch. & C.A.Mey.
C2613784|Astragalus jesdianus
C2613784|Astragalus jesdianus Boiss. & Buhse
C2613785|Astragalus jessenii
C2613785|Astragalus jessenii Bunge
C2613786|Astragalus khoshjailensis
C2613786|Astragalus khoshjailensis Sirj. & Rech.f.
C2613787|Astragalus kirrindicus
C2613787|Astragalus kirrindicus Boiss.
C2613788|Astragalus lagopoides
C2613788|Astragalus lagopodioides Vahl
C2613789|Astragalus lamprocarpus
C2613789|Astragalus lamprocarpus Maassoumi
C2613790|Astragalus latifolius
C2613790|Astragalus latifolius Lam.
C2613791|Astragalus ledinghamii
C2613791|Astragalus ledinghamii Barneby
C2613792|Astragalus macrobotrys
C2613792|Astragalus macrobotrys Bunge
C2613793|Astragalus macrosemius
C2613793|Astragalus macrosemius Boiss. & Hohen.
C2613794|Astragalus macrostachys
C2613794|Astragalus macrostachys DC.
C2613795|Astragalus magistratus
C2613795|Astragalus magistratus Maassoumi, Ghahr. & Mozaff.
C2613796|Astragalus masanderanus
C2613796|Astragalus masanderanus Bunge
C2613797|Astragalus migpo
C2613797|Astragalus migpo Kamelin
C2613798|Astragalus mucronifolius
C2613798|Astragalus mucronifolius Boiss.
C2613799|Astragalus multijugus
C2613799|Astragalus multijugus DC.
C2613800|Astragalus murinus
C2613800|Astragalus murinus Boiss.
C2613801|Astragalus nephtonensis
C2613802|Astragalus obtusifolius
C2613803|Astragalus ochreatus
C2613804|Astragalus odoratus
C2613805|Astragalus oleifolius
C2613806|Astragalus ophiocarpus
C2613807|Astragalus ornithopodioides
C2613808|Astragalus oxyglottis
C2613809|Astragalus paradoxus
C2613810|Astragalus peltatus
C2613811|Astragalus perpexus
C2613812|Astragalus persepolitanus
C2613813|Astragalus piptocephalus
C2613814|Astragalus pishchakensis
C2613815|Astragalus pseudorhacodes
C2613816|Astragalus retamocarpus
C2613816|Astragalus retamocarpus Boiss. & Hohen. ex Boiss.
C2613817|Astragalus rhodosemius
C2613817|Astragalus rhodosemius Boiss. & Hausskn.
C2613818|Astragalus robustus
C2613818|Astragalus robustus Bunge
C2613819|Astragalus sahendi
C2613819|Astragalus sahendi Buhse
C2613820|Astragalus scaberrimus
C2613820|stragalus scaberrimus Bunge
C2613821|Astragalus schistocalyx
C2613821|Astragalus schistocalyx Bunge
C2613822|Astragalus schmalhausenii
C2613822|Astragalus schmalhauseni Bunge
C2613823|Astragalus sesamoides
C2613823|Astragalus sesamoides Boiss.
C2613824|Astragalus shelkovnikovii
C2613824|Astragalus shelkovnikovii Grossh.
C2613825|Astragalus siliquosus
C2613825|Astragalus siliquosus Boiss.
C2613826|Astragalus squarrosus
C2613826|Astragalus squarrosus Bunge
C2613827|Astragalus stenolepis
C2613827|Astragalus stenolepis Fisch.
C2613828|Astragalus stocksii
C2613828|Astragalus stocksii Benth. ex Bunge
C2613829|Astragalus straussii
C2613829|Astragalus straussii Hausskn. ex Bornm.
C2613830|Astragalus submitis
C2613830|Astragalus submitis Boiss. & Hohen.
C2613831|Astragalus subsecundus
C2613831|Astragalus subsecundus Boiss. & Hohen.
C2613832|Astragalus tawilicus
C2613832|Astragalus tawilicus C.C.Towns.
C2613833|Astragalus teheranicus
C2613833|Astragalus teheranicus Boiss. & Hohen.
C2613834|Astragalus trachyacanthos
C2613834|Astragalus trachyacanthos Fisch.
C2613835|Astragalus tricholobus
C2613835|Astragalus tricholobus DC.
C2613836|Astragalus urmiensis
C2613836|Astragalus urmiensis Bunge
C2613837|Astragalus vereskensis
C2613837|Astragalus vereskensis Maassoumi & Podlech
C2613838|Astragalus verus
C2613838|Astragalus verus Olivier
C2613839|Astragalus vicarius
C2613839|Astragalus vicarius Lipsky
C2613840|Astragalus vulcanicus
C2613840|Astragalus vulcanicus Bornm.
C2613841|Astragalus xiphidioides
C2613841|Astragalus xiphidioides Freyn & Sint.
C2613842|Astragalus zerdanus
C2613842|Astragalus zerdanus Boiss.
C2613621|Astragalus anserinaefolius
C2613621|Astragalus anserinifolius
C2613621|Astragalus anserinifolius Boiss.
C2613622|Astragalus askius
C2613622|Astragalus askius Bunge
C2613623|Astragalus atricapillus
C2613623|Astragalus atricapillus Bornm.
C2613624|Astragalus austriacus
C2613624|Astragalus austriacus Jacq.
C2613625|Astragalus botryophorus
C2613625|Astragalus botryophorus Maassoumi & Podlech
C2613626|Astragalus brevidens Rydb.
C2613626|Astragalus brevidens
C2613627|Astragalus callistachys Buhse
C2613627|Astragalus callistachys
C2613628|Astragalus campylotrichus
C2613628|Astragalus campylotrichus Bunge
C2613629|Astragalus catacamptus
C2613629|Astragalus catacamptus Bunge
C2613630|Astragalus chartostegius
C2613630|Astragalus chartostegius Boiss. & Hausskn.
C2613631|Astragalus coluteocarpus
C2613631|Astragalus coluteocarpus Boiss.
C2613632|Astragalus compactus Lam.
C2613632|Astragalus compactus
C2613632|Astracantha compacta (Lam.) Podlech
C2613632|Astracantha compacta
C2613633|Astragalus cyclophyllon
C2613633|Astragalus cyclophyllon G.Beck ex Stapf
C2613633|Astragalus cyclophyllon Beck ex Stapf
C2613634|Astragalus depressus
C2613634|Astragalus depressus L.
C2613635|Astragalus echidna
C2613635|Astragalus echidna Bunge
C2613636|Astragalus eriosphaerus
C2613636|Astragalus eriosphaerus Boiss. & Hausskn.
C2613637|Astragalus floccosus
C2613637|Astragalus floccosus Boiss.
C2613638|Astragalus frigidus
C2613638|Astragalus frigidus (L.) A.Gray
C2613639|Astragalus glaux
C2613639|Astragalus glaux L.
C2613640|Astragalus glochideus
C2613640|Astragalus stevenianus subsp. glochideus
C2613640|Astragalus glochideus Boriss.
C2613640|Astragalus stevenianus subsp. glochideus Scischk. ex Sobolevsk.
C2613641|Astragalus glumaceus
C2613641|Astragalus glumaceus Boiss.
C2613642|Astragalus gossypinus
C2613642|Astragalus gossypinus Fisch.
C2613643|Astragalus hololeios
C2613643|Astragalus hololeios Bornm.
C2613644|Astragalus hymenostegis
C2613644|Astragalus hymenostegis Fisch. & C.A.Mey.
C2613645|Astragalus icmadophilus
C2613645|Astragalus icmadophilus Hand.-Mazz.
C2613646|Astragalus kahiricus
C2613646|Astragalus kahiricus DC.
C2613647|Astragalus kerkukiensis
C2613647|Astragalus kerkukiensis Bornm.
C2613648|Astragalus kohrudicus
C2613648|Astragalus kohrudicus Bunge
C2613649|Astragalus koschukensis
C2613649|Astragalus koschukensis Boiss.
C2613650|Astragalus krauseanus
C2613650|Astragalus krauseanus Regel
C2613651|Astragalus laristanicus
C2613651|Astragalus laristanicus Bornm. & Gauba
C2613652|Astragalus leiophyllus
C2613652|Astragalus leiophyllus Freyn & Bornm.
C2613653|Astragalus leptynticus A.A.Maassoumi
C2613653|Astragalus leptynticus
C2613653|Astragalus leptynticus Maassoumi
C2613654|Astragalus leucocephalus
C2613654|Astragalus leucocephalus Graham ex Benth.
C2613655|Astragalus lilacinus
C2613655|Astragalus lilacinus Boiss.
C2613656|Astragalus macrourus
C2613656|Astragalus macrourus Fischer & C.A.Mey.
C2613656|Astragalus macrourus Fisch. & C.A.Mey.
C2613657|Astragalus meyeri
C2613657|Astragalus meyeri Boiss.
C2613658|Astragalus neurophyllus Franch.
C2613658|Astragalus neurophyllus
C2613659|Astragalus ochrochlorus
C2613659|Astragalus ocrochlorus
C2613659|Astragalus ochrochlorus Boiss. & Hohen.
C2613660|Astragalus paralipomenus
C2613660|Astragalus paralipomenus Bunge
C2613661|Astragalus paralurges
C2613661|Astragalus paralurges Bunge
C2613662|Astragalus pauperiflorus
C2613662|Astragalus pauperiflorus Bornm.
C2613663|Astragalus pellitus
C2613663|Astragalus pellitus Bunge
C2613664|Astragalus penetratus
C2613664|Astragalus penetratus A.A.Maassoumi
C2613665|Astragalus plagiophacos
C2613665|Astragalus plagiophacos Maassoumi & Podlech
C2613666|Astragalus podocarpus C.A.Mey.
C2613666|Astragalus podocarpus
C2613667|Astragalus pseudonobilis
C2613667|Astragalus pseudonobilis Popov
C2613668|Astragalus pycnocephalus
C2613668|Astragalus pycnocephalus Fisch.
C2613669|Astragalus recognitus
C2613669|Astragalus recognitus Fisch.
C2613670|Astragalus refractus
C2613670|Astragalus refractus C.A.Mey.
C2613671|Astragalus ruscifolius
C2613671|Astragalus ruscifolius Boiss.
C2613672|Astragalus saxifractor
C2613672|Astragalus saxifractor Rech.f. & Gilli
C2613672|Astragalus saxifractor Rech.f. & Gil
C2613673|Astragalus sciureus
C2613673|Astragalus sciureus Boiss. & Hohen.
C2613674|Astragalus semnanensis
C2613674|Astragalus semnanensis Bornm. & Rech.f.
C2613675|Astragalus sphaeranthus
C2613675|Astragalus sphaeranthus Boiss.
C2613676|Astragalus stevenianus
C2613676|Astragalus stevenianus DC.
C2613677|Astragalus supervisus
C2613677|Astragalus supervisus (Kuntze) E.Sheld.
C2613678|Astragalus talimansurensis
C2613678|Astragalus talimansurensis Sirj. & Rech.f.
C2613679|Astragalus tarumensis
C2613679|Astragalus tarumensis Sirj. & Rech.f.
C2613680|Astragalus thlaspi
C2613680|Astragalus thlaspi Lipsky
C2613681|Astragalus ulodjensis
C2613681|Astragalus ulodjensis Sirj. & Rech.f.
C2613682|Astragalus xanthomeloides
C2613682|Astragalus xanthomeloides Korovin & Popov
C2757825|Astragalus membranaceus var. mongholicus (Bunge) P.K.Hsiao
C2757825|Astragalus penduliflorus subsp. mongholicus
C2757825|Astragalus penduliflorus var. mongholicus
C2757825|Astragalus penduliflorus var. mongholicus (Bunge) X.Y.Zhu
C2757825|Astragalus mongholicus Bunge
C2757825|Astragalus penduliflorus subsp. mongholicus var. mongholicus
C2757825|Astragalus penduliflorus subsp. mongholicus (Bunge) X.Y.Zhu
C2757825|Astragalus mongholicus
C2757825|Astragalus membranaceus var. mongholicus
C2761350|Astragalus alopecuroides
C2761350|non Astragalus alopecuroides Ledeb., nom. illeg.
C2761350|Astragalus alopecuroides L.
C2761350|non Astragalus alopecuroides Pall., nom. illeg.
C2761351|Astragalus exscapus L
C2761351|Astragalus exscapus
C2763835|Astragalus variabilis Bunge ex Maxim.
C2763835|Astragalus variabilis
C2773106|Astragalus memoriosus
C2773106|Astragalus memoriosus M.Pakravan, Y.Nasseh & Maassoumi
C2775661|Astragalus camptodontoides N.D. Simpson
C2775661|Astragalus camptodontoides
C2775662|Astragalus camptodontus
C2775662|Phyllolobium camptodontum
C2775662|Phyllolobium camptodontum (Franch.) M.L.Zhang & Podl.
C2775662|Astragalus camptodontus Franch.
C2775663|Astragalus craibianus
C2775663|Astragalus craibianus N.D.Simpson
C2775664|Phyllolobium flavovirens (K.T.Fu) M.L.Zhang & Podl.
C2775664|Astragalus flavovirens
C2775664|Astragalus flavovirens K.T.Fu
C2775664|Phyllolobium flavovirens
C2775665|Astragalus heydei
C2775665|Phyllolobium heydei (Baker) M.L.Zhang & Podl.
C2775665|Astragalus heydei Baker
C2775665|Phyllolobium heydei
C2775666|Astragalus lasaensis
C2775666|Phyllolobium lasaense
C2775666|Astragalus lasaensis C.C.Ni & P.C.Li
C2775666|Phyllolobium lasaense (C.C.Ni & P.C.Li) M.L.Zhang & Podl.
C2775667|Phyllolobium pastorium (Tsai & T.T.Yu) M.L.Zhang & Podl.
C2775667|Phyllolobium pastorium
C2775667|Astragalus pastorius
C2775667|Astragalus pastorius Tsai & T.T.Yu
C2775668|Phyllolobium prodigiosum
C2775668|Astragalus prodigiosus K.T.Fu
C2775668|Astragalus prodigiosus
C2775668|Phyllolobium prodigiosum (K.T.Fu) M.L.Zhang & Podl.
C2775669|Astragalus sanbilingensis Tsai & T.T.Yu
C2775669|Astragalus sanbilingensis
C2775669|Phyllolobium sanbilingense
C2775669|Phyllolobium sanbilingense (Tsai & T.T.Yu) M.L.Zhang & Podl.
C2775670|Phyllolobium siccaneum (P.C.Li) M.L.Zhang & Podl.
C2775670|Astragalus siccaneus
C2775670|Astragalus siccaneus P.C.Li
C2775670|Phyllolobium siccaneum
C2775671|Phyllolobium turgidocarpum (K.T.Fu) M.L.Zhang & Podl.
C2775671|Phyllolobium turgidocarpum
C2775671|Astragalus turgidocarpus K.T.Fu
C2775671|Astragalus turgidocarpus
C2776091|Astragalus devesae Talavera, A.Gonzalaez & G.Lopez
C2776091|Astragalus devesae
C2791632|Astragalus angustifoliolatus
C2791632|Astragalus angustifoliolatus K.T.Fu
C2791871|Astragalus ansinii Uzun, Terzioglu & Palabas-Uzun
C2791871|Astragalus ansinii
C2791872|Astragalus viridissimus Freyn & Sint.
C2791872|Astragalus viridissimus
C2792644|Astragalus drummondii
C2792644|Astragalus drummondii Douglas ex Hook.
C2792645|Astragalus leptocarpus
C2792645|Astragalus leptocarpus Torr. & A.Gray
C2792646|Astragalus pectinatus
C2792646|Astragalus pectinatus (Hook.) Douglas ex G.Don
C2792647|Astragalus racemosus Pursh
C2792647|Astragalus racemosus
C2793359|Astragalus schelichowii Turcz.
C2793359|Astragalus schelichowii
C2793360|Astragalus eucosmus subsp. sealei
C2793360|Astragalus eucosmus subsp. sealei (Lepage) Hulten
C2793360|Astragalus sealei
C2793360|Astragalus sealei Lepage
C2793361|Astragalus tolmaczevii
C2793361|Astragalus tolmaczevii Jurtzev
C2797066|Astragalus chrysochlorus Boiss. & Kotschy
C2797066|Astragalus chrysochlorus
C2809829|Astragalus candolleanus Benth.
C2809829|Astragalus rhizanthus subsp. candolleanus
C2809829|Astragalus candolleanus
C2809829|non Astragalus candolleanus Boiss., nom. illeg.
C2809829|Astragalus rhizanthus subsp. candolleanus (Benth.) Podlech
C2809829|Astragalus rhizanthus subsp. candolleanus (Royle ex Benth.) Podlech
C2809829|Astragalus candolleanus Royle ex Benth.
C2809830|Astragalus malacophyllus
C2809830|Astragalus malacophyllus Bunge
C2809830|Astragalus malacophyllus Benth. ex Bunge
C2809831|Astragalus candolleanus var. pindreensis
C2809831|Astragalus pindreensis
C2809831|Astragalus pindreensis (Benth. ex Baker f.) Ali
C2809831|Astragalus candolleanus var. pindreensis Benth. ex Baker f.
C2816029|Astragalus vesicarius
C2816029|Astragalus vesicarius L.
C2816559|Astragalus hancockii
C2816559|Astragalus hancockii Bunge ex Maxim.
C2822816|Astragalus crotalariae
C2822816|Astragalus crotalariae A.Gray
C2989006|Astragalus melilotoides
C2989006|Astragalus melilotoides Pall.
C2989306|Astragalus capillipes M.E.Jones
C2989306|Astragalus capillipes
C2989306|Astragalus trichopodus
C2989306|Astragalus trichopodus (Nutt.) A.Gray
C3053096|Astragalus tragacantha
C3053096|Astragalus tragacantha L.
C3081056|Astragalus borealimongolicus
C3081056|Astragalus borealimongolicus Y.Z.Zhao
C3081057|Astragalus zacharensis Bunge
C3081057|Astragalus zacharensis
C3084604|Astragalus striatus
C3084604|Astragalus striatus Nutt.
C3086465|Astragalus bifidus
C3086465|Astragalus bifidus Turcz. ex Ledeb.
C3086466|Astragalus olchonensis Gontsch.
C3086466|Astragalus olchonensis
C3086467|Astragalus versicolor Pall.
C3086467|Astragalus versicolor
C3127924|Astragalus stereocalyx Bornm.
C3127924|Astragalus stereocalyx
C3357778|Astragalus antalyensis
C3357778|Astragalus antalyensis A.Duran & Podl.
C3357779|Astragalus apricus Bunge
C3357779|Astragalus apricus
C3357780|Astragalus avicennicus Parsa
C3357780|Astragalus avicennicus
C3357781|Astragalus caprinus L.
C3357781|Astragalus caprinus
C3357782|Astragalus chrysanthus Boiss. & Hohen.
C3357782|Astragalus chrysanthus
C3357783|Astragalus echinops
C3357783|Astragalus echinops Aucher ex Boiss.
C3357784|Astragalus gaubae
C3357784|Astragalus gaubae Bornm.
C3357785|Astragalus gypsocola
C3357785|Astragalus gypsocola Maassoumi & Mozaff.
C3357786|Astragalus impexus Podlech
C3357786|Astragalus impexus
C3357787|Astragalus ischredensis
C3357787|Astragalus ischredensis Bunge
C3357788|Astragalus johannis
C3357788|Astragalus johannis Boiss.
C3357789|Astragalus kashmarensis
C3357789|Astragalus kashmarensis Maassoumi & Podlech
C3357790|Astragalus kermanschahensis Bornm.
C3357790|Astragalus kermanschahensis
C3357791|Astragalus kirpicznikovii
C3357791|Astragalus kirpicznikovii Grossh.
C3357792|Astragalus leonardii
C3357792|Astragalus leonardii Maassoumi
C3357793|Astragalus macropelmatus Bunge
C3357793|Astragalus macropelmatus
C3357794|Astragalus mozaffarianii
C3357794|Astragalus mozaffarianii Maassoumi
C3357795|Astragalus neopodlechii
C3357795|Astragalus neopodlechii Maassoumi
C3357796|Astragalus ovinus
C3357796|Astragalus ovinus Boiss.
C3357797|Astragalus pinetorum
C3357797|Astragalus pinetorum Boiss.
C3357798|Astragalus ponticus
C3357798|Astragalus ponticus Pall.
C3357799|Astragalus pseudobrachystachys Sirj. & Rech.f.
C3357799|Astragalus pseudobrachystachys
C3357800|Astragalus pseudoibicinus
C3357800|Astragalus pseudoibicinus Maassoumi & Podlech
C3357801|Astragalus remotijugus Boiss. & Hohen.
C3357801|Astragalus remotijugus
C3357802|Astragalus reshadensis
C3357802|Astragalus reshadensis Podlech
C3357802|Astragalus reshadianus
C3357803|Astragalus rufescens Freyn & Bornm.
C3357803|Astragalus rufescens
C3357804|Astragalus touranicus
C3357804|Astragalus touranicus Freitag & Podlech
C3357805|Astragalus vanillae
C3357805|Astragalus vanillae Boiss.
C3388311|Astragalus albicaulis
C3388311|Astragalus albicaulis DC.
C3388312|Astragalus asper Jacq.
C3388312|Astragalus asper
C3388313|Astragalus pallescens
C3388313|Astragalus pallescens M.Bieb.
C3388314|Astragalus peterfii
C3388314|Astragalus peterfii Javorka
C3388315|Astragalus tarchankuticus
C3388315|Astragalus tarchankuticus Boriss.
C3388316|Astragalus ucrainicus Popov & Klokov
C3388316|Astragalus ucrainicus
C3388317|Astragalus varius
C3388317|Astragalus varius S.G.Gmel.
C3389177|Astragalus holmgreniorum
C3389177|Astragalus holmgreniorum Barneby
C3395328|Astragalus onobrychis L.
C3395328|Astragalus onobrychis
C3457541|Astragalus danicus Retz.
C3457541|Astragalus danicus
C3900926|Astragalus strictus Graham ex Benth.
C3900926|Astragalus strictus
C3336430|Astragalus aboriginum var. richardsonii (E.Sheld.) B.Boivin
C3336430|Astragalus richardsonii E.Sheld.
C3336430|Astragalus aboriginum var. richardsonii
C3336430|Astragalus richardsonii
C3586109|Astragalus macrocephalus
C3586109|Astragalus macrocephalus Willd.
C3617674|Astragalus umbraticus E.Sheld.
C3617674|Astragalus umbraticus
C3617674|Astragalus sylvaticus S.Watson, 1888, non Willd., 1802
C3617670|Astragalus oniciformis Barneby
C3617670|Astragalus oniciformis
C3586113|Astragalus neoassadianus Ranjbar
C3586113|Astragalus neoassadianus
C3564626|Astragalus sulcatus
C3564626|Astragalus sulcatus L.
C3617668|Astragalus howellii A.Gray
C3617668|Astragalus howellii
C3586114|Astragalus phlomoides Boiss.
C3586114|Astragalus phlomoides
C3617669|Astragalus misellus
C3617669|Astragalus misellus S.Watson
C3586118|Astragalus turbinatus
C3586118|Astragalus turbinatus Bunge
C3617666|Astragalus agnicidus
C3617666|Astragalus agnicidus Barneby
C3564624|Astragalus scopiformis Ledeb.
C3564624|Astragalus scopaeformis
C3564624|Astragalus scopiformis
C3586111|Astragalus melanophrurius Boiss.
C3586111|Astragalus melanophrurius
C3564622|Astragalus hispanicus
C3564622|Astragalus hispanicus Coss. ex Bunge
C3564625|Astragalus spruneri
C3564625|Astragalus spruneri Boiss.
C3609914|Astragalus wolgensis
C3609914|Astragalus wolgensis Bunge
C3564620|Astragalus contortuplicatus L.
C3564620|Astragalus contortuplicatus
C3594871|Astragalus nakaianus Y.N.Lee
C3594871|Astragalus nakaianus
C3586116|Astragalus schahrudensis Bunge
C3586116|Astragalus schahrudensis
C3586102|Astragalus ajubensis Bunge
C3586102|Astragalus ajubensis
C3586120|Astragalus zarjabadensis Ranjbar
C3586120|Astragalus zarjabadensis
C3586106|Astragalus foliosus
C3586106|Astragalus foliosus Podlech, Maassoumi & Ranjbar
C3574165|Astragalus hymenocalyx Boiss.
C3574165|Astragalus hymenocalyx
C3586104|Astragalus bezudensis
C3586104|Astragalus bezudensis Sirj. & Rech.f.
C3617672|Astragalus peckii
C3617672|Astragalus peckii Piper
C3586107|Astragalus hamadanus
C3586107|Astragalus hamadanus Boiss.
C3564623|Astragalus nummularius Lam., non Desf., 1799
C3564623|Astragalus nummularius
C3617667|Astragalus congdonii S.Watson
C3617667|Astragalus congdonii
C3586110|Astragalus megalotropis C.A.Mey. ex Bunge
C3586110|Astragalus megalotropis
C3586103|Astragalus alopecurus Pall.
C3586103|Astragalus alopecurus
C3586115|Astragalus saetiger
C3586115|Astragalus saetiger Becht
C3586117|Astragalus speciosus
C3586117|Astragalus speciosus Boiss. & Hohen.
C3617671|Astragalus paysonii (Rydb.) Barneby
C3617671|Astragalus paysonii
C3586105|Astragalus caryolobus Bunge
C3586105|Astragalus caryolobus
C3564621|Astragalus dasyanthus
C3564621|Astragalus dasyanthus Pall.
C3558102|Astragalus vesicarius subsp. pseudoglaucus Ciocarlan & Serb.
C3558102|Astragalus vesicarius subsp. pseudoglaucus
C3558102|Astragalus pseudoglaucus
C3558102|Astragalus pseudoglaucus Klokov
C3586108|Astragalus maabudii Ranjbar
C3586108|Astragalus maabudii
C3589903|Astragalus helmii
C3589903|Astragalus helmii Fisch. ex DC.
C3586119|Astragalus victoriae
C3586119|Astragalus victoriae (Podl. & Kirchhoff) Podl. & Kirchhoff
C3586112|Astragalus meridionalis Bunge
C3586112|Astragalus meridionalis
C3617673|Astragalus toquimanus
C3617673|Astragalus toquimanus Barneby
C3725786|Astragalus scholerianus
C3725786|Astragalus scholerianus Bornm.
C3797027|Astragalus tortuosus DC.
C3797027|Astragalus tortuosus
C3731256|Astragalus lepidanthus
C3731007|Astragalus nutzotinensis
C3731007|Astragalus nutzotinensis J.Rousseau
C3731007|Gynophoraria falcata Rydb., non Astragalus falcatus Lam.
C3720512|Astragalus brevipes
C3720512|Astragalus brevipes Bunge
C3797003|Astragalus bodeanus Fisch.
C3797003|Astragalus bodeanus
C3731242|Astragalus angustifolius
C3725767|Astragalus gladiatus
C3725767|Astragalus gladiatus Boiss.
C3725756|Astragalus brevidentatus
C3725756|Astragalus brevidentatus C.H.Wright
C3797029|Astragalus veiskaramii Zarre, Podl. & Sabaii
C3797029|Astragalus veiskaramii
C3797007|Astragalus crassispinus
C3797007|Astragalus crassispinus Bunge
C3720324|Astragalus juladakensis Maassoumi
C3720324|Astragalus juladakensis
C3720333|Astragalus xiphidium Bunge
C3720333|Astragalus xiphidium
C3725763|Astragalus dasycarpus D.F.Chamb.
C3725763|Astragalus dasycarpus
C3726053|Astragalus sp. A20
C3731257|Astragalus macrocarpus
C3720321|Astragalus djenarensis
C3720321|Astragalus djenarensis Sirj. & Rech.f.
C3725790|Astragalus tigridis
C3725790|Astragalus tigridis Boiss.
C3731255|Astragalus kurnet-es-saudae
C3725766|Astragalus germanicopolitanus Bornm.
C3725766|Astragalus germanicopolitanus
C3720316|Astragalus aestimabilis Podlech
C3720316|Astragalus aestimabilis
C3731246|Astragalus cedreti
C3725771|Astragalus lasioglottis M.Bieb.
C3725771|Astragalus lasioglottis
C3720323|Astragalus husseinovii
C3720323|Astragalus husseinovii Rzazade
C3725788|Astragalus subulatus Desf.
C3725788|Astragalus subulatus
C3804432|Astragalus sp. A108
C3797008|Astragalus cymbostegis Bunge
C3797008|Astragalus cymbostegis
C3720319|Astragalus baraftabensis Maassoumi & Podlech
C3720319|Astragalus baraftabensis
C3720521|Astragalus psoraloides Lam.
C3720521|Astragalus psoraloides
C3725755|Astragalus brachycarpus M.Bieb.
C3725755|Astragalus brachycarpus
C3720513|Astragalus effusus Bunge
C3720513|Astragalus effusus
C3720516|Astragalus jodostachys
C3720516|Astragalus jodostachys Boiss. & Buhse
C3725787|Astragalus sigmoideus
C3725787|Astragalus sigmoideus Bunge
C3797010|Astragalus dipodurus
C3797010|Astragalus dipodurus Bunge
C3720523|Astragalus sevangensis
C3720523|Astragalus sevangensis Grossh.
C3725784|Astragalus scabrifolius
C3725784|Astragalus scabrifolius Boiss.
C3725750|Astragalus achundovii
C3725750|Astragalus achundovii Grossh.
C3725775|Astragalus nezaketiae
C3725775|Astragalus nezaketiae A.Duran & Aytac
C3725775|Astragalus nezaketae
C3725760|Astragalus clavatus
C3725760|Astragalus clavatus DC.
C3722957|Astragalus flexuosus (Hook.) Douglas ex G.Don
C3722957|Astragalus flexuosus
C3720332|Astragalus viridis
C3720332|Astragalus viridis Bunge
C3725769|Astragalus hartvigii Kit Tan
C3725769|Astragalus hartvigii
C3731241|Astragalus angulosus
C3720329|Astragalus saadatabadensis Podlech
C3720329|Astragalus saadatabadensis
C3797002|Astragalus aureus
C3797002|Astragalus aureus Willd.
C3797024|Astragalus rubrolineatus
C3797024|Astragalus rubrolineatus Sirj. & Rech.f.
C3725774|Astragalus micrancistrus
C3725774|Astragalus micrancistrus Boiss. & Hausskn.
C3797005|Astragalus clusianus
C3797005|Astragalus clusianus (Boiss.) Soldano, nom. illeg.
C3797005|Astragalus clusii Boiss.
C3797005|Astragalus clusii
C3720526|Astragalus vegetus
C3720526|Astragalus vegetus Bunge
C3725770|Astragalus kastamonuensis D.F.Chamb. & V.A.Matthews
C3725770|Astragalus kastamonuensis
C3797030|Astragalus wagneri
C3797030|Astragalus wagneri Bartl. ex Bunge
C3720325|Astragalus juratzkanus Freyn & Sint.
C3720325|Astragalus juratzkanus
C3720514|Astragalus goktschaicus
C3720514|Astragalus goktschaicus Grossh.
C3725762|Astragalus czorochensis
C3725762|Astragalus czorochensis Kharadze
C3731254|Astragalus hirsutissimus
C3731250|Astragalus dictyocarpus
C3781921|Astragalus spinosus
C3781921|Astragalus spinosus (Forssk.) Muschl.
C3725794|Astragalus yildirimlii Aytac & Ekici
C3725794|Astragalus yildirimlii
C3725776|Astragalus nigrifructus Podlech & Aytac
C3725776|Astragalus nigrifructus
C3725753|Astragalus bachmarensis
C3725753|Astragalus bachmarensis Grossh.
C3720520|Astragalus parvarensis
C3720520|Astragalus parvarensis Podl. & Sytin
C3725779|Astragalus oreades
C3725779|Astragalus oreades C.A.Mey.
C3797021|Astragalus raddei Basil.
C3797021|Astragalus raddei
C3731253|Astragalus emarginatus
C3725781|Astragalus polhillii
C3725781|Astragalus polhillii Podlech
C3720328|Astragalus pravitzii
C3720328|Astragalus pravitzii Podlech
C3720517|Astragalus lunatus Gilib.
C3720517|Astragalus lunatus
C3720517|Astragalus lunatus Pall.
C3725758|Astragalus cedreticola
C3725758|Astragalus cedreticola A.Duran & Podlech
C3720320|Astragalus dendroproselius
C3720320|Astragalus dendroproselius Rech.f.
C3731251|Astragalus ehdenensis
C3725780|Astragalus ovatus
C3725780|Astragalus ovatus DC.
C3723004|Astragalus keredjensis (Bornm. & Gauba) Podl.
C3723004|Astragalus keredjensis
C3731258|Astragalus psilodontius
C3720318|Astragalus aucheri Boiss.
C3720318|Astragalus aucheri
C3720509|Astragalus arguricus Bunge
C3720509|Astragalus arguricus
C3731245|Astragalus bethlehemiticus
C3797011|Astragalus distans Fisch.
C3797011|Astragalus distans
C3720326|Astragalus melanocalyx
C3720326|Astragalus melanocalyx Boiss. & Buhse
C3731259|Astragalus trichopterus
C3731259|Astragalus nummularius subsp. trichopterus
C3797019|Astragalus megalocystis
C3797019|Astragalus megalocystis Bunge
C3797009|Astragalus diphtherites
C3797009|Astragalus diphtherites Fenzl
C3725768|Astragalus glaucophyllus
C3725768|Astragalus glaucophyllus Bunge
C3726052|Astragalus sp. A2
C3797006|Astragalus coluteopsis Parsa
C3797006|Astragalus coluteopsis
C3797014|Astragalus ghashghaicus
C3797014|Astragalus ghashghaicus Tietz & Zarre
C3797012|Astragalus ebenoides Boiss.
C3797012|Astragalus ebenoides
C3797023|Astragalus remotiflorus Boiss.
C3797023|Astragalus remotiflorus
C3797001|Astragalus anthylloides
C3797001|Astragalus anthylloides Lam.
C3726055|Astragalus sp. A35
C3797020|Astragalus microphysa Boiss.
C3797020|Astragalus microphysa
C3720524|Astragalus sufianicus
C3720524|Astragalus sufianicus Podl. & Sytin
C3797025|Astragalus susianus
C3797025|Astragalus susianus Boiss.
C3720334|Astragalus zoshkensis
C3720334|Astragalus zoshkensis Ghahr.-Nejad
C3725795|Astragalus zaraensis Podlech
C3725795|Astragalus zaraensis
C3725783|Astragalus sanguinolentus M.Bieb.
C3725783|Astragalus sanguinolentus
C3725777|Astragalus nitens Boiss. & Heldr.
C3725777|Astragalus nitens
C3720330|Astragalus sitiens
C3720330|Astragalus sitiens Bunge
C3731247|Astragalus cephalotes
C3725752|Astragalus ancistrocarpus
C3725752|Astragalus ancistrocarpus Boiss. & Hausskn.
C3720522|Astragalus scapiger Ranjbar & Maassoumi
C3720522|Astragalus scapiger
C3720327|Astragalus nigrolineatus
C3720327|Astragalus nigrolineatus Sirj. & Rech.f.
C3725754|Astragalus beypazaricus
C3725754|Astragalus beypazaricus Podlech & Aytac
C3720525|Astragalus trifoliolatus
C3720525|Astragalus trifoliolatus Boiss.
C3725761|Astragalus cornutus
C3725761|Astragalus cornutus Pall.
C3726054|Astragalus sp. A3
C3731243|Astragalus baalbekensis
C3720508|Astragalus aduncus Willd.
C3720508|Astragalus aduncus
C3725793|Astragalus viciifolius DC.
C3725793|Astragalus viciaefolius
C3725793|Astragalus viciifolius
C3725764|Astragalus elongatus Willd.
C3725764|Astragalus elongatus
C3797022|Astragalus raswendicus Hausskn. & Bornm.
C3797022|Astragalus raswendicus
C3797026|Astragalus szovitsii
C3797026|Astragalus szovitsii Fisch. & C.A.Mey.
C3731244|Astragalus berytheus
C3725773|Astragalus melanocarpus
C3725773|Astragalus melanocarpus Richardson
C3726049|Astragalus sp. A109
C3725782|Astragalus saganlugensis Trautv.
C3725782|Astragalus saganlugensis
C3725759|Astragalus cinereus Willd.
C3725759|Astragalus cinereus
C3797016|Astragalus keratensis
C3797016|Astragalus keratensis Bunge
C3720510|Astragalus bijarensis Podl. & Sytin
C3720510|Astragalus bijarensis
C3725792|Astragalus vexillaris Boiss.
C3725792|Astragalus vexillaris
C3797018|Astragalus lumsdenianus Aitch.
C3797018|Astragalus lumsdenianus
C3797017|Astragalus lalesarensis
C3797017|Astragalus lalesarensis Bornm.
C3726058|Astragalus sp. A66
C3797028|Astragalus vaginans
C3797028|Astragalus vaginans DC.
C3720331|Astragalus sumbari Popov
C3720331|Astragalus sumbari
C3731260|Astragalus zachlensis
C3726051|Astragalus sp. A16
C3720518|Astragalus neochaldoranicus
C3720518|Astragalus neochaldoranicus Podlech & Maassoumi
C3720518|Astragalus chaldoranicus Podlech & Maassoumi, non Astragalus chaldiranicus Kit Tan & Sorger
C3720519|Astragalus oligoflorus
C3720519|Astragalus oligoflorus Maassoumi, Ghahrem. & Javadi
C3734172|Astragalus drusorum
C3720317|Astragalus argyroides Beck ex Stapf
C3720317|Astragalus argyroides
C3725751|Astragalus akmanii
C3725751|Astragalus akmanii Aytac & H.Duman
C3725789|Astragalus taochius Woronow
C3725789|Astragalus taochius
C3725778|Astragalus olurensis
C3725778|Astragalus olurensis Podlech
C3720322|Astragalus eburneus Bornm. & Gauba
C3720322|Astragalus eburneus
C3726057|Astragalus sp. A65
C3720515|Astragalus huthianus
C3720515|Astragalus huthianus Freyn & Bornm.
C3797004|Astragalus chardini
C3797004|Astragalus chardinii
C3797004|Astragalus chardinii Boiss.
C3720527|Astragalus xerophilus
C3720527|Astragalus xerophilus Ledeb.
C3725785|Astragalus schizopterus
C3725785|Astragalus schizopterus Boiss.
C3726056|Astragalus sp. A52
C3797013|Astragalus gevashensis
C3797013|Astragalus gevashensis D.F.Chamb. & V.A.Matthews
C3720511|Astragalus brachyodontus
C3720511|Astragalus brachyodontus Boiss.
C3725765|Astragalus frickii
C3725765|Astragalus frickii Bunge
C3731248|Astragalus coluteoides
C3781920|Astragalus sieberi
C3781920|Astragalus sieberi DC.
C3797015|Astragalus halicacabus Lam.
C3797015|Astragalus halicacabus
C3731252|Astragalus ehrenbergii
C3722958|Astragalus laxmannii Jacq.
C3722958|Astragalus laxmannii
C3726050|Astragalus sp. A110
C3725791|Astragalus turkmenensis
C3725791|Astragalus turkmenensis Dural, Tugay & Ertugrul
C3725772|Astragalus longisubulatus Podlech
C3725772|Astragalus longisubulatus
C3731249|Astragalus cruentiflorus
C3725757|Astragalus cariensis Boiss.
C3725757|Astragalus cariensis
C3908984|Astragalus oligophyllus
C3908984|Astragalus oligophyllus Boiss.
C3908979|Astragalus joharchii
C3908979|Astragalus joharchii F.Ghahrem. & Gaskin
C3908967|Astragalus baharensis
C3908967|Astragalus baharensis F.Ghahrem.
C3908990|Astragalus sangonensis Sirj. & Rech.f.
C3908990|Astragalus sangonensis
C3908966|Astragalus ammodendron
C3908966|Astragalus ammodendron Bunge
C3908965|Astragalus akhundzadahensis
C3908965|Astragalus akhundzadahensis Podl. & Zarre
C3908972|Astragalus erwinii-gaubae Sirj. & Rech.f.
C3908972|Astragalus erwinii-gaubae
C3959806|Astragalus davuricus (Pall.) DC.
C3959806|Astragalus davuricus
C3908975|Astragalus ghamishluensis
C3908975|Astragalus ghamishluensis Dastpak, Maassoumi & Kaz.Osaloo
C3908986|Astragalus podoloboides Maassoumi
C3908986|Astragalus podoloboides
C3908982|Astragalus nigricans
C3908982|Astragalus nigrescens Popov, 1947, non Pall., 1800
C3908982|Astragalus nigricans Barneby
C3908980|Astragalus kavirensis
C3908980|Astragalus kavirensis Freitag
C3956686|Astragalus arenarius
C3956686|Astragalus arenarius L.
C3908976|Astragalus griffithii
C3908976|Astragalus griffithii Benth. ex Bunge
C3908988|Astragalus pseudoarvatensis
C3908988|Astragalus pseudoarvatensis Podl. & Sytin
C3908994|Astragalus tabrizianus
C3908994|Astragalus tabrizianus Buhse
C3908981|Astragalus karakugensis
C3908981|Astragalus karakugensis Bunge
C3908968|Astragalus bazarganii Podl. & Zarre
C3908968|Astragalus bazarganii
C3908977|Astragalus inchebroonensis Maassoumi
C3908977|Astragalus inchebroonensis
C3908973|Astragalus farsicus Sirj. & Rech.f.
C3908973|Astragalus farsicus
C3999434|Astragalus trifoliastrum Hub.-Mor. & V.A.Matthews
C3999434|Astragalus trifoliastrum
C3908970|Astragalus brevicalycinus Maassoumi
C3908970|Astragalus brevicalycinus
C3999432|Astragalus assadabadensis F.Ghahrem. & Podlech
C3999432|Astragalus assadabadensis
C3908971|Astragalus darrehbidensis
C3908971|Astragalus darrehbidensis Podl. & Zarre
C3908978|Astragalus jaskensis
C3908978|Astragalus jaskensis Maassoumi
C3908991|Astragalus semiglabricarpus Maassoumi
C3908991|Astragalus semiglabricarpus
C3908987|Astragalus podolobus Boiss. & Hohen.
C3908987|Astragalus podolobus
C3966917|Astragalus sp. PMD-2014
C3999433|Astragalus laguriformis Freyn
C3999433|Astragalus laguriformis
C3908993|Astragalus tenuiramosus
C3908993|Astragalus tenuiramosus Podl. & Zarre
C3908974|Astragalus gebleri Bong.
C3908974|Astragalus gebleri
C3908969|Astragalus biarjmandicus
C3908969|Astragalus biarjmandicus Podl. & Zarre
C3908989|Astragalus pseudonigrescens Maassoumi
C3908989|Astragalus pseudonigrescens
C3909260|Astragalus acutifolius Bunge, 1868
C3909260|Astragalus acutifolius
C3908985|Astragalus ovalis Boiss. & Balansa
C3908985|Astragalus ovalis
C3908983|Astragalus oldenburgii B.Fedtsch.
C3908983|Astragalus oldenburgii
C3908992|Astragalus sympileicalycinus Maassoumi & Nasseh
C3908992|Astragalus sympileicalycinus
C0330847|Astragalus lentiginosus
C0330847|Astragalus lentiginosus Douglas ex Hook.
C0330847|Astragalus lentiginosus (organism)
C0330846|Astragalus pubentissimus
C0330846|Astragalus pubentissimus (organism)
C1040224|Astragalus australis
C1040224|Astragalus australis (L.) Lam.
C1040219|Astragalus alvordensis
C1040219|Astragalus alvordensis M.E.Jones
C1001107|Astragalus brandegei
C1001107|Astragalus brandegeei Porter
C1092198|Astragalus penduliflorus Lam.
C1092198|Astragalus penduliflorus
C1031852|Astragalus sparsus
C1031852|Astragalus sparsus Decne.
C1001111|Astragalus cremnophylax
C1001111|Astragalus cremnophylax Barneby
C1075622|Astragalus austrosibiricus
C1075622|Astragalus austrosibiricus Schischk.
C1040276|Astragalus umbellatus
C1040276|Astragalus umbellatus Bunge
C1013040|Astragalus complanatus
C1013040|Astragalus complanatus R.Br. ex Bunge
C1040240|Astragalus eremiticus
C1040240|Astragalus eremiticus E.Sheld.
C1001105|Astragalus asterias
C1001105|Astragalus asterias Steven
C1086980|Astragalus williamsii
C1086980|Astragalus williamsii Britton & Rydb.
C1040229|Astragalus chamaemeniscus
C1040229|Astragalus chamaemeniscus Barneby
C1040226|Astragalus calycosus
C1040226|Astragalus calycosus Torr. ex S.Watson
C1086972|Astragalus molybdenus
C1086972|Astragalus molybdenus Barneby
C1094369|Astragalus tener
C1094369|Astragalus tener A.Gray
C1075621|Astragalus aksuensis
C1075621|Astragalus aksuensis Bunge
C1001119|Astragalus pulchellus
C1001122|Astragalus thurberi
C1001122|Astragalus thurberi A.Gray
C1001108|Astragalus chaborasicus
C1001108|Astragalus chaborasicus Boiss. & Hausskn.
C1081363|Astragalus tribuloides
C1081363|Astragalus tribuloides Delile
C1040220|Astragalus arizonicus
C1040220|Astragalus arizonicus A.Gray
C1040246|Astragalus kentrophyta A.Gray
C1040246|Astragalus kentrophyta
C1040271|Astragalus sheldonii
C1040271|Astragalus sheldonii (Rydb.) Barneby
C1086976|Astragalus polaris
C1040234|Astragalus curvicarpus
C1040234|Astragalus curvicarpus (E.Sheld.) J.F.Macbr.
C1082960|Astragalus peristereus
C1040241|Astragalus eucosmus
C1040241|Astragalus eucosmus B.L.Rob.
C1013031|Astragalus americanus
C1013031|Astragalus americanus (Hook.) M.E.Jones
C1001123|Astragalus utahensis
C1001123|Astragalus utahensis (Torr.) Torr. & A.Gray
C1040235|Astragalus cymbicarpos
C1040235|Astragalus cymbicarpos Brot.
C1001114|Astragalus humillimus
C1001114|Astragalus humillimus A.Gray
C1086975|Astragalus paposanus
C1040264|Astragalus polycladus
C1040273|Astragalus spatulatus
C1040273|Astragalus spatulatus E.Sheld.
C1040273|Homalobus caespitosus Nutt. 1838, non Pall., 1803
C1040252|Astragalus moyanoi
C1040252|Astragalus moyanoi Speg.
C1075625|Astragalus sieversianus Pall.
C1075625|Astragalus sieversianus
C1075624|Astragalus membranaceus f. propinquus
C1075624|Astragalus propinquus Schischkin
C1075624|Astragalus membranaceus f. propinquus (Schischkin) Kitag.
C1075624|Astragalus propinquus
C1086974|Astragalus oreganus
C1013048|Astragalus cerasocrenus
C1013048|Astracantha cerasocrena (Bunge) Podlech
C1013048|Astragalus cerasocrenus Bunge
C1001113|Astragalus hamosus
C1001113|Astragalus hamosus L.
C1001104|Astragalus aretioides
C1001104|Orophaca aretioides (M.E.Jones) Rydb.
C1001104|Astragalus aretioides (M.E.Jones) Barneby
C1001115|Astragalus lobophorus
C1001115|Astragalus lobophorus Boiss.
C1013053|Astragalus bodinii
C1013053|Astragalus bodinii E.Sheld.
C1001118|Astragalus oocalycis
C1001112|Astragalus hallii
C1001112|Astragalus hallii A.Gray
C1001106|Astragalus bisulcatus
C1001106|Astragalus bisulcatus (Hook.) A.Gray
C1040244|Astragalus gilviflorus
C1040244|Astragalus gilviflorus E.Sheld.
C1460814|Astragalus tribulifolius Benth. ex Bunge
C1460814|Astragalus tribulifolius
C1040233|Astragalus collinus
C1040233|Astragalus collinus (Hook.) Douglas ex G.Don
C1013047|Astragalus atropilosulus
C1013047|Astragalus atropilosulus (Hochst.) Bunge
C1040228|Astragalus ceramicus
C1040228|Astragalus ceramicus E.Sheld.
C1927453|Astragalus layneae
C1927453|Astragalus layneae Greene
C1040269|Astragalus sabulonum
C1040269|Astragalus sabulonum A.Gray
C1501916|Astragalus monspessulanus L.
C1501916|Astragalus monspessulanus
C1040250|Astragalus mollissimus
C1040250|Astragalus mollissimus Torr.
C1082965|Astragalus echinatus
C1082965|Astragalus echinatus Murray
C1086977|Astragalus reventus
C1086977|Astragalus reventus A.Gray
C1040275|Astragalus tetrapterus
C1040275|Astragalus tetrapterus A.Gray
C1040331|Astragalus sp. Sanderson 2509
C1040260|Astragalus palanae
C1089563|Astragalus lehmannianus
C1089563|Astragalus lehmannianus Bunge
C1040223|Astragalus asymmetricus
C1040223|Astragalus asymmetricus E.Sheld.
C1040253|Astragalus nankotaizanensis
C1040256|Astragalus nuttallii
C1040245|Astragalus inyoensis
C1040245|Astragalus inyoensis E.Sheld.
C1460810|Astragalus balfourianus N.D.Simpson
C1460810|Astragalus balfourianus
C1460813|Astragalus tanguticus Batalin
C1460813|Astragalus tanguticus
C1040248|Astragalus lindheimeri
C1040248|Astragalus lindheimeri Engelm. ex A.Gray
C1001117|Astragalus nuttallianus DC.
C1001117|Astragalus nuttallianus
C1040265|Astragalus praelongus
C1086971|Astragalus linifolius
C1086971|Astragalus linifolius Osterh.
C1040227|Astragalus caricinus
C1040227|Astragalus caricinus (M.E.Jones) Barneby
C1040277|Astragalus woodruffii
C1040277|Astragalus woodruffii M.E.Jones
C1040237|Astragalus didymocarpus
C1040237|Astragalus didymocarpus Hook. & Arn.
C1040259|Astragalus pachypus
C1040222|Astragalus arthurii M.E.Jones
C1040222|Astragalus arthurii
C1040222|Astragalus arthuri
C1040258|Astragalus oxyphysus
C1013030|Astragalus robbinsii (Oakes) A.Gray
C1013030|Astragalus robbinsii
C1001121|Astragalus scopulorum
C1001121|Astragalus scopulorum Porter
C1086392|Astragalus glycyphyllos L.
C1086392|liquorice milk-vetch
C1086392|Astragalus glycyphyllos
C1040218|Astragalus allochrous
C1040218|Astragalus allochrous A.Gray
C1040266|Astragalus preussii
C1013041|Astragalus sinicus
C1013041|Astragalus sinicus L.
C1001110|Astragalus corrugatus
C1001110|Astragalus corrugatus Bertol.
C1460812|Astragalus milingensis C.C.Ni & P.C.Li
C1460812|Astragalus milingensis
C1075623|Astragalus lepsensis
C1075623|Astragalus lepsensis Bunge
C1927452|Astragalus jaegerianus
C1927452|Astragalus jaegerianus Munz
C1040239|Astragalus edulis
C1040239|Astragalus edulis Durieu ex Coss.
C1093436|Astragalus echidnaeformis
C1093436|Astragalus echidniformis
C1093436|Astragalus echidniformis Sirj.
C1040243|Astragalus garbancillo
C1040243|Astragalus garbancillo Cav.
C1040267|Astragalus rattanii
C1040267|Astragalus rattanii A.Gray
C1040261|Astragalus patagonicus
C1013064|Astragalus vogelii
C1013064|Astragalus vogelii (Webb) Bornm.
C1094367|Astragalus asclepiadoides
C1094367|Astragalus asclepiadoides M.E.Jones
C1040249|Astragalus lonchocarpus
C1040249|Astragalus lonchocarpus Torr.
C1040221|Astragalus arnottianus
C1040221|Astragalus arnottianus (Gillies ex Hook. & Arn.) Reiche
C1040270|Astragalus salmonis
C1040270|Astragalus salmonis M.E.Jones
C1040247|Astragalus leptaleus
C1040247|Astragalus leptaleus A.Gray
C1001101|Astragalus adsurgens
C1001101|Astragalus adsurgens Pall.
C1040238|Astragalus douglasii
C1040238|Astragalus douglasii (Torr. & A.Gray) A.Gray
C1086979|Astragalus speirocarpus
C1086979|Astragalus speirocarpus A.Gray
C1460811|Astragalus hendersonii Baker
C1460811|Astragalus hendersonii
C1040274|Astragalus tenellus
C1040274|Astragalus tenellus Pursh
C1040251|Astragalus monoensis
C1040251|Astragalus monoensis Barneby
C1001102|Astragalus agrestis
C1001102|Astragalus agrestis G.Don
C1040263|Astragalus pickeringii
C1040272|Astragalus shultziorum
C1040272|Astragalus shultziorum Barneby
C1093072|Astragalus canadensis
C1093072|Astragalus canadensis L.
C1086978|Astragalus sesquiflorus
C1086978|Astragalus sesquiflorus S.Watson
C1040232|Astragalus cobrensis
C1040232|Astragalus cobrensis A.Gray
C1082971|Astragalus epiglottis
C1082971|Astragalus epiglottis L.
C1040225|Astragalus boeticus
C1040225|Astragalus boeticus L.
C1040242|Astragalus filipes
C1040242|Astragalus filipes Torr. ex A.Gray
C1040255|Astragalus nothoxys
C1040268|Astragalus rubyi
C1040268|Astragalus rubyi Greene & Morris
C1460815|Astragalus yatungensis C.C.Ni & P.C.Li
C1460815|Astragalus yatungensis
C1040262|Astragalus pehuenches
C1013019|Astragalus falcatus
C1013019|Astragalus falcatus Lam.
C1001109|Astragalus cicer
C1001109|Astragalus cicer L.
C1094368|Astragalus miser
C1094368|Astragalus miser Douglas
C1040231|Astragalus cibarius
C1040231|Astragalus cibarius E.Sheld.
C1040230|Astragalus chinensis
C1040230|Astragalus chinensis L.f.
C1086973|Astragalus neuquenensis
C1040254|Astragalus neglectus
C1040257|Astragalus obscurus
C1001103|Astragalus alpinus
C1001103|Astragalus alpinus L.
C1040236|Astragalus cysticalyx
C1040236|Astragalus cysticalyx Ledeb.
C1001120|Astragalus purshii
C1001116|Astragalus monumentalis
C1001116|Astragalus monumentalis Barneby
C1013090|Astragalus alopecias
C1013090|Astragalus alopecias Pall.
C1057531|Astragalus hoantchy
C1057531|Astragalus hoantchy Franch.
C2271918|Astragalus oophorus
C2285393|Astragalus uliginosus
C2285393|Astragalus uliginosus L.
C2287240|Astragalus acutirostris
C2287240|Astragalus acutirostris S.Watson
C2287241|Astragalus casei
C2287241|Astragalus casei A.Gray ex Brewer & S.Watson
C2287242|Astragalus coccineus
C2287242|Astragalus coccineus (Parry) Brandegee
C2287243|Astragalus geyeri
C2287243|Astragalus geyeri A.Gray
C2287244|Astragalus malacus
C2287244|Astragalus malacus A.Gray
C2287245|Astragalus newberryi
C2287245|Astragalus newberryi A.Gray
C2287246|Astragalus platytropis A.Gray
C2287246|Astragalus platytropis
C2287247|Astragalus serenoi
C2287247|Astragalus serenoi (Kuntze) E.Sheld.
C2287248|Astragalus wootonii
C2287248|Astragalus wootonii E.Sheld.
C2301324|Astragalus amatus Clos
C2301324|Astragalus amatus
C2301325|Astragalus berteroanus (Moris) Reiche
C2301325|Astragalus berterianus
C2301325|Astragalus berteroanus
C2301326|Astragalus cruckshanksii (Hook. & Arn.) Griseb.
C2301326|Astragalus cruikschankii
C2301326|Astragalus cruckshanksii
C2301327|Astragalus cryptobotrys
C2301327|Phaca clandestina Phil.
C2301327|Astragalus cryptobotrys I.M.Johnst.
C2301328|Astragalus curvicaulis
C2301328|Astragalus curvicaulis (Clos) Reiche
C2301329|Astragalus darumbium (Bertero ex Colla) Clos
C2301329|Astragalus darumbium
C2301330|Astragalus edmonstonei
C2301330|Astragalus edmondstonei (Hook.f.) B.L.Rob.
C2301330|Astragalus edmondstonei
C2301331|Astragalus johnstonii
C2301331|Astragalus johnstonii Gomez-Sosa
C2301332|Astragalus looseri
C2301332|Astragalus looserii
C2301332|Astragalus looseri I.M.Johnst.
C2301333|Astragalus monticola Phil.
C2301333|Astragalus monticola
C2301334|Astragalus nivicola
C2301334|Astragalus nivicola Gomez-Sosa
C2301335|Astragalus uniflorus
C2301335|Astragalus uniflorus DC.
C2301336|Astragalus vagus
C2301336|Astragalus vagus Reiche
C2301858|Astragalus rhizanthus
C2301858|Astragalus rhizanthus Royle ex Benth.
C2310493|Astragalus armatus
C2310493|Astragalus armatus Willd.
C1095897|Astragalus preparation
C1095897|ASTRAGALUS
C1095897|astragalus (medication)
C1095897|ASTRAGALUS EXTRACT
C1177063|ASTRAGALUS EXTRACT PWDR
C1177063|ASTRAGALUS EXTRACT PWDR [VA Product]
C3864824|paritaprevir
C3864824|Paritaprevir (product)
C3864824|Paritaprevir (substance)
C3883274|PARITAPREVIR DIHYDRATE
C4046856|Technivie
C3864967|ombitasvir / paritaprevir / Ritonavir
C3864967|ombitasvir/paritaprevir/ritonavir
C3864967|ombitasvir + paritaprevir + ritonavir
C3864967|ombitasvir + paritaprevir + ritonavir (medication)
C3864967|Ombitasvir + paritaprevir + ritonavir (product)
C4075296|Oral form paritaprevir (product)
C4075296|Oral form paritaprevir
C3865211|ombitasvir / paritaprevir / Ritonavir Oral Product
C3865211|Oral form ombitasvir + paritaprevir + ritonavir
C3865211|Oral form ombitasvir + paritaprevir + ritonavir (product)
C4046961|ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG [Technivie]
C3865125|ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet
C3865125|Ombitasvir/Paritaprevir/Ritonavir 12.5 MG-75 MG-50 MG Oral Tablet
C3865125|Ombitasvir, Paritaprevir, Ritonavir 12.5-75-50mg Oral tablet
C3865125|Ombitasvir-Paritaprevir-Ritonavir Tab 12.5-75-50 MG
C3865188|ombitasvir / paritaprevir / Ritonavir Oral Tablet
C4047089|Technivie Pill
C4047040|ombitasvir / paritaprevir / Ritonavir Oral Tablet [Technivie]
C4047090|Technivie Oral Product
C3854281|{2 (dasabuvir 250 MG Oral Tablet) / 2 (ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet) } Pack [Viekira Pak]
C3854281|Viekira Pak
C3854281|Viekira Pak KIT
C3854281|Viekira Pak, oral kit
C3854281|Dasabuvir;Ombitasvir/Paritaprevir/Ritonavir NA Oral Tablet [VIEKIRA PAK]
C3864964|{2 (dasabuvir 250 MG Oral Tablet) / 2 (ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet) } Pack
C3864964|Ombitas-Paritapre-Riton & Dasab Tab Pak 12.5-75-50 & 250 MG
C3864964|DASABUVIR/OMBITASVIR/PARITAPREVIR/RITONAVIR DAILY DOSE PACK [VA Product]
C3864964|VIEKIRA DAILY PAK
C3864964|DASABUVIR/OMBITASVIR/PARITAPREVIR/RITONAVIR DAILY DOSE PACK
C3864964|TECHNIVIE DOSE PACK,56
C3864964|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56
C3864964|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DOSE PACK,56 [VA Product]
C3864964|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK [VA Product]
C3864964|OMBITASVIR 12.5/PARITAPREVIR 75/RITONAVIR 50MG TAB DAILY PACK
C3864964|TECHNIVIE DAILY PACK
C4046169|technivie 12.5 MG / 75 MG / 50 MG Oral Tablet
C4046169|Technivie KIT
C4046169|RITONAVIR 50 mg / OMBITASVIR HEMINONAHYDRATE 12.5 mg / PARITAPREVIR DIHYDRATE 75 mg ORAL TABLET, FILM COATED [Technivie]
C4046169|Technivie 12.5mg-75mg-50mg Tablet
C4046169|Ombitasvir/Paritaprevir/Ritonavir 12.5 MG-75 MG-50 MG Oral Tablet [TECHNIVIE]
C4046169|ombitasvir 12.5 MG / paritaprevir 75 MG / Ritonavir 50 MG Oral Tablet [Technivie]
C4046169|Technivie, 12.5 mg-75 mg-50 mg oral tablet
C4080053|grazoprevir
C4080455|Zepatier
C4080456|elbasvir 50 MG / grazoprevir 100 MG [Zepatier]
C4080458|Zepatier Oral Product
C4080452|elbasvir / grazoprevir Oral Tablet
C4080454|Elbasvir, Grazoprevir 50-100mg Oral tablet
C4080454|Elbasvir/Grazoprevir 50 MG-100 MG Oral Tablet
C4080454|elbasvir 50 MG / grazoprevir 100 MG Oral Tablet
C4080459|Zepatier Pill
C4080457|elbasvir / grazoprevir Oral Tablet [Zepatier]
C4080460|ZEPATIER 50mg-100mg Tablet
C4080460|Zepatier 50 MG / 100 MG Oral Tablet
C4080460|Zepatier (elbasvir 50 MG / grazoprevir 100 MG) Oral Tablet
C4080460|ELBASVIR 50 mg / GRAZOPREVIR 100 mg ORAL TABLET, FILM COATED [ZEPATIER]
C4080460|Elbasvir/Grazoprevir 50 MG-100 MG Oral Tablet [ZEPATIER]
C4080460|elbasvir 50 MG / grazoprevir 100 MG Oral Tablet [Zepatier]
C2976304|PSI-7977
C2976304|7977, PSI
C2976304|PSI7977
C2976304|PSI 7977
C3530149|GS-7977
C3530149|GS7977
C3530149|GS 7977
C2976303|L-Alanine, N-[[P(S),2'R]-2'-deoxy-2'-fluoro-2'-methyl-P-phenyl-5'-uridylyl]-, 1-methylethyl Ester
C2976303|Sofosbuvir
C2976303|antivirals sofosbuvir
C2976303|sofosbuvir (medication)
C2976303|Sofosbuvir (substance)
C2976303|2-((5-(2,4-dioxo-3,4-dihydro-2H-pyrimidin-1-yl)-4-fluoro-3-hydroxy-4-methyltetrahydrofuran-2-ylmethoxy)phenoxyphosphorylamino)propionic acid isopropyl ester
C2976303|Sofosbuvir [Chemical/Ingredient]
C2976303|Sofosbuvir (product)
C3700471|Sovaldi
C3858025|Harvoni
C3858051|ledipasvir / sofosbuvir
C3858051|ledipasvir-sofosbuvir
C3858051|LEDIPASVIR/SOFOSBUVIR
C3858051|ledipasvir + sofosbuvir
C3858051|antiviral ledipasvir + sofosbuvir
C3858051|ledipasvir + sofosbuvir (medication)
C3858051|ledipasvir, sofosbuvir drug combination
C3858051|ledipasvir - sofosbuvir
C3858051|Ledipasvir + sofosbuvir (product)
C3696724|sofosbuvir Oral Product
C3696724|Oral form sofosbuvir
C3696724|Oral form sofosbuvir (product)
C3857383|ledipasvir 90 MG / sofosbuvir 400 MG Oral Tablet [Harvoni]
C3857383|LEDIPASVIR 90 mg / SOFOSBUVIR 400 mg ORAL TABLET, FILM COATED [Harvoni]
C3857383|Harvoni 90 MG / 400 MG Oral Tablet
C3857383|Harvoni (ledipasvir 90 MG / sofosbuvir 400 MG) Oral Tablet
C3857383|Harvoni 90mg-400mg Tablet
C3857383|Ledipasvir/Sofosbuvir 90 MG-400 MG Oral Tablet [HARVONI]
C3857383|Harvoni, 90 mg-400 mg oral tablet
C3857383|LEDIPASVIR 90 mg / SOFOSBUVIR 400 mg ORAL TABLET, FILM COATED [Harvoni Access]
C3858162|ledipasvir / sofosbuvir Oral Tablet [Harvoni]
C3852670|ombitasvir
C3852670|Ombitasvir (substance)
C3852670|Ombitasvir (product)
C3883273|OMBITASVIR HEMINONAHYDRATE
C4075325|Oral form ombitasvir
C4075325|Oral form ombitasvir (product)
C4080052|elbasvir
C3252090|daclatasvir
C3252090|DCV
C3252090|Daclatasvir (substance)
C3252090|daclatasvir (medication)
C3252090|antiviral daclatasvir
C3252090|Daclatasvir (product)
C3892852|daclatasvir dihydrochloride
C3892852|daclatasvir (as dihydrochloride)
C4046850|Daklinza
C4047230|daclatasvir Oral Product
C4047230|Oral form daclatasvir
C4047230|Oral form daclatasvir (product)
C4047078|Daklinza Pill
C3857361|Daclatasvir 30 MG Oral Tablet
C3857361|DACLATASVIR DIHYDROCHLORIDE 30 mg ORAL TABLET
C3857361|daclatasvir (as daclatasvir dihydrochloride 33 mg) 30 MG Oral Tablet
C3857361|Daclatasvir 30mg Oral tablet
C3857361|DACLATASVIR 30MG TAB
C3857361|Daclatasvir Dihydrochloride Tab 30 MG (Base Equivalent)
C3857361|DACLATASVIR 30MG TAB [VA Product]
C4047197|daclatasvir Oral Tablet
C3892515|DACLATASVIR DIHYDROCHLORIDE 60 mg ORAL TABLET
C3892515|daclatasvir 60 MG Oral Tablet
C3892515|Daclatasvir 60mg Oral tablet
C3892515|daclatasvir (as daclatasvir dihydrochloride 66 mg) 60 MG Oral Tablet
C3892515|DACLATASVIR 60MG TAB
C3892515|Daclatasvir Dihydrochloride Tab 60 MG (Base Equivalent)
C3892515|DACLATASVIR 60MG TAB [VA Product]
C3852655|GS-5885
C3851350|ledipasvir
C3851350|Ledipasvir (substance)
C3851350|Ledipasvir (product)
C4075037|Oral form ledipasvir (product)
C4075037|Oral form ledipasvir
C3858322|ledipasvir / sofosbuvir Oral Product
C3858322|Oral form ledipasvir + sofosbuvir
C3858322|Oral form ledipasvir + sofosbuvir (product)
C3858113|ledipasvir 90 MG / sofosbuvir 400 MG [Harvoni]
C3858080|ledipasvir 90 MG / sofosbuvir 400 MG Oral Tablet
C3858080|Ledipasvir, Sofosbuvir 90-400mg Oral tablet
C3858080|Ledipasvir-Sofosbuvir Tab 90-400 MG
C3858080|ledipasvir-sofosbuvir 90 mg-400 mg oral tablet
C3858080|Ledipasvir/Sofosbuvir 90 MG-400 MG Oral Tablet
C3858080|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB
C3858080|LEDIPASVIR 90MG/SOFOSBUVIR 400MG TAB [VA Product]
C3858300|ledipasvir / sofosbuvir Oral Tablet
C3858199|Harvoni Pill
C3858200|Harvoni Oral Product
