C0201916|Bilirubin, direct measurement
C0236556|Direct reacting bilirubin
C1883011|Serum Direct Bilirubin Measurement
C1883011|serum direct bilirubin measurement (lab test)
C0428439|Conjugated bilirubin level
C0428439|Conjugated bilirubin level (procedure)
C1278035|Plasma conjugated bilirubin level
C1278035|Plasma conjugated bilirubin level (procedure)
C1278035|Plasma conjugated bilirubin measurement (procedure)
C1278035|Plasma conjugated bilirubin measurement
C1278038|Serum conjugated bilirubin level
C1278038|Serum conjugated bilirubin level (procedure)
C1278038|Serum Direct (Conjugated) Bilirubin Test
C1278038|Serum conjugated bilirubin measurement (procedure)
C1278038|Serum conjugated bilirubin measurement
C0580935|Serum conjugated:total bilirubin ratio (& level)
C0580935|Serum conjugated:total bilirubin ratio (& level) (procedure)
C0580935|Se conj total bilirubin ratio
C0580935|Serum conjugated:total bilirubin ratio
C0580935|Serum conjugated/total bilirubin ratio
C0580935|Serum conjugated/total bilirubin ratio measurement (procedure)
C0580935|Serum conjugated/total bilirubin ratio measurement
C0006678|Bilirubinate, Calcium
C0006678|Calcium bilirubinate
C0006678|Salt Bilirubin, Calcium
C0006678|Calcium Salt Bilirubin
C0006678|Bilirubin, Calcium Salt
C0006678|Calcium bilirubinate (substance)
C0053592|21H-biline-8,12-dipropanoic acid, 2,17-diethenyl-1,10-19,22,23,24-hexahydro-3,7,13,18-tetramethyl-1,19-dioxo-, mono-beta-D-glucopyranuronosyl ester
C0053592|bilirubin glucuronate
C0053592|bilirubin glucuronide
C0053592|bilirubin, glucuronic acid conjugates
C0053592|Bilirubin glucuronide (substance)
