C0021682|Health Insurance
C0018717|Medicare
C0018717|Medicare coverage
C3530230|Private health insurance
C3530230|Private health insurance--other commercial Indemnity
C4069202|Private Insurance (includes "no-fault", BCBS, United Health, etc)
C2347682|Private Health Insurance
C1955981|Blue Cross Blue Shield
C1955981|Blue Cross Blue Shield Insurance
C1955981|Blue Cross Blue Shield Insurance Plans
C0005864|Blue Cross
C0021681|Insurance, Dental
C0021681|dental health insurance
C0021681|INSURANCE DENT
C0021681|DENT INSURANCE
C0021681|Dental insurance
C0596896|Medicare/Medicaid
C0018717|Medicare
C0018717|HEALTH INSURANCE AGED DISABLED
C0018717|HEALTH INSURANCE AGED DISABLED TITLE 18
C0018717|HEALTH INSURANCE AGED TITLE 18
C0018717|Medicare Program
C0018717|Medicare coverage (finding)
C0018717|Medicare coverage
C0018717|Health Insurance for Aged, Disabled, Title 18
C0018717|Health Insurance for Aged, Title 18
C0018717|Health Insurance for Aged and Disabled, Title 18
C0018720|Health Maintenance Organizations
C0018720|HMO
C0018720|Organization, Health Maintenance
C0018720|health maintenance organization
C0018720|GROUP HEALTH ORGAN PREPAID
C0018720|ORGAN HEALTH MAINTENANCE
C0018720|HEALTH MAINTENANCE ORGAN
C0018720|PREPAID GROUP HEALTH ORGAN
C0018720|Organizations, Health Maintenance
C0018720|Prepaid Group Health Organizations
C0018720|Group Health Organizations, Prepaid
C0018720|Prepaid healthcare organization
C0018720|Health maintenance organisation
C0018720|Health maintenance organization (environment)
C0018720|Prepaid healthcare organisation
C0021684|Health Insurance Reimbursements
C0021684|Insurance Reimbursement, Health
C0021684|Insurance Reimbursements, Health
C0021684|Insurance, Health, Reimbursement
C0021684|Payment, Third-Party
C0021684|Payments, Third-Party
C0021684|Reimbursements, Health Insurance
C0021684|Third Party Payments
C0021684|Third-Party Payment
C0021684|Health Insurance Reimbursement
C0021684|Third-Party Payments
C0021684|Reimbursement, Health Insurance
C0021684|Third Party Payment
C0021694|Insurance, Psychiatric
C0021694|Insurances, Psychiatric
C0021694|Psychiatric Insurance
C0021694|Psychiatric Insurances
C0021694|Mental health insurance
C0025071|Medicaid
C0025071|Medicaid Program
C0025071|Medicaid coverage (finding)
C0025071|Medicaid coverage
C0042613|Claim, Veterans Disability
C0042613|Claims, Veterans Disability
C0042613|Disability Claim, Veterans
C0042613|Disability Claims, Veterans
C0042613|Veterans Disability Claim
C0042613|Veterans Disability Claims
C0043233|Compensation, Workman's
C0043233|Compensation, Workmen's
C0043233|Compensations, Workman's
C0043233|Compensations, Workmen's
C0043233|Workman Compensation
C0043233|Workman's Compensations
C0043233|Workmans Compensation
C0043233|Workmen Compensation
C0043233|Workmen's Compensations
C0043233|Workmens Compensation
C0043233|Workers' Compensation
C0043233|Compensation, Worker's
C0043233|Compensation, Workers'
C0043233|Compensations, Worker's
C0043233|Compensations, Workers'
C0043233|Worker Compensation
C0043233|Worker's Compensations
C0043233|Workers Compensation
C0043233|Workers' Compensations
C0043233|workmen's compensation
C0043233|Workers Compensation Plan
C0043233|Worker's Compensation
C0043233|Workman's Compensation
C0242816|Fee for Service Plans
C0242816|Fee for Services
C0242816|Fee-for-Service Plan
C0242816|Fee-for-Service Plans
C0242816|Fees for Services
C0242816|Plan, Fee-for-Service
C0242816|Plans, Fee-for-Service
C0242816|Service, Fee for
C0242816|Service, Fees for
C0242816|Services, Fee for
C0242816|Services, Fees for
C0242816|FEE SERV
C0242816|Fee for Service Payment Method
C0242816|Fee-for-Service
C0242816|Fee for Service
C0242816|FFS
C0242816|Fees for Service
C0242816|Fee for Service payment plan
C0681104|Employee Health Insurance
C0086599|MED ASSISTANCE TITLE 19
C0086599|Medical Assistance, Title 19
C0021680|Accident Insurances
C0021680|Insurance, Accident
C0021680|Insurances, Accident
C0021680|Accident insurance
C0021685|Insurance, Hospitalization
C0021685|Hospitalization insurance
C0024679|Managed Care Program
C0024679|Managed Care Programs
C0024679|Program, Managed Care
C0024679|Programs, Managed Care
C0024679|Managed Health Care Insurance Plans
C0085563|Health Plan, Prepaid
C0085563|Plan, Prepaid Health
C0085563|Plans, Prepaid Health
C0085563|Prepaid Health Plan
C0085563|Prepaid Health Plans
C0085563|Health Plans, Prepaid
C0282485|Managed Competition
C0282485|Competition, Managed
C0600593|PUBLIC LAW 104 191
C0600593|PL 104 191
C0600593|Kassebaum Kennedy Act
C0600593|PL 104-191
C0600593|HIPAA
C0600593|Public Law 104-191
C0600593|United States Health Insurance Portability and Accountability Act
C0600593|Health Insurance Portability and Accountability Act
C0600593|PL104 191
C0600593|Kennedy Kassebaum Act
C0600593|PL104-191
C0021682|Insurance, Health
C0021682|health insurance
C0018688|Health Benefit Plans, Employee
C0018688|Employee Health Benefit Plans
C0021688|Insurance, Long Term Care
C0021688|Insurance, Long-Term Care
C0021688|Long Term Care Insurance
C0021688|Long-term Care Insurance
C0021690|Insurance, Nursing Services
C0021690|Insurances, Nursing Services
C0021690|Nursing Services Insurances
C0021690|Services Insurance, Nursing
C0021690|Services Insurances, Nursing
C0021690|INSURANCE NURS SERV
C0021690|NURS SERV INSURANCE
C0021690|Nursing Services Insurance
C0021691|Insurance, Pharmaceutical Services
C0021691|PHARM SERV INSURANCE
C0021691|INSURANCE PHARM SERV
C0021691|Pharmaceutical services insurance
C0021691|Insurance, Pharmacy Services
C0021691|Pharmacy Services Insurance
C0021691|Insurance, Pharmaceutic Services
C0021691|Pharmaceutic Services Insurance
C0085558|Insurance, Medigap
C0085558|Medigap Policies
C0085558|Policies, Medigap
C0085558|Policy, Medigap
C0085558|Medigap Insurance
C0085558|Medigap Policy
C0600588|SAVINGS ACCOUNTS MED
C0600588|ACCOUNTS MED SAVINGS
C0600588|MED SAVINGS ACCOUNTS
C0600588|Account, Medical Savings
C0600588|Medical Savings Account
C0600588|Medical Savings Accounts
C0600588|Savings Account, Medical
C0600588|Accounts, Medical Savings
C0600588|Savings Accounts, Medical
C0021689|Insurance, Major Medical
C0021689|INSURANCE MAJOR MED
C0021689|MAJOR MED INSURANCE
C0021689|MED INSURANCE MAJOR
C0021689|Medical Insurance, Major
C0021689|Major Medical Insurance
C0021693|Insurance, Physician Services
C0021693|Insurances, Physician Services
C0021693|Physician Services Insurance
C0021693|Physician Services Insurances
C0021693|Services Insurances, Physician
C0021693|Insurance Physician Service
C0021693|Insurance Physician Services
C0021693|Physician Service, Insurance
C0021693|Service, Insurance Physician
C0021693|Services, Insurance Physician
C0021693|INSURANCE PHYSICIAN SERV
C0021693|SERV INSURANCE PHYSICIAN
C0021693|PHYSICIAN SERV INSURANCE
C0021693|Services Insurance, Physician
C0021693|Physician Services, Insurance
C0021695|Insurance, Surgical
C0021695|Insurances, Surgical
C0021695|Surgical Insurances
C0021695|INSURANCE SURG
C0021695|SURG INSURANCE
C0021695|Surgical Insurance
C0027454|National Health Insurance, United States
C0027454|NATL HEALTH INSUR US
C0027454|National health insurance--United States
C0027454|United States National Health Insurance
C0027454|Federal Health Insurance Plans, United States
C0282487|Single Payer System
C0282487|Single-Payer System
C0282487|Single-Payer Systems
C0282487|System, Single-Payer
C0282487|Systems, Single-Payer
C0018256|Health Insurance, Group
C0018256|Insurance, Group Health
C0018256|Group Health Insurance
C0018718|Insurance, Voluntary Health
C0018718|Voluntary Health Insurance
C0018718|Health Insurance, Voluntary
C2936611|PL111 148
C2936611|111-148, PL
C2936611|Public Law 111 148
C2936611|Patient Protection and Affordable Care Act
C2936611|PL 111 148
C2936611|Care Act, Affordable (ACA)
C2936611|Acts, Affordable Care (ACA)
C2936611|Care Act, Affordable
C2936611|Acts, Affordable Care
C2936611|Act, Affordable Care
C2936611|Affordable Care Acts
C2936611|Care Acts, Affordable
C2936611|Affordable Care Act
C2936611|PL 111-148
C2936611|Obamacare
C2936611|Public Law 111-148
C2936611|Affordable Care Act (ACA)
C2936611|Health Care Reform Act
C2936611|PL111-148
C2936638|For Profit Insurance Plans
C2936638|Insurance Plans, For-Profit
C2936638|Insurance Plan, For-Profit
C2936638|For-Profit Insurance Plan
C2936638|Plans, For-Profit Insurance
C2936638|For-Profit Insurance Plans
C2936639|Plans, Not-For-Profit Insurance
C2936639|Not-For-Profit Insurance Plan
C2936639|Not-For-Profit Insurance Plans
C2936639|Insurance Plan, Not-For-Profit
C2936639|Insurance Plans, Not-For-Profit
C2936639|Plan, Not-For-Profit Insurance
C2936639|Not For Profit Insurance Plans
C2347682|Private Health Insurance
C2347682|Health Insurance
C3494321|Purchasings, Value-Based
C3494321|Value-Based Purchasing
C3494321|Value Based Purchasing
C3494321|Value-Based Purchasings
C3494321|Purchasing, Value-Based
C4042889|Children's Health Insurance Program
C0079817|Medicare Part A
C0079817|Part A, Medicare
C0079817|MEDICARE HOSP INSURANCE PROGRAM
C0079817|MEDICARE A
C0079817|HOSP INSURANCE PROGRAM MEDICARE
C0079817|Hospital Insurance Program, Medicare
C0079817|Medicare Hospital Insurance Program
C0079818|Medicare Part B
C0079818|Part B, Medicare
C0079818|Program, SMI
C0079818|Programs, SMI
C0079818|SMI Programs
C0079818|MEDICARE SUPPLEMENTARY MED INSURANCE PROGRAM
C0079818|MEDICARE B
C0079818|SUPPLEMENTARY MED INSURANCE PROGRAM MEDICARE
C0079818|Supplementary Medical Insurance Program, Medicare
C0079818|SMI Program
C0079818|Medicare Supplementary Medical Insurance Program
C0025114|Assignment, Medicare
C0025114|Assignments, Medicare
C0025114|Medicare Assignment
C0025114|Medicare Assignments
C0600580|MEDICARE C
C0600580|Medicare Part C
C0600580|Part C, Medicare
C0600580|Choice, Medicare Plus
C0600580|Plus Choice, Medicare
C0600580|Programs, Medicare+Choice (US)
C0600580|Medicare+Choice Programs (US)
C0600580|Program, Medicare+Choice (US)
C0600580|Medicare+Choice Program (US)
C0600580|Medicare Plus Choice Program (US)
C0600580|Medicare Choice
C0600580|Medicare Plus Choice
C1955953|Medicare Part D
C1955953|Part D, Medicare
C3530305|Medicare (Managed Care)
C3530300|Medicare (Non-managed Care)
C3530295|Medicare Other
C3530238|Managed Care (Private)
C3530234|Private Health Insurance - Indemnity
C3530229|Managed Care (private) or private health insurance (indemnity), not otherwise specified
C3530228|Organized Delivery System
C3530227|Small Employer Purchasing Group
C3530226|Other Private Insurance
C1955981|Blue Cross Blue Shield Insurance Plans
C1955981|BLUE CROSS/BLUE SHIELD
C0005864|Blue Cross
C0005864|Blue Crosses
C0005864|Cross, Blue
C0005864|Crosses, Blue
C0005865|Shields, Blue
C0005865|Shield, Blue
C0005865|Blue Shield
C0005865|Blue Shields
C3530225|BC Managed Care
C3530220|BC Indemnity
C3530219|BC (Indemnity or Managed Care) - Out of State
C3530218|BC (Indemnity or Managed Care) - Unspecified
C3530217|BC (Indemnity or Managed Care) - Other
