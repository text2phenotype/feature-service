C1990758|INR platelet poor plasma
C0005790|Blood coagulation tests
C0525032|International Normalized Ratio
C0525032|INR
C0525032|LOINC LP20762-8
C0525032|LOINC 20762-8
C2360882|Coagulation tissue factor induced.INR^post heparin adsorption:RelTime:Pt:PPP:Qn:Coag
C2360882|INR in Platelet poor plasma by Coagulation assay --post heparin adsorption
C2360882|INR p heparin adsorption PPP
C2360882|Coagulation tissue factor induced.INR^post heparin adsorption:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482691|INR in Platelet poor plasma by Coagulation assay
C0482691|INR PPP
C0482691|Coagulation tissue factor induced.INR:RelTime:Pt:PPP:Qn:Coag
C0482691|Coagulation tissue factor induced.INR:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0033707|Prothrombin Time
C0033707|Prothrombin Times
C0033707|Time, Prothrombin
C0033707|Times, Prothrombin
C0033707|Prothrombin time (PT)
C0033707|PT
C0033707|Prothrombin Time Test
C0033707|prothrombin time (PT) (lab test)
C0033707|Test;prothrombin time
C0033707|Prothrombin time assay
C0033707|PT assay
C0033707|Protime
C0033707|PTT - Prothrombin time
C0033707|Quick one stage prothrombin time
C0033707|PT - Prothrombin time
C0033707|Prothrombin time (procedure)
C0033707|One stage prothrombin time
C0033707|One stage prothrombin time (procedure)
C0033707|Pro-thrombin time
C0033707|Prothrombin test
C0033707|Plasma Prothrombin Test
C0005729|Bleeding Time
C0005729|Bleeding Times
C0005729|Time, Bleeding
C0005729|Times, Bleeding
C0005729|bleeding time (lab test)
C0005729|Test;bleeding time
C0005729|BLEEDING TIME TEST
C0005729|Measurement of bleeding time
C0005729|Bleeding time (finding)
C0005729|BLEEDT
C0005729|Clotting Time Homeostasis
C0005729|Bleeding time (procedure)
C0005729|Bleeding time - observation
C0005729|Bleeding time procedure
C0005729|Bleeding time, NOS
C0005729|test bleeding time
C0040017|Thrombelastography
C0040017|THROMBELASTOGR
C0040017|THROMBOELASTOGR
C0040017|thromboelastography (lab test)
C0040017|thromboelastography
C0040017|Thromboelastogram
C0040017|Thromboelastography (procedure)
C0043159|Whole Blood Coagulation Time
C0043159|Coagulation time; Lee and White
C0043159|ACTIVATED COAG TIME WHOLE BLOOD
C0043159|WHOLE BLOOD COAG TIME
C0043159|BLOOD COAG TIME WHOLE
C0043159|COAG TIME WHOLE BLOOD
C0043159|COAGULATION TIME LEE AND WHITE
C0043159|COAGULATION TIME LEE & WHITE
C0043159|Lee and White coagulation time test
C0043159|Whole blood clotting time (procedure)
C0043159|Whole blood clotting time
C0043159|whole blood clotting time (lab test)
C0043159|Activated Coagulation Time, Whole Blood
C0043159|Coagulation Time, Whole Blood
C0043159|Blood Coagulation Time, Whole
C0043159|Coagulation time, Lee White
C0043159|Lee White coagulation time
C0043159|Blood coagulation time
C0043159|WBCT - Whole blood clotting time
C0043159|Coagulation time, Lee White (procedure)
C0043159|Whole blood clotting time procedure (procedure)
C0043159|Whole blood clotting time procedure
C1255157|Sonoclot Coagulation Rate Test
C1255158|Sonoclot Peak Time Test
C1255159|Whole Blood Clot Onset Time Test
C0005790|Blood Coagulation Test
C0005790|Blood Coagulation Tests
C0005790|Coagulation Test, Blood
C0005790|Test, Blood Coagulation
C0005790|coagulation studies
C0005790|TESTS BLOOD COAG
C0005790|BLOOD COAG TESTS
C0005790|COAG TESTS BLOOD
C0005790|Coagulation Study
C0005790|Coagulation
C0005790|Coag
C0005790|Clotting screening
C0005790|Blood coagulation test (procedure)
C0005790|Clotting screening (procedure)
C0005790|Clotting
C0005790|Coagulation Tests, Blood
C0005790|Tests, Blood Coagulation
C0005790|Bleeding Time Test
C0005790|Clotting screen
C0005790|Coagulation system screening
C0005790|Blood coagulation panel (procedure)
C0005790|Blood coagulation panel
C0005790|Blood coagulation screen
C0005790|Blood coagulation panel, NOS
C0005790|Blood coagulation screen, NOS
C0030605|APTT
C0030605|PTT
C0030605|partial thromboplastin time: PTT
C0030605|Partial Thromboplastin Time
C0030605|Activated partial thromboplastin time
C0030605|partial thromboplastin time (PTT) (lab test)
C0030605|partial thromboplastin time (PTT)
C0030605|activated PTT
C0030605|activated partial thromboplastin time (aPTT)
C0030605|activated partial thromboplastin time (aPTT) (lab test)
C0030605|Partial thromboplastin time activated
C0030605|Activated partial thromboplastin time (procedure)
C0030605|Partial thromboplastin time activated (procedure)
C0030605|Thromboplastin time, partial (PTT)
C0030605|Thromboplastin Time, Partial
C0030605|Plasma Thromboplastin Test
C0030605|Partial thromboplastin time, activated
C0030605|PTT, activated
C0030605|PTT assay
C0030605|APTT - Activated partial thromboplastin time
C0030605|PTT - Partial thromboplastin time
C0030605|Partial thromboplastin time, activated (procedure)
C0030605|Activated Partial Thromboplastin Time measurement
C0677634|Reptilase Times
C0677634|Thrombin Time
C0677634|Thrombin Times
C0677634|Time, Reptilase
C0677634|Time, Thrombin
C0677634|Times, Reptilase
C0677634|Times, Thrombin
C0677634|Thrombin time; plasma
C0677634|TCT
C0677634|thrombin clotting time
C0677634|reptilase time
C0677634|reptilase time (lab test)
C0677634|Thrombin Time Assay
C0677634|thrombin time (lab test)
C0677634|reptilase time test
C0677634|TT
C0677634|THROMBIN TIME PLASMA
C0677634|Test;thrombin time
C0677634|Thrombin time test on plasma
C0677634|Reptilase clotting time (procedure)
C0677634|Reptilase clotting time
C0677634|Thrombin time (procedure)
C0677634|Plasma Thrombin Test
C0677634|Fibrin time
C0677634|TT - Thrombin time
C0677634|Reptilase time (procedure)
C0677634|Thrombin time - observation
C0677634|thrombin time test
C0525032|International Normalized Ratio
C0525032|International Normalized Ratios
C0525032|Normalized Ratio, International
C0525032|Normalized Ratios, International
C0525032|Ratio, International Normalized
C0525032|Ratios, International Normalized
C0525032|INR
C0525032|international normalized ratio (INR)
C0525032|international normalized ratio (INR) (lab test)
C0525032|International normalised ratio
C0525032|BCR
C0525032|coagulation studies: INR
C0525032|International normalised ratio (procedure)
C0525032|Prothrombin Intl. Normalized Ratio
C0525032|INR (International normalised ratio)
C0525032|INR (International normalized ratio)
C0525032|International normalized ratio (qualifier value)
C0525032|INR - Internationalised ratio
C0525032|Internationalised ratio
C0525032|International normalized ratio (observable entity)
C0525032|INR - Internationalized ratio
C0525032|Internationalized ratio
C0200416|Antithrombin III
C0200416|antithrombin III assay (lab test)
C0200416|antithrombin III assay
C0200416|Antithrombin III Measurement
C0200416|Antithrombin Activity Measurement
C0200416|Antithrombin III level
C0200416|Antithrombin III level (procedure)
C0200416|Antithrombin
C0200416|Antithrombin III Activity
C0200416|Antithrombin Activity
C0200416|ANTHRM
C0200416|Antithrombin III assay (procedure)
C0200416|Antithrombin III assay, NOS
C2825855|Factor III Measurement
C2825855|Tissue Factor, CD142
C2825855|Factor III
C2825855|FACTIII
C2825856|Factor VII Measurement
C2825856|FACTVII
C2825856|Stable Factor
C2825856|Factor VII
C2825856|Proconvertin
C2825857|Factor VIII Measurement
C2825857|Factor VIII
C2825857|FACTVIII
C2825857|Anti-hemophilic Factor
C3274375|Anti-Factor Xa Activity Measurement
C3274375|Anti-Factor Xa Activity
C3274375|AFACTXAA
C0200408|factor IX assay
C0200408|factor IX assay (lab test)
C0200408|factor IX level
C0200408|Coagulation factor IX level
C0200408|Clotting; factor IX (PTC or Christmas)
C0200408|Coagulation factor IX measurement
C0200408|CLOTTING FACTOR IX PTC/CHRISTMAS
C0200408|Factor IX Measurement
C0200408|CLOT FACTOR IX PTC/CHRSTMAS
C0200408|Assay for clotting factor IX (PTC)
C0200408|Clotting factor IX (PTC or Christmas) measurement
C0200408|Factor IX assay (procedure)
C0200408|Christmas Factor
C0200408|Factor IX
C0200408|FACTIX
C0200408|Clotting factor IX assay
C0200408|Christmas disease factor assay
C0200408|Hemophilia B assay
C0200408|Plasma thromboplastin component assay
C0200408|Haemophilia B assay
C0200408|Clotting factor IX assay (procedure)
C0200408|Autoprothrombin II assay
C3274393|Factor V Measurement
C3274393|Factor V
C3274393|FACTV
C3274393|Labile Factor
C3274394|Factor X Measurement
C3274394|Factor X
C3274394|FACTX
C3274435|Prothrombin Activity Measurement
C3274435|Factor II Activity
C3274435|Prothrombin Activity
C3274435|PTA
C2239219|von Willebrand's factor (lab test)
C2239219|von Willebrand Factor Measurement
C2239219|Clotting factor VIII (von Willebrand factor) measurement
C2239219|von Willebrand Factor
C2239219|von Willebrand Factor Antigen
C2239219|FACTVW
C2239219|von Willebrand factor (lab test)
C2239219|von Willebrand's factor
C3640656|Endogenous Thrombin Potential Measurement
C3640656|Endogenous Thrombin Potential
C3640656|ETP
C3272912|Reptilase Time Measurement
C3272912|Reptilase Time
C3272912|RPTLTIME
C3640663|Lupus Anticoagulant Sensitive APTT Measurement
C3640663|Lupus Anticoagulant Sensitive APTT
C3640663|APTTLAS
C3640663|APTT-LA
C3541350|Factor V Activity Measurement
C3541350|FACTVA
C3541350|Factor V Activity
C3541350|Labile Factor Activity
C3640659|Endogenous Thrombin Potential Time to Peak Measurement
C3640659|ETP Time to Peak
C3640659|Endogenous Thrombin Potential Time to Peak
C3640659|ETPTP
C3641237|Dilute Russell's Viper Venom Time to Control Ratio Measurement
C3641237|DRVVTRT
C3641237|Lupus Anticoagulant Ratio
C3641237|Dilute Russell's Viper Venom Time Ratio
C3640654|Endogenous Thrombin Potential Lag Time Measurement
C3640654|Endogenous Thrombin Potential Lag Time
C3640654|ETPLT
C3640654|ETP Lag Time
C3641245|Factor VIIa Activity Measurement
C3641245|Factor VIIa Activity
C3641245|FCTVIIAA
C3641244|Factor VII Activity Measurement
C3641244|FACTVIIA
C3641244|Stable Factor Activity
C3641244|Proconvertin Activity
C3641244|Factor VII Activity
C0427611|Coagulation time; activated
C0427611|clotting time, activated
C0427611|activated clotting time (lab test)
C0427611|activated clotting time
C0427611|activated coagulation time
C0427611|COAGULATION TIME ACTIVATED
C0427611|Activated coagulation time test
C0427611|ACT
C0427611|ACT - activated clotting time
C0427611|Activated Clot Time
C0427611|Coagulation Activated
C0427611|Coagulation time, activated
C0427611|Ground glass clotting time
C0427611|Whole blood activated clotting time
C0427611|Coagulation time, activated (procedure)
C0427611|Activated clotting time measurement
C3640660|Endogenous Thrombin Potential Time to Peak Relative Measurement
C3640660|ETP Time to Peak Relative
C3640660|Endogenous Thrombin Potential Time to Peak Relative
C3640660|ETPTPR
C3640653|Endogenous Thrombin Potential Area Under Curve Measurement
C3640653|Endogenous Thrombin Potential Area Under Curve
C3640653|ETPAUC
C3640653|ETP Area Under Curve
C3641246|Factor VIII Activity Measurement
C3641246|Factor VIII Activity
C3641246|Anti-hemophilic Factor Activity
C3641246|FCTVIIIA
C3542419|Factor V Leiden Measurement
C3542419|FACTVL
C3542419|Factor V Leiden
C2199618|ecarin clotting time
C2199618|ecarin clotting time (lab test)
C2199618|clotting time, ecarin
C2199618|Ecarin Clotting Time Measurement
C2199618|ECT
C0920267|platelet aggregation
C0920267|platelet aggregation (lab test)
C0920267|Platelet aggr
C0920267|Platelet aggregation measurement
C0920267|Platelet aggregation test (procedure)
C0920267|Platelet aggregation assay (qualifier value)
C0920267|Platelet aggregation assay
C0920267|Platelet aggregation test
C0920267|PLATAGGR
C0920267|Platelet Function
C0920267|Platelet aggregation NOS
C0920267|Aggregometer test
C0920267|Platelet aggregation test, NOS
C0920267|Aggregometer test, NOS
C3640658|Endogenous Thrombin Potential Peak Height Relative Measurement
C3640658|ETP Peak Height Relative
C3640658|ETPPHR
C3640658|Endogenous Thrombin Potential Peak Height Relative
C3640655|Endogenous Thrombin Potential Lag Time Relative Measurement
C3640655|ETP Lag Time Relative
C3640655|ETPLTR
C3640655|Endogenous Thrombin Potential Lag Time Relative
C3642159|Factor XIV Activity Measurement
C3642159|Factor XIV Activity
C3642159|Protein C Function
C3642159|FACTXIVA
C3642159|Protein C Activity
C1168438|Protein C Measurement
C1168438|Factor XIV Measurement
C1168438|Autoprothrombin IIA
C1168438|Protein C Antigen
C1168438|FACTXIV
C1168438|Protein C
C1168438|Factor XIV
C1168438|Protein C antigen measurement
C3640657|Endogenous Thrombin Potential Peak Height Measurement
C3640657|ETP Peak Height
C3640657|ETPPH
C3640657|Endogenous Thrombin Potential Peak Height
C3538955|Factor IX Activity Measurement
C3538955|Christmas Factor Activity Measurement
C3538955|Factor IX Activity
C3538955|Christmas Factor Activity
C3538955|FACTIXA
C1271595|Other coagulation/bleeding tests (procedure)
C1271595|Other coagulation/bleeding tests
C0364172|Cardiolipin [Mass/volume] in Serum
C0364172|Cardiolipin Ser-mCnc
C0364172|Cardiolipin:MCnc:Pt:Ser:Qn
C0364172|Cardiolipin:Mass Concentration:Point in time:Serum:Quantitative
C0945541|Prot S Act/Nor PPP
C0945541|Protein S actual/normal in Platelet poor plasma by Coagulation assay
C0945541|Protein S actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0945541|Protein S actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0943668|von Willebrand factor Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C0943668|von Willebrand factor Ag:ACnc:Pt:PPP:Qn:EIA
C0943668|Deprecated vWF Ag PPP EIA-aCnc
C0943668|Deprecated von Willebrand factor (vWf) Ag [Units/volume] in Platelet poor plasma by EIA
C0945642|Plasminogen actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C0945642|Plasminogen actual/normal in Platelet poor plasma by Chromogenic method
C0945642|PLG Act/Nor PPP Chro
C0945642|Plasminogen actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0365431|Fibrin.soluble:ACnc:Pt:Ser:Qn:Coag
C0365431|Fibrin Sol Ser-aCnc
C0365431|Fibrin.soluble [Units/volume] in Serum by Coagulation assay
C0365431|Fibrin.soluble:Arbitrary Concentration:Point in time:Serum:Quantitative:Coagulation Assay
C0482705|Fibrinogen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:COAGULATION ASSAY
C0482705|Fibrinogen PPP-mCnc
C0482705|Fibrinogen [Mass/volume] in Platelet poor plasma by Coagulation assay
C0482705|Fibrinogen:MCnc:Pt:PPP:Qn:Coag
C1316351|Coagulation surface induced.factor substitution^1H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316351|Coagulation surface induced.factor substitution^1 hour post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316351|aPTT 1h p 1:4 NP Cont PPP
C1316351|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --1H post incubation with 1:4 normal plasma
C1316353|Coagulation surface induced.factor substitution^2H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1316353|Coagulation surface induced.factor substitution^2 hours post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1316353|aPTT 2h NP PPP
C1316353|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --2H post incubation with normal plasma
C1316354|Coagulation surface induced.factor substitution^2H post incubation after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316354|Coagulation surface induced.factor substitution^2 hours post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316354|aPTT 2h NP Cont PPP
C1316354|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --2H post incubation with normal plasma
C0482711|Fibrinopeptide B beta (1-42) Ag:MCnc:Pt:PPP:Qn:Imm
C0482711|FpB Beta1-42 Ag PPP Imm-mCnc
C0482711|Fibrinopeptide B beta (1-42) Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482711|Fibrinopeptide B beta (1-42) Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1315990|PA Coll lo dose PRP
C1315990|Platelet aggregation.collagen induced^low dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1315990|Platelet aggregation.collagen induced^low dose:RelACnc:Pt:PRP:Qn
C1315990|Platelet aggregation collagen induced in Platelet rich plasma --Low dose
C0482605|Antithrombin Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482605|Antithrombin Ag:ACnc:Pt:PPP:Qn:Imm
C0482605|AT III Ag PPP Imm-aCnc
C0482605|Antithrombin Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1147716|Phosphatidylserine IgG Ab [Units/volume] in Serum by Immunoassay
C1147716|Phosphatidylserine Ab.IgG:ACnc:Pt:Ser:Qn:EIA
C1147716|PS IgG Ser EIA-aCnc
C1147716|Phosphatidylserine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0482636|Coagulation factor VIII Activity.Xa activator [Units/volume] in Platelet poor plasma by Chromogenic method
C0482636|Coagulation factor VIII activity.X(little a) activator:ACnc:Pt:PPP:Qn:Chromo
C0482636|Fact VIII Xa Act PPP Chro-aCnc
C0482636|Coagulation factor VIII activity.X(a) activator:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1624141|Cardiolipin Ab.IgA.B2GP1 independent:MoM:Pt:Ser:Qn
C1624141|Cardiolipin IgA B2GP1 indep MoM Ser
C1624141|Cardiolipin IgA Ab B2GP1 independent [Multiple of the median] in Serum
C1624141|Cardiolipin Antibody.immunoglobulin A.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C2361182|Clot formation.extrinsic coagulation system activated.fibrinolysis suppressed:Time:Pt:Bld:Qn:Thromboelastography
C2361182|Clot formation.extrinsic coagulation system activated.fibrinolysis suppressed [Time] in Blood by Thromboelastography
C2361182|Clot formation.extrinsic coagulation system activated.fibrinolysis suppressed:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361182|CFT.fibinolysis sup Bld TEG
C1978764|Coagulation surface induced.lupus sensitive.factor substitution^1H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1978764|Coagulation surface induced.lupus sensitive.factor substitution^1 hour post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1978764|aPTT-LA 1h NP PPP
C1978764|aPTT.lupus sensitive.factor substitution in Platelet poor plasma by Coagulation assay --1H post incubation with normal plasma
C1978252|Prothrombin time (PT) circulating inhibitor [Presence] in Platelet poor plasma
C1978252|PTcirculating inhib PPP Ql
C1978252|Coagulation tissue factor induced circulating inhibitor:ACnc:Pt:PPP:Ord
C1978252|Coagulation tissue factor induced circulating inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C0482679|Coagulation surface induced normal/Actual:RelTime:Pt:PPP:Qn:Coag
C0482679|aPTT Inv Ratio PPP
C0482679|Coagulation surface induced normal/Actual:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482679|aPTT normal/actual in Platelet poor plasma by Coagulation assay
C0482669|Deprecated Russell viper venom time in Platelet poor plasma from control by Coagulation assay
C0482669|Coagulation Russell viper venom induced:Time:Pt:PPP^control:Qn:Tilt tube
C0482669|Deprecated Coag RVV Ind PPP Cont Qn
C0482669|Coagulation Russell viper venom induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Tilt tube
C0482677|COAGULATION SURFACE INDUCED.FACTOR SUBSTITUTION^IMMEDIATELY AFTER ADDITION OF NORMAL PLASMA:TIME:POINT IN TIME:PLATELET POOR PLASMA:QUANTITATIVE:COAGULATION ASSAY
C0482677|Deprecated aPTT imm NP PPP Qn
C0482677|Deprecated Activated partial thrombplastin time (aPTT).factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C0482677|Coagulation surface induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C0482677|Deprecated Activated partial thrombplastin time (aPTT).factor substitution in Platelet poor plasma by Coagulation assay --immediately after 1:1 addition of normal plasma
C0482677|aPTT imm NP PPP
C0482677|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C2708583|Hirudin [Mass/volume] in Platelet poor plasma by Chromogenic method
C2708583|Hirudin PPP Chro-mCnc
C2708583|Hirudin:MCnc:Pt:PPP:Qn:Chromo
C2708583|Hirudin:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C2598758|von Willebrand factor cleaving protease actual/normal:RelCCnc:Pt:PPP:Qn:Chromo
C2598758|von Willebrand factor (vWf) cleaving protease actual/normal in Platelet poor plasma by Chromogenic method
C2598758|vWF Cp Act/Nor PPP Chro
C2598758|von Willebrand factor cleaving protease actual/normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3259767|Heparin/kg body weight:Mass Content:Point in time:Whole blood:Quantitative
C3259767|Heparin/kg body weight:MCnt:Pt:Bld:Qn
C3259767|Heparin/kg body weight [Mass/mass] in Blood
C3259767|Heparin/kg BW Bld-mCnt
C3259776|Clot strength:ArEnrg:Pt:Bld:Qn:Thromboelastography
C3259776|Clot strength in Blood by Thromboelastography
C3259776|Clot strength:Energy/Area:Point in time:Whole blood:Quantitative:Thromboelastography
C3259776|Clot strength Bld TEG
C3259338|Clot firmness reduction [Length fraction] in Blood by Thromboelastography --60M post maximum clot amplitude
C3259338|CF reduc 60M p MA LenFr Bld TEG
C3259338|Clot firmness reduction^60M post maximum clot amplitude:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C3259338|Clot firmness reduction^60M post maximum clot amplitude:LenFr:Pt:Bld:Qn:Thromboelastography
C0482745|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex [Mass/volume] in Platelet poor plasma by Immunologic method --10 minutes post venistasis
C0482745|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex^10M post venistasis:MCnc:Pt:PPP:Qn:Imm
C0482745|tPA-PAI1 10M PPP Imm-mCnc
C0482745|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex^10 minutes post venistasis:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0365496|PA Epineph PRP
C0365496|Platelet aggregation.epinephrine induced:RelACnc:Pt:PRP:Qn
C0365496|Platelet aggregation epinephrine induced in Platelet rich plasma
C0365496|Platelet aggregation.epinephrine induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0482774|von Willebrand factor multimers:Prid:Pt:PPP:Nom:IB
C0482774|von Willebrand factor (vWf) multimers in Platelet poor plasma by Immunoblot (IB)
C0482774|vWF multimers PPP IB
C0482774|von Willebrand factor multimers:Presence or Identity:Point in time:Platelet poor plasma:Nominal:Immune Blot
C0484869|Phospholipid Ab [Units/volume] in Serum
C0484869|Phospholipid Ab Ser-aCnc
C0484869|Phospholipid Ab:ACnc:Pt:Ser:Qn
C0484869|Phospholipid Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C1980609|Acarboxyprothrombin &#x7C; Bld-Ser-Plas
C0800003|Fibrinopeptide B beta (43-47) Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0800003|Fibrinopeptide B beta (43-47) Ag:ACnc:Pt:PPP:Qn:Imm
C0800003|FpB Beta43-47 Ag PPP Imm-aCnc
C0800003|Fibrinopeptide B beta (43-47) Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0551336|Phosphatidylglycerol Ab.IgA:ACnc:Pt:Ser:Qn
C0551336|PG IgA Ser-aCnc
C0551336|Phosphatidylglycerol IgA Ab [Units/volume] in Serum
C0551336|Phosphatidylglycerol Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C0802066|Phospholipid Ab:ACnc:Pt:Ser:Ord
C0802066|Phospholipid Ab Ser Ql
C0802066|Phospholipid Ab [Presence] in Serum
C0802066|Phospholipid Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C0943513|Protein C actual/normal in Platelet poor plasma by Chromogenic method
C0943513|Prot C Act/Nor PPP Chro
C0943513|Protein C actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C0943513|Protein C actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0365452|Heparin.unfractionated:MRat:24H:Urine:Qn
C0365452|Heparin unfractionated [Mass/time] in 24 hour Urine
C0365452|Heparin.unfractionated:Mass Rate:24 hours:Urine:Quantitative
C0365452|UFH 24h Ur-mRate
C1316134|Platelet aggregation.collagen induced lag^high dose:Time:Pt:PRP:Qn
C1316134|Platelet aggregation collagen induced lag [Time] in Platelet rich plasma --High dose
C1316134|Platelet aggregation.collagen induced lag^high dose:Time:Point in time:Platelet rich plasma:Quantitative
C1316134|PA Coll Lag time hi dose PRP
C1315987|PA ADP hi dose PRP
C1315987|Platelet aggregation.adenosine diphosphate induced^high dose:RelACnc:Pt:PRP:Qn
C1315987|Platelet aggregation.adenosine diphosphate induced^high dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1315987|Platelet aggregation ADP induced in Platelet rich plasma --High dose
C1146844|Heparin anti Xa:ACnc:Pt:Flu.nonbiological:Qn
C1146844|Heparin Anti Xa Fld.NB-aCnc
C1146844|Heparin anti Xa [Units/volume] in Nonbiological fluid
C1146844|Heparin anti Xa:Arbitrary Concentration:Point in time:Flu.nonbiological:Quantitative
C1625225|PS IgA B2GP1 indep MoM Ser
C1625225|Phosphatidylserine Ab.IgA.B2GP1 independent:MoM:Pt:Ser:Qn
C1625225|Phosphatidylserine IgA Ab B2GP1 independent [Multiple of the median] in Serum
C1625225|Phosphatidylserine Antibody.immunoglobulin A.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1632957|Fibrin D-dimer:ACnc:Pt:CSF:Ord
C1632957|D Dimer CSF Ql
C1632957|Fibrin D-dimer [Presence] in Cerebral spinal fluid
C1632957|Fibrin D-dimer:Arbitrary Concentration:Point in time:Cerebral spinal fluid:Ordinal
C1623602|Cardiolipin Ab.IgA.B2GP1 dependent:MoM:Pt:Ser:Qn
C1623602|Cardiolipin IgA Ab B2GP1 dependent [Multiple of the median] in Serum
C1623602|Cardiolipin IgA B2GP1 dep MoM Ser
C1623602|Cardiolipin Antibody.immunoglobulin A.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C2925953|Fact VIII Ab PPP Ql Imm
C2925953|Coagulation factor VIII Ab [Presence] in Platelet poor plasma by Immunologic method
C2925953|Coagulation factor VIII Ab:ACnc:Pt:PPP:Ord:Imm
C2925953|Coagulation factor VIII Antibody:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Imm
C0482667|Coagulation Russell viper venom induced:Time:Pt:PPP^control:Qn:Coag
C0482667|Coagulation Russell viper venom induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482667|Russell viper venom time in control Platelet poor plasma by Coagulation assay
C0482667|RVV time Cont PPP
C0482676|Coagulation surface induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP^control:Qn:Tilt tube
C0482676|Deprecated Activated partial thrombplastin time (aPTT).factor substitution in Platelet poor plasma from control by Coagulation assay --immediately after addition of normal plasma
C0482676|Deprecated aPTT imm NP PPP Cont Qn
C0482676|Coagulation surface induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Tilt tube
C0482742|Plasminogen activator inhibitor 2 Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482742|PAI2 Ag PPP Imm-mCnc
C0482742|Plasminogen activator inhibitor 2 Ag:MCnc:Pt:PPP:Qn:Imm
C0482742|Plasminogen activator inhibitor 2 Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C2708576|Coagulation ecarin induced:Time:Pt:Bld:Qn:Coag
C2708576|Ecarin clotting time (ECT) [Time] in Blood by Coagulation assay
C2708576|Coagulation ecarin induced:Time:Point in time:Whole blood:Quantitative:Coagulation Assay
C2708576|ECT Bld
C2733735|PA Rist 250 ug/mL Bld
C2733735|Platelet aggregation.ristocetin induced^250 ug/mL:RelACnc:Pt:Bld:Qn
C2733735|Platelet aggregation.ristocetin induced^250 ug/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733735|Platelet aggregation ristocetin induced in Blood --250 ug/mL
C3259770|Clotting time of Blood by Heparin protamine titration
C3259770|Clotting time:Time:Pt:Bld:Qn:Heparin protamine titration
C3259770|Clotting time:Time:Point in time:Whole blood:Quantitative:Heparin protamine titration
C3259770|Clotting time Bld HPT
C0482753|Plasminogen Ag:ACnc:Pt:PPP:Qn:Imm
C0482753|PLG Ag PPP Imm-aCnc
C0482753|Plasminogen Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482753|Plasminogen Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0798350|Fibrin D-dimer [Presence] in Platelet poor plasma
C0798350|D Dimer PPP Ql
C0798350|Fibrin D-dimer:ACnc:Pt:PPP:Ord
C0798350|Fibrin D-dimer:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C0550593|Protein C/Coagulation factor IX:Mass Ratio:Point in time:Platelet poor plasma:Quantitative
C0550593|Protein C/Coagulation factor IX:MRto:Pt:PPP:Qn
C0550593|Prot C/Fact IX PPP
C0550593|Protein C/Coagulation factor IX [Mass Ratio] in Platelet poor plasma
C0551341|PI IgM Ser-aCnc
C0551341|Phosphatidylinositol Ab.IgM:ACnc:Pt:Ser:Qn
C0551341|Phosphatidylinositol IgM Ab [Units/volume] in Serum
C0551341|Phosphatidylinositol Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0800567|Phosphatidylethanolamine Ab.IgA:ACnc:Pt:Ser:Ord
C0800567|PE IgA Ser Ql
C0800567|Phosphatidylethanolamine IgA Ab [Presence] in Serum
C0800567|Phosphatidylethanolamine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Ordinal
C0800575|Phosphatidylinositol Ab.IgM:ACnc:Pt:Ser:Ord
C0800575|Phosphatidylinositol IgM Ab [Presence] in Serum
C0800575|PI IgM Ser Ql
C0800575|Phosphatidylinositol Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482662|Coagulation factor XIII Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482662|Coagulation factor XIII Ag actual/normal in Platelet poor plasma by Immunologic method
C0482662|Fact XIII Ag Act/Nor PPP Imm
C0482662|Coagulation factor XIII Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1316347|Coagulation tissue factor induced.factor substitution^1H post incubation after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316347|Coagulation tissue factor induced.factor substitution^1 hour post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316347|Prothrombin time (PT) factor substitution in control Platelet poor plasma by Coagulation assay --1H post incubation with normal plasma
C1316347|PT 1h NP Cont PPP
C0482709|Fibrinogen fragments Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482709|Fibrinogen Frg Ag PPP Imm-aCnc
C0482709|Fibrinogen fragments Ag:ACnc:Pt:PPP:Qn:Imm
C0482709|Fibrinogen fragments Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1114192|Coagulation surface induced.factor substitution^1H post incubation:Time:Pt:PPP:Qn
C1114192|Coagulation surface induced.factor substitution^1 hour post incubation:Time:Point in time:Platelet poor plasma:Quantitative
C1114192|aPTT 1h p Inc PPP
C1114192|aPTT.factor substitution in Platelet poor plasma --1 hour post incubation
C0482614|Fact IX Ag Act/Nor PPP Imm
C0482614|Coagulation factor IX Ag actual/normal in Platelet poor plasma by Immunologic method
C0482614|Coagulation factor IX Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482614|Coagulation factor IX Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482649|Coagulation factor XI activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482649|Coagulation factor XI activity actual/normal in Platelet poor plasma by Coagulation assay
C0482649|Fact XI Act/Nor PPP
C0482649|Coagulation factor XI activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482651|Coagulation factor XI Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482651|Coagulation factor XI Ag:ACnc:Pt:PPP:Qn:Imm
C0482651|Fact XI Ag PPP Imm-aCnc
C0482651|Coagulation factor XI Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1544102|Coagulation tissue factor induced^1D post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544102|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --1 day post XXX challenge
C1544102|Coagulation tissue factor induced^1 day post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544102|PT 1D p chal PPP
C1544429|Clot Lysis [Presence] in Platelet poor plasma by Coagulation assay
C1544429|Coagulum lysis:ACnc:Pt:PPP:Ord:Coag
C1544429|Clot Lysis PPP Ql
C1544429|Coagulum lysis:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C1978749|Platelet factor 4 Ag:ACnc:Pt:PPP:Ord:Imm
C1978749|PF4 Ag PPP Ql Imm
C1978749|Platelet factor 4 Ag [Presence] in Platelet poor plasma by Immunologic method
C1978749|Platelet factor 4 Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Imm
C0482681|Deprecated TT PPP Qn
C0482681|Coagulation thrombin induced:Time:Pt:PPP:Qn:Tilt tube
C0482681|Deprecated Thrombin time in Platelet poor plasma by Coagulation assay
C0482681|Coagulation thrombin induced:Time:Point in time:Platelet poor plasma:Quantitative:Tilt tube
C0482735|Plasminogen:ACnc:Pt:PPP:Qn:Chromo
C0482735|Plasminogen [Units/volume] in Platelet poor plasma by Chromogenic method
C0482735|PLG PPP Chro-aCnc
C0482735|Plasminogen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C2708571|PA Rist 1000 ug/mL PRP
C2708571|Platelet aggregation ristocetin induced in Platelet rich plasma --1000 ug/mL
C2708571|Platelet aggregation.ristocetin induced^1000 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C2708571|Platelet aggregation.ristocetin induced^1000 ug/mL:RelACnc:Pt:PRP:Qn
C2733734|PA Coll 5 ug/mL Bld
C2733734|Platelet aggregation.collagen induced^5 ug/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733734|Platelet aggregation.collagen induced^5 ug/mL:RelACnc:Pt:Bld:Qn
C2733734|Platelet aggregation collagen induced in Blood --5 ug/mL
C3259335|Clotting time^after addition of heparinase:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C3259335|Clotting time^after addition of heparinase:Time:Pt:Bld:Qn:Thromboelastography
C3259335|Clotting time of Blood by Thromboelastography --after addition of heparinase
C3259335|Clotting time Heparinase Bld TEG
C3533726|Protein S Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C3533726|Prot S Ag PPP Imm-aCnc
C3533726|Protein S Ag [Units/volume] in Platelet poor plasma by Immunologic method
C3533726|Protein S Ag:ACnc:Pt:PPP:Qn:Imm
C0799300|Beta 2 glycoprotein 1 IgG Ab [Units/volume] in Serum
C0799300|B2 Glycoprot1 IgG Ser-aCnc
C0799300|Beta 2 glycoprotein 1 Ab.IgG:ACnc:Pt:Ser:Qn
C0799300|Beta 2 glycoprotein 1 Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0551327|Phosphatidate IgA Ab [Units/volume] in Serum
C0551327|Phosphatidate Ab.IgA:ACnc:Pt:Ser:Qn
C0551327|Phosphatidate IgA Ser-aCnc
C0551327|Phosphatidate Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C0551337|Phosphatidylglycerol Ab.IgG:ACnc:Pt:Ser:Qn
C0551337|Phosphatidylglycerol IgG Ab [Units/volume] in Serum
C0551337|PG IgG Ser-aCnc
C0551337|Phosphatidylglycerol Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0796812|Deprecated TT Qn
C0796812|Coagulation thrombin induced:Time:Pt::Qn:Coag
C0796812|Deprecated Thrombin time in Platelet poor plasma from control by Coagulation assay
C0796812|Coagulation thrombin induced:Time:Point in time::Quantitative:Coagulation Assay
C0365449|Heparin.low molecular weight:MRat:24H:Urine:Qn
C0365449|LMW Heparin [Mass/time] in 24 hour Urine
C0365449|Heparin.low molecular weight:Mass Rate:24 hours:Urine:Quantitative
C0365449|LMWH 24h Ur-mRate
C0482722|Heparin unfractionated [Units/volume] in Platelet poor plasma by Chromogenic method
C0482722|UFH PPP Chro-aCnc
C0482722|Heparin.unfractionated:ACnc:Pt:PPP:Qn:Chromo
C0482722|Heparin.unfractionated:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482716|Heparin Ab PPP Qn Pl Agg
C0482716|Heparin Ab:Threshold:Pt:PPP:Qn:Platelet aggr
C0482716|Heparin Ab [Threshold] in Platelet poor plasma by Platelet aggregation
C0482716|Heparin Antibody:Threshold:Point in time:Platelet poor plasma:Quantitative:Platelet aggr
C1316023|PA Rist 300 ug/mL PRP
C1316023|Platelet aggregation.ristocetin induced^300 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1316023|Platelet aggregation ristocetin induced in Platelet rich plasma --300 ug/mL
C1316023|Platelet aggregation.ristocetin induced^300 ug/mL:RelACnc:Pt:PRP:Qn
C2361202|MCF.fibrinolysis supp Bld TEG
C2361202|Maximum clot firmness.extrinsic coagulation system activated.fibrinolysis suppressed [Length] in Blood by Thromboelastography
C2361202|Maximum clot firmness.extrinsic coagulation system activated.fibrinolysis suppressed:Length:Point in time:Whole blood:Quantitative:Thromboelastography
C2361202|Maximum clot firmness.extrinsic coagulation system activated.fibrinolysis suppressed:Len:Pt:Bld:Qn:Thromboelastography
C2361210|MCF.extrinsic Bld TEG
C2361210|Maximum clot firmness.extrinsic coagulation system activated [Length] in Blood by Thromboelastography
C2361210|Maximum clot firmness.extrinsic coagulation system activated:Len:Pt:Bld:Qn:Thromboelastography
C2361210|Maximum clot firmness.extrinsic coagulation system activated:Length:Point in time:Whole blood:Quantitative:Thromboelastography
C2361216|Maximum lysis.extrinsic coagulation system activated:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C2361216|ML.extrinsic LenFr Bld TEG
C2361216|Maximum lysis.extrinsic coagulation system activated:LenFr:Pt:Bld:Qn:Thromboelastography
C2361216|Maximum lysis.extrinsic coagulation system activated [Length fraction] in Blood by Thromboelastography
C1976964|Platelet function:Imp:Pt:Bld:Nar
C1976964|Closure Tme Bld-Imp
C1976964|Platelet function:Impression/interpretation of study:Point in time:Whole blood:Narrative
C1976964|Platelet function (closure time) [Interpretation] in Blood Narrative
C1953451|Fibrin D-dimer DDU:MCnc:Pt:PPP:Qn
C1953451|D dimer DDU PPP-mCnc
C1953451|Fibrin D-dimer DDU [Mass/volume] in Platelet poor plasma
C1953451|Fibrin D-dimer DDU:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C0482736|Plasminogen activator tissue type Ag [Mass/volume] in Platelet poor plasma by Immunologic method --10 minutes post venistasis
C0482736|Plasminogen activator tissue type Ag^10M post venistasis:MCnc:Pt:PPP:Qn:Imm
C0482736|tPA Ag 10M PPP Imm-mCnc
C0482736|Plasminogen activator tissue type Antigen^10 minutes post venistasis:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0365493|PA AA PRP
C0365493|Platelet aggregation arachidonate induced in Platelet rich plasma
C0365493|Platelet aggregation.arachidonate induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0365493|Platelet aggregation.arachidonate induced:RelACnc:Pt:PRP:Qn
C0482762|Protein C+Acarboxy Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482762|Prot C+ACA Ag PPP Imm-aCnc
C0482762|Protein C+Acarboxy Ag:ACnc:Pt:PPP:Qn:Imm
C0482762|Protein C+Acarboxy Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0485836|Cardiolipin Ab:ACnc:Pt:Ser:Qn
C0485836|Cardiolipin Ab [Units/volume] in Serum
C0485836|Cardiolipin Ab Ser-aCnc
C0485836|Cardiolipin Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C3481507|Coagulation reptilase induced actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3481507|Coagulation reptilase induced actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3481507|Reptilase time/normal
C3481507|Reptilase time actual/Normal
C3481709|Rosner index in Platelet poor plasma by Coagulation assay
C3481709|Rosner index:RelTime:Pt:PPP:Qn:Coag
C3481709|Rosner index PPP
C3481709|Rosner index:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0040053|Thromboses
C0040053|Thrombosis
C0040053|Blood vessel thrombosis
C0040053|Thrombotic disorder (disorder)
C0040053|Thrombotic disorder (navigational concept)
C0040053|Thrombosis (disorder)
C0040053|Thrombosis [Disease/Finding]
C0040053|Thrombosis NOS
C0040053|Thrombosis (qualifier value)
C0040053|Thrombotic disorder
C0040053|Thrombosis, NOS
C0485826|Phosphatidylserine IgG Ab [Presence] in Serum by Immunoassay
C0485826|PS IgG Ser Ql EIA
C0485826|Phosphatidylserine Ab.IgG:ACnc:Pt:Ser:Ord:EIA
C0485826|Phosphatidylserine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal:Enzyme Immunoassay
C0484863|Coagulation factor VIII Ag:ACnc:Pt:Tiss:Ord:Immune stain
C0484863|Coagulation factor VIII Ag [Presence] in Tissue by Immune stain
C0484863|Fact VIII Ag Tiss Ql ImStn
C0484863|Coagulation factor VIII Antigen:Arbitrary Concentration:Point in time:Tissue, unspecified:Ordinal:Immune stain
C0798530|Coagulation surface induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C0798530|Coagulation surface induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0798530|aPTT imm 1:4 NP PPP
C0798530|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after 1:4 addition of normal plasma
C0800572|Phosphatidylglycerol IgM Ab [Presence] in Serum
C0800572|Phosphatidylglycerol Ab.IgM:ACnc:Pt:Ser:Ord
C0800572|PG IgM Ser Ql
C0800572|Phosphatidylglycerol Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal
C0882498|Cardiolipin IgG Ser Ql EIA
C0882498|Cardiolipin IgG Ab [Presence] in Serum by Immunoassay
C0882498|Cardiolipin Ab.IgG:ACnc:Pt:Ser:Ord:EIA
C0882498|Cardiolipin Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1316076|Phosphatidylethanolamine Ab:ACnc:Pt:Ser:Qn
C1316076|PE Ab Ser-aCnc
C1316076|Phosphatidylethanolamine Ab [Units/volume] in Serum
C1316076|Phosphatidylethanolamine Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C1315775|Phosphatidate Ab Ser Ql
C1315775|Phosphatidate Ab:ACnc:Pt:Ser:Ord
C1315775|Phosphatidate Ab [Presence] in Serum
C1315775|Phosphatidate Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C1315777|Phosphatidylethanolamine Ab:ACnc:Pt:Ser:Ord
C1315777|Phosphatidylethanolamine Ab [Presence] in Serum
C1315777|PE Ab Ser Ql
C1315777|Phosphatidylethanolamine Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482698|Fibrin D-dimer:ACnc:Pt:PPP:Qn:EIA
C0482698|Fibrin D-dimer [Units/volume] in Platelet poor plasma by Immunoassay
C0482698|D Dimer PPP EIA-aCnc
C0482698|Fibrin D-dimer:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C0482621|Fact VIIa PPP-aCnc
C0482621|Coagulation factor VII activated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482621|Coagulation factor VII activated activity:ACnc:Pt:PPP:Qn:Coag
C0482621|Coagulation factor VII activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482637|Coagulation factor VIII Ag [Units/volume] in Platelet poor plasma by Immunoelectrophoresis
C0482637|Coagulation factor VIII Ag:ACnc:Pt:PPP:Qn:Immunoelectrophoresis
C0482637|Fact VIII Ag PPP IEP-aCnc
C0482637|Coagulation factor VIII Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Immunoelectrophoresis
C0482653|Coagulation factor XII inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482653|Coagulation factor XII inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482653|Fact XII Inhib PPP-aCnc
C0482653|Coagulation factor XII inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1831367|Phosphatidate IgM Ab [Units/volume] in Serum by Immunoassay
C1831367|Phosphatidate Ab.IgM:ACnc:Pt:Ser:Qn:EIA
C1831367|Phosphatidate IgM Ser EIA-aCnc
C1831367|Phosphatidate Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C2360411|PA ADP 10 umol/L PRP Ql
C2360411|Platelet aggregation.adenosine diphosphate induced^10 umol/L:Pr:Pt:PRP:Ord
C2360411|Platelet aggregation ADP induced [Presence] in Platelet rich plasma --10 umol/L
C2360411|Platelet aggregation.adenosine diphosphate induced^10 umol/L:Presence:Point in time:Platelet rich plasma:Ordinal
C1977080|Protein C/Coagulation factor X:MRto:Pt:PPP:Qn
C1977080|Protein C/Coagulation factor X:Mass Ratio:Point in time:Platelet poor plasma:Quantitative
C1977080|Protein C/Coagulation factor X [Mass Ratio] in Platelet poor plasma
C1977080|Prot C/Fact X PPP
C1953385|Coagulation surface induced.lupus sensitive actual/Normal:RelTime:Pt:PPP:Qn
C1953385|Coagulation surface induced.lupus sensitive actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative
C1953385|aPTT.lupus sensitive actual/normal (normalized LA screen)
C1953385|Screen aPTT/normal
C0482682|Coagulation tissue factor induced actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482682|Coagulation tissue factor induced actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482682|Prothrombin time (PT) actual/Normal
C0482682|Prothrombin time/nomal
C2708405|Coagulation surface induced.factor substitution^5M post incubation after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C2708405|Coagulation surface induced.factor substitution^5 minutes post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C2708405|aPTT 5M p NP Cont PPP
C2708405|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --5 minutes post incubation after addition of normal plasma
C0365500|Platelet aggregation thrombin induced [Units threshold] in Platelet rich plasma
C0365500|PA Thrombin PRP
C0365500|Platelet aggregation.thrombin induced:ThrACnc:Pt:PRP:Qn
C0365500|Platelet aggregation.thrombin induced:Threshold Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0482756|Platelet factor 4 Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482756|PF4 Ag PPP Imm-mCnc
C0482756|Platelet factor 4 Ag:MCnc:Pt:PPP:Qn:Imm
C0482756|Platelet factor 4 Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0798330|Extrins clotting path PPP-Imp
C0798330|Coagulation factor.extrinsic pathway:Imp:Pt:PPP:Nar
C0798330|Coagulation factor.extrinsic pathway:Impression/interpretation of study:Point in time:Platelet poor plasma:Narrative
C0798330|Coagulation factor extrinsic pathway [Interpretation] in Platelet poor plasma Narrative
C0798362|Lupus anticoagulant neutralization dilute phospholipid [Presence] in Platelet poor plasma
C0798362|Lupus anticoagulant neutralization.dilute phospholipid:ACnc:Pt:PPP:Ord
C0798362|Lupus anticoagulant neutralization.dilute phospholipid:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C0798362|LA Nt dPL PPP Ql
C0550595|Protein S/Coagulation factor IX [Mass Ratio] in Platelet poor plasma by Coagulation assay
C0550595|Protein S/Coagulation factor IX:Mass Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0550595|Protein S/Coagulation factor IX:MRto:Pt:PPP:Qn:Coag
C0550595|Prot S/Fact IX PPP
C0550588|Coagulation surface induced^2nd specimen:Time:Pt:PPP:Qn:Coag
C0550588|Coagulation surface induced^2nd specimen:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0550588|aPTT sp2 PPP
C0550588|aPTT in Platelet poor plasma by Coagulation assay --2nd specimen
C0943512|Beta 2 glycoprotein 1 Ab:ACnc:Pt:Ser:Ord:EIA
C0943512|Beta 2 glycoprotein 1 Ab [Presence] in Serum by Immunoassay
C0943512|B2 Glycoprot1 Ab Ser Ql EIA
C0943512|Beta 2 glycoprotein 1 Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal:Enzyme Immunoassay
C0881643|Platelet aggregation ADP induced [Presence] in Platelet rich plasma
C0881643|Platelet aggregation.adenosine diphosphate induced:ACnc:Pt:PRP:Ord
C0881643|PA ADP PRP Ql
C0881643|Platelet aggregation.adenosine diphosphate induced:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C0881651|Cardiolipin Ab.IgM:ACnc:Pt:Ser:Ord:EIA
C0881651|Cardiolipin IgM Ser Ql EIA
C0881651|Cardiolipin IgM Ab [Presence] in Serum by Immunoassay
C0881651|Cardiolipin Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1316077|PI Ab Ser-aCnc
C1316077|Phosphatidylinositol Ab [Units/volume] in Serum
C1316077|Phosphatidylinositol Ab:ACnc:Pt:Ser:Qn
C1316077|Phosphatidylinositol Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C1316906|Acarboxyprothrombin SerPl-mCnc
C1316906|Acarboxyprothrombin:MCnc:Pt:Ser/Plas:Qn
C1316906|Acarboxyprothrombin [Mass/volume] in Serum or Plasma
C1316906|Acarboxyprothrombin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0482664|Coagulation factor XIII coagulum dissolution at 24H:ACnc:Pt:PPP:Ord:Coag
C0482664|Coagulation factor XIII coagulum dissolution at 24H:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C0482664|Fact XIII Clot Dis 24h PPP Ql
C0482664|Coagulation factor XIII coagulum dissolution at 24 hours [Presence] in Platelet poor plasma by Coagulation assay
C0482703|FSP PPP LA-aCnc
C0482703|Fibrin+Fibrinogen fragments:ACnc:Pt:PPP:Qn:LA
C0482703|Fibrin+Fibrinogen fragments [Units/volume] in Platelet poor plasma by Latex agglutination
C0482703|Fibrin+Fibrinogen fragments:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Latex Agglutination
C1315998|PA ADP lo dose PRP Cont
C1315998|Platelet aggregation.adenosine diphosphate induced^low dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma^Control:Quantitative
C1315998|Platelet aggregation.adenosine diphosphate induced^low dose:RelACnc:Pt:PRP^control:Qn
C1315998|Platelet aggregation ADP induced in control Platelet rich plasma --Low dose
C0482618|Coagulation factor V Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482618|Coagulation factor V Ag:ACnc:Pt:PPP:Qn:Imm
C0482618|Fact V Ag PPP Imm-aCnc
C0482618|Coagulation factor V Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482633|Coagulation factor VIII activity actual/normal in Platelet poor plasma by Coagulation assay
C0482633|Coagulation factor VIII activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482633|Fact VIII Act/Nor PPP
C0482633|Coagulation factor VIII activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1114317|Cardiolipin IgA Ser Ql
C1114317|Cardiolipin Ab.IgA:ACnc:Pt:Ser:Ord
C1114317|Cardiolipin IgA Ab [Presence] in Serum
C1114317|Cardiolipin Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Ordinal
C0366903|PK PPP-mCnc
C0366903|Prekallikrein (Fletcher Factor) [Mass/volume] in Platelet poor plasma
C0366903|Prekallikrein:MCnc:Pt:PPP:Qn
C0366903|Prekallikrein:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C1624144|Phosphatidylcholine IgM Ab B2GP1 independent [Multiple of the median] in Serum
C1624144|PC IgM B2GP1 indep MoM Ser
C1624144|Phosphatidylcholine Ab.IgM.B2GP1 independent:MoM:Pt:Ser:Qn
C1624144|Phosphatidylcholine Antibody.immunoglobulin M.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1623608|PE IgM B2GP1 indep MoM Ser
C1623608|Phosphatidylethanolamine Ab.IgM.B2GP1 independent:MoM:Pt:Ser:Qn
C1623608|Phosphatidylethanolamine IgM Ab B2GP1 independent [Multiple of the median] in Serum
C1623608|Phosphatidylethanolamine Antibody.immunoglobulin M.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1978978|Platelet aggregation.adenosine diphosphate induced^2 umol/L:Pr:Pt:PRP:Ord
C1978978|Platelet aggregation ADP induced [Presence] in Platelet rich plasma --2 umol/L
C1978978|PA ADP 2 umol/L PRP Ql
C1978978|Platelet aggregation.adenosine diphosphate induced^2 umol/L:Presence:Point in time:Platelet rich plasma:Ordinal
C0482769|Prot S PPP-aCnc
C0482769|Protein S [Units/volume] in Platelet poor plasma by Coagulation assay
C0482769|Protein S:ACnc:Pt:PPP:Qn:Coag
C0482769|Protein S:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3699646|Fondaparinux [Mass/volume] in Platelet poor plasma by Chromogenic method
C3699646|Fondaparinux:MCnc:Pt:PPP:Qn:Chromo
C3699646|Fondaparinux PPP Chro-mCnc
C3699646|Fondaparinux:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0799777|Coagulation surface induced:Time:Pt:Bld^control:Qn:Coag.saline 1:1
C0799777|Coagulation surface induced:Time:Point in time:Whole blood^Control:Quantitative:Coagulation Assay.saline 1:1
C0799777|aPTT Cont Bld 1:1 saline
C0799777|aPTT in control Blood by Coagulation 1:1 saline
C0551340|Phosphatidylinositol Ab.IgG:ACnc:Pt:Ser:Qn
C0551340|Phosphatidylinositol IgG Ab [Units/volume] in Serum
C0551340|PI IgG Ser-aCnc
C0551340|Phosphatidylinositol Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0804258|Plasminogen activator urokinase type:ACnc:Pt:Tiss:Ord
C0804258|Plasminogen activator urokinase type [Presence] in Tissue
C0804258|uPA Tiss Ql
C0804258|Plasminogen activator urokinase type:Arbitrary Concentration:Point in time:Tissue, unspecified:Ordinal
C0941825|Prothrombin Fragment 1.2 [Moles/volume] in Serum or Plasma
C0941825|Prothrombin fragment 1+2:SCnc:Pt:Ser/Plas:Qn
C0941825|Pro Frg1+2 SerPl-sCnc
C0941825|Prothrombin fragment 1+2:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1316061|Platelet factor 4 [Presence] in Platelet poor plasma
C1316061|Platelet factor 4:ACnc:Pt:PPP:Ord
C1316061|PF4 PPP Ql
C1316061|Platelet factor 4:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C1316350|Coagulation tissue factor induced.factor substitution^2H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1316350|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --2H post incubation with normal plasma
C1316350|Coagulation tissue factor induced.factor substitution^2 hours post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1316350|PT 2h NP PPP
C1316000|PA AA PRP Cont
C1316000|Platelet aggregation arachidonate induced in control Platelet rich plasma
C1316000|Platelet aggregation.arachidonate induced:RelACnc:Pt:PRP^control:Qn
C1316000|Platelet aggregation.arachidonate induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma^Control:Quantitative
C1316019|PA Rist 1500 ug/mL PRP
C1316019|Platelet aggregation.ristocetin induced^1500 ug/mL:RelACnc:Pt:PRP:Qn
C1316019|Platelet aggregation ristocetin induced in Platelet rich plasma --1500 ug/mL
C1316019|Platelet aggregation.ristocetin induced^1500 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1114191|Coagulation surface induced.factor substitution^1H post incubation:Time:Pt:PPP^control:Qn:Coag
C1114191|Coagulation surface induced.factor substitution^1 hour post incubation:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1114191|aPTT 1h p Inc Cont PPP
C1114191|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --1 hour post incubation
C1146843|Fibrinogen Ag/Fibrinogen:MRto:Pt:PPP:Qn
C1146843|Fibrinogen Ag/Fibrinogen [Mass Ratio] in Platelet poor plasma
C1146843|Fibrinogen Ag/Func PPP
C1146843|Fibrinogen Antigen/Fibrinogen:Mass Ratio:Point in time:Platelet poor plasma:Quantitative
C0365327|Clotting time:Time:Pt:Bld:Qn:Lee White
C0365327|Clotting time of Blood by Lee White method
C0365327|Clotting time:Time:Point in time:Whole blood:Quantitative:Lee White
C0365327|Clotting time Bld Lee White
C0482613|Coagulation factor IX Ag:ACnc:Pt:PPP:Qn:Imm
C0482613|Coagulation factor IX Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482613|Fact IX Ag PPP Imm-aCnc
C0482613|Coagulation factor IX Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1147715|Phosphatidylserine IgA Ab [Units/volume] in Serum by Immunoassay
C1147715|PS IgA Ser EIA-aCnc
C1147715|Phosphatidylserine Ab.IgA:ACnc:Pt:Ser:Qn:EIA
C1147715|Phosphatidylserine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1544678|Heparin Ab PPP Ql Pl Agg
C1544678|Heparin Ab [Presence] in Platelet poor plasma by Platelet aggregation
C1544678|Heparin Ab:ACnc:Pt:PPP:Ord:Platelet aggr
C1544678|Heparin Antibody:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Platelet aggr
C2361733|Coagulation factor XI activated [Units/volume] in Platelet poor plasma by Coagulation assay
C2361733|Fact XIa PPP-aCnc
C2361733|Coagulation factor XI activated activity:ACnc:Pt:PPP:Qn:Coag
C2361733|Coagulation factor XI activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1978231|Lupus anticoagulant neutralization dilute phospholipid actual/normal in Platelet poor plasma by Coagulation assay
C1978231|Lupus anticoagulant neutralization.dilute phospholipid actual/Normal:RelTime:Pt:PPP:Qn:Coag
C1978231|Lupus anticoagulant neutralization.dilute phospholipid actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1978231|LA Nt dPL Act/Nor PPP
C0482671|Coagulation surface induced.factor substitution^20M post incubation after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C0482671|Coagulation surface induced.factor substitution^20 minutes post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482671|aPTT 20M NP Cont PPP
C0482671|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --20M post incubation with normal plasma
C0482689|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C0482689|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C0482689|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482689|PT imm NP PPP
C0365471|Plasminogen activator tissue type Ag:MCnc:Pt:PPP:Qn:Imm
C0365471|Plasminogen activator tissue type Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0365471|tPA Ag PPP Imm-mCnc
C0365471|Plasminogen activator tissue type Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482738|Plasminogen activator inhibitor 1 [Units/volume] in Platelet poor plasma by Chromogenic method
C0482738|Plasminogen activator inhibitor 1:ACnc:Pt:PPP:Qn:Chromo
C0482738|PAI1 PPP Chro-aCnc
C0482738|Plasminogen activator inhibitor 1:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482740|PAI2 PPP Chro-aCnc
C0482740|Plasminogen activator inhibitor 2:ACnc:Pt:PPP:Qn:Chromo
C0482740|Plasminogen activator inhibitor 2 [Units/volume] in Platelet poor plasma by Chromogenic method
C0482740|Plasminogen activator inhibitor 2:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C2736262|Coagulation dilute Russell viper venom induced.excess phospholipid:Time:Pt:PPP:Qn
C2736262|Coagulation dilute Russell viper venom induced.excess phospholipid:Time:Point in time:Platelet poor plasma:Quantitative
C2736262|Confirm dRVVT
C2736262|dRVVT W excess phospholipid (LA confirm)
C2733975|PA Rist 1.0 mg/mL Bld
C2733975|Platelet aggregation.ristocetin induced^1.0 mg/mL:RelACnc:Pt:Bld:Qn
C2733975|Platelet aggregation.ristocetin induced^1.0 mg/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733975|Platelet aggregation ristocetin induced in Blood --1.0 mg/mL
C0178635|fibrinopeptide
C0178635|Fibrinopeptide (substance)
C0800574|PI IgG Ser Ql
C0800574|Phosphatidylinositol IgG Ab [Presence] in Serum
C0800574|Phosphatidylinositol Ab.IgG:ACnc:Pt:Ser:Ord
C0800574|Phosphatidylinositol Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C0800578|Phospholipid IgA Ser EIA-aCnc
C0800578|Phospholipid IgA Ab [Units/volume] in Serum by Immunoassay
C0800578|Phospholipid Ab.IgA:ACnc:Pt:Ser:Qn:EIA
C0800578|Phospholipid Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1316450|Heparin CF II Act/Nor PPP Chro
C1316450|Heparin cofactor II actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C1316450|Heparin cofactor II actual/normal in Platelet poor plasma by Chromogenic method
C1316450|Heparin cofactor II actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482725|Kininogen HMW actual/normal in Platelet poor plasma by Immunologic method
C0482725|HMWK Act/Nor PPP Imm
C0482725|Kininogen.high molecular weight actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482725|Kininogen.high molecular weight actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0365457|Kininogen.low molecular weight:MCnc:Pt:Ser:Qn:Imm
C0365457|LMWK Ser Imm-mCnc
C0365457|Kininogen LMW [Mass/volume] in Serum by Immunologic method
C0365457|Kininogen.low molecular weight:Mass Concentration:Point in time:Serum:Quantitative:Imm
C1315825|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --1H post incubation with normal plasma
C1315825|Coagulation tissue factor induced.factor substitution^1H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1315825|Coagulation tissue factor induced.factor substitution^1 hour post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1315825|PT 1h NP PPP
C1316343|Coagulation tissue factor induced.factor substitution^2H post incubation after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316343|Coagulation tissue factor induced.factor substitution^2 hours post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316343|Prothrombin time (PT) factor substitution in control Platelet poor plasma by Coagulation assay --2H post incubation with normal plasma
C1316343|PT 2h NP Cont PPP
C1315994|Coagulation thrombin induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1315994|Thrombin time.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C1315994|Coagulation thrombin induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1315994|TT imm NP PPP
C0482606|AT III PPP Chro-sCnc
C0482606|Antithrombin:SCnc:Pt:PPP:Qn:Chromo
C0482606|Antithrombin [Moles/volume] in Platelet poor plasma by Chromogenic method
C0482606|Antithrombin:Substance Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482642|Coagulation factor X activity:ACnc:Pt:PPP:Qn:Chromo
C0482642|Fact X PPP Chro-aCnc
C0482642|Coagulation factor X activity [Units/volume] in Platelet poor plasma by Chromogenic method
C0482642|Coagulation factor X activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482650|Coagulation factor XI activity:ACnc:Pt:PPP:Qn:Chromo
C0482650|Coagulation factor XI activity [Units/volume] in Platelet poor plasma by Chromogenic method
C0482650|Fact XI PPP Chro-aCnc
C0482650|Coagulation factor XI activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1544092|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --baseline
C1544092|Coagulation tissue factor induced^baseline:Time:Pt:PPP:Qn:Coag
C1544092|Coagulation tissue factor induced^baseline:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544092|PT BS PPP
C1544100|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --8 hours post XXX challenge
C1544100|Coagulation tissue factor induced^8H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544100|Coagulation tissue factor induced^8 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544100|PT 8h p chal PPP
C1543631|Coagulation factor X inhibitor [Presence] in Platelet poor plasma by Coagulation assay
C1543631|Coagulation factor X inhibitor:ACnc:Pt:PPP:Ord:Coag
C1543631|Fact X Inhib PPP Ql
C1543631|Coagulation factor X inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C1830306|Prothrombin time (PT) in Capillary blood by Coagulation assay
C1830306|Coagulation tissue factor induced:Time:Pt:BldC:Qn:Coag
C1830306|Coagulation tissue factor induced:Time:Point in time:Blood capillary:Quantitative:Coagulation Assay
C1830306|PT BldC
C1624709|Phosphatidylcholine Ab.IgG.B2GP1 dependent:MoM:Pt:Ser:Qn
C1624709|Phosphatidylcholine IgG Ab B2GP1 dependent [Multiple of the median] in Serum
C1624709|PC IgG B2GP1 dep MoM Ser
C1624709|Phosphatidylcholine Antibody.immunoglobulin G.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C1714709|Cardiolipin Ab.IgG:MCnc:Pt:Ser:Qn
C1714709|Cardiolipin IgG Ser-mCnc
C1714709|Cardiolipin IgG Ab [Mass/volume] in Serum
C1714709|Cardiolipin Antibody.immunoglobulin G:Mass Concentration:Point in time:Serum:Quantitative
C2361192|Clotting time.extrinsic coagulation system activated.fibrinolysis suppressed:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361192|Clotting time.extrinsic coagulation system activated.fibrinolysis suppressed of Blood by Thromboelastography
C2361192|Clotting time.extrinsic coagulation system activated.fibrinolysis suppressed:Time:Pt:Bld:Qn:Thromboelastography
C2361192|CT.fibinolysis supp Bld TEG
C1954716|Coagulum retraction:VFr:Pt:Bld:Qn
C1954716|Clot Retraction [Volume Fraction] in Blood
C1954716|Clot Retract VFr Bld
C1954716|Coagulum retraction:Volume Fraction:Point in time:Whole blood:Quantitative
C0482665|Coagulation reptilase induced:Time:Pt:PPP^control:Qn:Coag
C0482665|Coagulation reptilase induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482665|Reptilase time in control Platelet poor plasma by Coagulation assay
C0482665|Reptilase time Cont PPP
C2706768|Coagulation surface induced.factor substitution^immediately after addition of factor V depleted plasma:Time:Pt:PPP:Qn:Coag
C2706768|Coagulation surface induced.factor substitution^immediately after addition of factor V depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2706768|aPTT imm FV DP PPP
C2706768|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor V depleted plasma
C2733694|Platelet aggregation.ristocetin induced^1000 mg/L:ACnc:Pt:PRP:Ord
C2733694|PA Rist 1000 mg/L PRP Ql
C2733694|Platelet aggregation ristocetin induced [Presence] in Platelet rich plasma --1000 mg/L
C2733694|Platelet aggregation.ristocetin induced^1000 mg/L:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C2733958|PA Coll ATP secr 1 ug/mL Bld
C2733958|Platelet aggregation.collagen induced ATP secretion^1 ug/mL:RelACnc:Pt:Bld:Qn
C2733958|Platelet aggregation collagen induced ATP secretion in Blood --1 ug/mL
C2733958|Platelet aggregation.collagen induced ATP secretion^1 ug/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C0482751|Plasminogen activator tissue type^10M post venistasis:MCnc:Pt:PPP:Qn:Chromo
C0482751|tPA 10M PPP Chro-mCnc
C0482751|Plasminogen activator tissue type [Mass/volume] in Platelet poor plasma by Chromogenic method --10 minutes post venistasis
C0482751|Plasminogen activator tissue type^10 minutes post venistasis:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1979796|Platelet function header
C0798152|Coagulation surface induced:Time:Pt:PPP:Qn:Coag
C0798152|Coagulation surface induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0798152|aPTT PPP
C0798152|aPTT in Platelet poor plasma by Coagulation assay
C0797428|PC IgG Ser Ql
C0797428|Phosphatidylcholine Ab.IgG:ACnc:Pt:Ser:Ord
C0797428|Phosphatidylcholine IgG Ab [Presence] in Serum
C0797428|Phosphatidylcholine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C0798300|Deprecated Fibrin D-dimer:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:ENZYME IMMUNOASSAY
C0798300|Deprecated D Dimer PPP EIA-mCnc
C0798300|Fibrin D-dimer:MCnc:Pt:PPP:Qn:EIA
C0798300|Fibrin D-dimer:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C0798300|Deprecated Fibrin D-dimer EIA
C0551331|Phosphatidylcholine Ab.IgG:ACnc:Pt:Ser:Qn
C0551331|Phosphatidylcholine IgG Ab [Units/volume] in Serum
C0551331|PC IgG Ser-aCnc
C0551331|Phosphatidylcholine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0551330|Phosphatidylcholine IgA Ab [Units/volume] in Serum
C0551330|PC IgA Ser-aCnc
C0551330|Phosphatidylcholine Ab.IgA:ACnc:Pt:Ser:Qn
C0551330|Phosphatidylcholine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C0797198|PC IgA Ser EIA-aCnc
C0797198|Phosphatidylcholine Ab.IgA:ACnc:Pt:Ser:Qn:EIA
C0797198|Phosphatidylcholine IgA Ab [Units/volume] in Serum by Immunoassay
C0797198|Phosphatidylcholine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0800568|PE IgG Ser Ql
C0800568|Phosphatidylethanolamine Ab.IgG:ACnc:Pt:Ser:Ord
C0800568|Phosphatidylethanolamine IgG Ab [Presence] in Serum
C0800568|Phosphatidylethanolamine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482720|Heparin.low molecular weight:ACnc:Pt:PPP:Qn:Chromo
C0482720|LMWH PPP Chro-aCnc
C0482720|LMW Heparin [Units/volume] in Platelet poor plasma by Chromogenic method
C0482720|Heparin.low molecular weight:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1316652|Coagulation surface induced.factor substitution^30M post incubation after addition of normal plasma:Time:Pt:PPP:Qn
C1316652|Coagulation surface induced.factor substitution^30 minutes post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative
C1316652|aPTT 30M NP PPP
C1316652|aPTT.factor substitution in Platelet poor plasma --30M post incubation with normal plasma
C0482700|Fibrin fragments Ag:ACnc:Pt:PPP:Qn:Imm
C0482700|Fibrin Frg Ag PPP Imm-aCnc
C0482700|Fibrin fragments Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482700|Fibrin fragments Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1315991|PA Rist hi dose PRP
C1315991|Platelet aggregation.ristocetin induced^high dose:RelACnc:Pt:PRP:Qn
C1315991|Platelet aggregation.ristocetin induced^high dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1315991|Platelet aggregation ristocetin induced in Platelet rich plasma --High dose
C1316055|Phosphatidylethanolamine Ab [Units/volume] in Serum by Immunoassay
C1316055|Phosphatidylethanolamine Ab:ACnc:Pt:Ser:Qn:EIA
C1316055|PE Ab Ser EIA-aCnc
C1316055|Phosphatidylethanolamine Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1146941|Beta 2 glycoprotein 1 Ab:ACnc:Pt:Ser:Ord
C1146941|Beta 2 glycoprotein 1 Ab [Presence] in Serum
C1146941|B2 Glycoprot1 Ab Ser Ql
C1146941|Beta 2 glycoprotein 1 Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482623|Fact VII PPP Chro-aCnc
C0482623|Coagulation factor VII activity [Units/volume] in Platelet poor plasma by Chromogenic method
C0482623|Coagulation factor VII activity:ACnc:Pt:PPP:Qn:Chromo
C0482623|Coagulation factor VII activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482644|Coagulation factor X Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482644|Coagulation factor X Ag actual/normal in Platelet poor plasma by Immunologic method
C0482644|Fact X Ag Act/Nor PPP Imm
C0482644|Coagulation factor X Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1113919|Fibrin+Fibrinogen fragments:MCnc:Pt:Ser:Qn
C1113919|Fibrin+Fibrinogen fragments [Mass/volume] in Serum
C1113919|FSP Ser-mCnc
C1113919|Fibrin+Fibrinogen fragments:Mass Concentration:Point in time:Serum:Quantitative
C1544105|Coagulation surface induced^30M post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544105|Coagulation surface induced^30 minutes post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544105|aPTT 30M p chal PPP
C1544105|aPTT in Platelet poor plasma by Coagulation assay --30 minutes post XXX challenge
C1544779|von Willebrand factor cleaving protease inhibitor:ACnc:Pt:PPP:Qn
C1544779|vWF Cp Inhib PPP-aCnc
C1544779|von Willebrand factor (vWf) cleaving protease inhibitor [Units/volume] in Platelet poor plasma
C1544779|von Willebrand factor cleaving protease inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0366906|Protein C Ag:MCnc:Pt:PPP:Qn
C0366906|Protein C Ag [Mass/volume] in Platelet poor plasma
C0366906|Prot C Ag PPP-mCnc
C0366906|Protein C Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C1624707|Cardiolipin IgM Ab B2GP1 independent [Multiple of the median] in Serum
C1624707|Cardiolipin Ab.IgM.B2GP1 independent:MoM:Pt:Ser:Qn
C1624707|Cardiolipin IgM B2GP1 indep MoM Ser
C1624707|Cardiolipin Antibody.immunoglobulin M.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1714708|Cardiolipin IgA Ab [Mass/volume] in Serum
C1714708|Cardiolipin Ab.IgA:MCnc:Pt:Ser:Qn
C1714708|Cardiolipin IgA Ser-mCnc
C1714708|Cardiolipin Antibody.immunoglobulin A:Mass Concentration:Point in time:Serum:Quantitative
C2360096|Coagulation tissue factor induced^post heparin adsorption:Time:Pt:PPP:Qn:Coag
C2360096|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --post heparin adsorption
C2360096|Coagulation tissue factor induced^post heparin adsorption:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2360096|PT p heparin adsorption PPP
C2361181|Clot formation [Time] in Blood by Thromboelastography
C2361181|Clot formation:Time:Pt:Bld:Qn:Thromboelastography
C2361181|Clot formation:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361181|CFT Bld TEG
C1978235|von Willebrand factor (vWf).collagen binding activity/von Willebrand factor Ag [Ratio] in Platelet poor plasma by Immunoassay
C1978235|vWF CBA/vWF Ag PPP EIA-Rto
C1978235|von Willebrand factor.collagen binding activity/von Willebrand factor Ag:Ratio:Pt:PPP:Qn:EIA
C1978235|von Willebrand factor.collagen binding activity/von Willebrand factor Antigen:Ratio:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C0365519|Prothrombin fragment 1+2:ACnc:Pt:Ser/Plas:Qn
C0365519|Pro Frg1+2 SerPl-aCnc
C0365519|Prothrombin Fragment 1.2 [Units/volume] in Serum or Plasma
C0365519|Prothrombin fragment 1+2:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C0482675|Coagulation surface induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C0482675|Coagulation surface induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482675|aPTT imm NP Cont PPP
C0482675|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C2733663|Cardiolipin IgG MoM Ser
C2733663|Cardiolipin IgG Ab [Multiple of the median] in Serum
C2733663|Cardiolipin Ab.IgG:MoM:Pt:Ser:Qn
C2733663|Cardiolipin Antibody.immunoglobulin G:Multiple of the median:Point in time:Serum:Quantitative
C2598680|PA Epineph 0.1 ug/mL PRP
C2598680|Platelet aggregation.epinephrine induced^0.1 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C2598680|Platelet aggregation epinephrine induced in Platelet rich plasma --0.1 ug/mL
C2598680|Platelet aggregation.epinephrine induced^0.1 ug/mL:RelACnc:Pt:PRP:Qn
C0367248|Streptokinase Ab Ser-aCnc
C0367248|Streptokinase Ab:ACnc:Pt:Ser:Qn
C0367248|Streptokinase Ab [Units/volume] in Serum
C0367248|Streptokinase Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C0482752|Plasminogen activator tissue type^20M post venistasis:ACnc:Pt:PPP:Qn:Chromo
C0482752|Plasminogen activator tissue type [Units/volume] in Platelet poor plasma by Chromogenic method --20 minutes post venistasis
C0482752|tPA 20M PPP Chro-aCnc
C0482752|Plasminogen activator tissue type^20 minutes post venistasis:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0365497|PA Norepineph PRP
C0365497|Platelet aggregation.norepinephrine induced:RelACnc:Pt:PRP:Qn
C0365497|Platelet aggregation norepinephrine induced in Platelet rich plasma
C0365497|Platelet aggregation.norepinephrine induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0365498|PA Rist PRP
C0365498|Platelet aggregation.ristocetin induced:RelACnc:Pt:PRP:Qn
C0365498|Platelet aggregation ristocetin induced in Platelet rich plasma
C0365498|Platelet aggregation.ristocetin induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0484871|Phospholipid IgM Ab [Units/volume] in Serum
C0484871|Phospholipid IgM Ser-aCnc
C0484871|Phospholipid Ab.IgM:ACnc:Pt:Ser:Qn
C0484871|Phospholipid Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0803297|Cardiolipin IgM Ab [Titer] in Serum
C0803297|Cardiolipin Ab.IgM:Titr:Pt:Ser:Qn
C0803297|Cardiolipin IgM Titr Ser
C0803297|Cardiolipin Antibody.immunoglobulin M:Dilution Factor (Titer):Point in time:Serum:Quantitative
C0943510|Coagulation factor XIII activity actual/normal in Platelet poor plasma by Chromogenic method
C0943510|Coagulation factor XIII activity actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C0943510|Fact XIII Act/Nor PPP Chro
C0943510|Coagulation factor XIII activity actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1369548|Coagulation tissue factor induced.factor substitution^immediately after addition of factor V depleted plasma:Time:Pt:PPP:Qn:Coag
C1369548|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor V depleted plasma
C1369548|Coagulation tissue factor induced.factor substitution^immediately after addition of factor V depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1369548|PT imm FV DP PPP
C1369553|Coagulation surface induced.factor substitution^immediately after addition of factor XI depleted plasma:Time:Pt:PPP:Qn:Coag
C1369553|Coagulation surface induced.factor substitution^immediately after addition of factor XI depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1369553|aPTT imm FXI DP PPP
C1369553|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor XI depleted plasma
C1316344|Coagulation tissue factor induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316344|Coagulation tissue factor induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316344|Prothrombin time (PT) factor substitution in control Platelet poor plasma by Coagulation assay --immediately after 1:4 addition of normal plasma
C1316344|PT imm 1:4 NP Cont PPP
C0482632|Coagulation factor VIII activated activity:ACnc:Pt:PPP:Qn:Coag
C0482632|Coagulation factor VIII activated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482632|Fact VIIIa PPP-aCnc
C0482632|Coagulation factor VIII activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1526518|Coagulation surface induced.factor substitution^2H post incubation:Time:Pt:PPP:Qn
C1526518|Coagulation surface induced.factor substitution^2 hours post incubation:Time:Point in time:Platelet poor plasma:Quantitative
C1526518|aPTT 2h p Inc PPP
C1526518|aPTT.factor substitution in Platelet poor plasma --2 hours post incubation
C0366905|Protein C [Mass/volume] in Plasma
C0366905|Protein C:MCnc:Pt:Plas:Qn
C0366905|Prot C Plas-mCnc
C0366905|Protein C:Mass Concentration:Point in time:Plasma:Quantitative
C1715217|Beta 2 glycoprotein 1 IgM Ab [Presence] in Serum
C1715217|B2 Glycoprot1 IgM Ser Ql
C1715217|Beta 2 glycoprotein 1 Ab.IgM:ACnc:Pt:Ser:Ord
C1715217|Beta 2 glycoprotein 1 Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal
C2361214|Maximum lysis.extrinsic coagulation system activated.fibrinolysis suppressed [Length fraction] in Blood by Thromboelastography
C2361214|Maximum lysis.extrinsic coagulation system activated.fibrinolysis suppressed:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C2361214|ML.fibrinolysis supp LenFr Bld TEG
C2361214|Maximum lysis.extrinsic coagulation system activated.fibrinolysis suppressed:LenFr:Pt:Bld:Qn:Thromboelastography
C0482694|Coagulation tissue factor induced:Time:Pt:PPP:Qn:Coag
C0482694|Coagulation tissue factor induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482694|Prothrombin time
C0482694|Prothrombin time (PT)
C2735003|Fibrinogen fragments [Mass/volume] in Urine
C2735003|Fibrinogen fragments:MCnc:Pt:Urine:Qn
C2735003|Fibrinogen Frg Ur-mCnc
C2735003|Fibrinogen fragments:Mass Concentration:Point in time:Urine:Quantitative
C2736263|Coagulation kaolin induced:Time:Pt:PPP^control:Qn
C2736263|Coagulation kaolin induced:Time:Point in time:Platelet poor plasma^Control:Quantitative
C2736263|Kaolin activated time in control Platelet poor plasma
C2736263|KCT Cont PPP
C2706769|Coagulation surface induced.factor substitution^immediately after addition of factor V depleted plasma+APC:Time:Pt:PPP:Qn:Coag
C2706769|Coagulation surface induced.factor substitution^immediately after addition of factor V depleted plasma+APC:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2706769|aPTT imm FV DP+APC PPP
C2706769|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor V depleted plasma+APC
C2733693|Platelet aggregation ristocetin induced [Presence] in Platelet rich plasma --1125 mg/L
C2733693|PA Rist 1125 mg/L PRP Ql
C2733693|Platelet aggregation.ristocetin induced^1125 mg/L:ACnc:Pt:PRP:Ord
C2733693|Platelet aggregation.ristocetin induced^1125 mg/L:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C0482757|PK PPP-aCnc
C0482757|Prekallikrein (Fletcher Factor) [Units/volume] in Platelet poor plasma
C0482757|Prekallikrein:ACnc:Pt:PPP:Qn
C0482757|Prekallikrein:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0485838|Cardiolipin Ab.IgG:ACnc:Pt:Ser/Plas:Qn
C0485838|Cardiolipin Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C0485838|Cardiolipin IgG SerPl-aCnc
C0485838|Cardiolipin IgG Ab [Units/volume] in Serum or Plasma
C1979801|Routine coag
C0797196|Phosphatidylcholine IgG Ab [Units/volume] in Serum by Immunoassay
C0797196|Phosphatidylcholine Ab.IgG:ACnc:Pt:Ser:Qn:EIA
C0797196|PC IgG Ser EIA-aCnc
C0797196|Phosphatidylcholine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0801359|Coagulation of Semen by Visual observation
C0801359|Coag Smn Ql Visual
C0801359|Coagulation:ACnc:Pt:Semen:Ord:Visual
C0801359|Coagulation:Arbitrary Concentration:Point in time:Seminal fluid:Ordinal:Visual
C0800570|Phosphatidylglycerol Ab.IgA:ACnc:Pt:Ser:Ord
C0800570|Phosphatidylglycerol IgA Ab [Presence] in Serum
C0800570|PG IgA Ser Ql
C0800570|Phosphatidylglycerol Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Ordinal
C0943506|AT III Act/Nor PPP Chro
C0943506|Antithrombin actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C0943506|Antithrombin actual/normal in Platelet poor plasma by Chromogenic method
C0943506|Antithrombin actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0944759|Fibrin D-dimer [Presence] in Platelet poor plasma by Latex agglutination
C0944759|D Dimer PPP Ql LA
C0944759|Fibrin D-dimer:ACnc:Pt:PPP:Ord:LA
C0944759|Fibrin D-dimer:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Latex Agglutination
C0945508|Protein C Ag/Coagulation factor VII Ag Ag [Mass Ratio] in Platelet poor plasma by Immunologic method
C0945508|Protein C Antigen/Coagulation factor VII Antigen:Mass Ratio:Point in time:Platelet poor plasma:Quantitative:Imm
C0945508|Protein C Ag/Coagulation factor VII Ag:MRto:Pt:PPP:Qn:Imm
C0945508|Prot C Ag/Fact VII Ag PPP Imm
C0881647|Platelet aggregation arachidonate induced [Presence] in Platelet rich plasma
C0881647|PA AA PRP Ql
C0881647|Platelet aggregation.arachidonate induced:ACnc:Pt:PRP:Ord
C0881647|Platelet aggregation.arachidonate induced:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C1315776|PC Ab Ser Ql
C1315776|Phosphatidylcholine Ab [Presence] in Serum
C1315776|Phosphatidylcholine Ab:ACnc:Pt:Ser:Ord
C1315776|Phosphatidylcholine Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482697|Clot Lysis [Time] in Platelet poor plasma by Coagulation assay
C0482697|Coagulum lysis:Time:Pt:PPP:Qn:Coag
C0482697|Coagulum lysis:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482697|Clot Lysis PPP
C1315988|PA ADP lo dose PRP
C1315988|Platelet aggregation.adenosine diphosphate induced^low dose:RelACnc:Pt:PRP:Qn
C1315988|Platelet aggregation ADP induced in Platelet rich plasma --Low dose
C1315988|Platelet aggregation.adenosine diphosphate induced^low dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0482607|Antithrombin Ag [Moles/volume] in Platelet poor plasma by Immunologic method
C0482607|Antithrombin Ag:SCnc:Pt:PPP:Qn:Imm
C0482607|AT III Ag PPP Imm-sCnc
C0482607|Antithrombin Antigen:Substance Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482622|Fact VII Act/Nor PPP
C0482622|Coagulation factor VII activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482622|Coagulation factor VII activity actual/normal in Platelet poor plasma by Coagulation assay
C0482622|Coagulation factor VII activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482629|Coagulation factor VIII Ab [Units/volume] in Platelet poor plasma by Immunologic method
C0482629|Fact VIII Ab PPP Imm-aCnc
C0482629|Coagulation factor VIII Ab:ACnc:Pt:PPP:Qn:Imm
C0482629|Coagulation factor VIII Antibody:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482634|Fact VIII PPP Chro-aCnc
C0482634|Coagulation factor VIII activity:ACnc:Pt:PPP:Qn:Chromo
C0482634|Coagulation factor VIII activity [Units/volume] in Platelet poor plasma by Chromogenic method
C0482634|Coagulation factor VIII activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1544107|Coagulation surface induced^1.5H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544107|Coagulation surface induced^1 1/2 hour post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544107|aPTT 1.5h p chal PPP
C1544107|aPTT in Platelet poor plasma by Coagulation assay --1.5 hours post XXX challenge
C1544552|Prothrom IgG SerPl-aCnc
C1544552|Prothrombin IgG Ab [Units/volume] in Serum or Plasma
C1544552|Prothrombin Ab.IgG:ACnc:Pt:Ser/Plas:Qn
C1544552|Prothrombin Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C1544657|Fibrin Monomer PPP Ql HA
C1544657|Fibrin monomer [Presence] in Platelet poor plasma by Hemagglutination
C1544657|Fibrin monomer:ACnc:Pt:PPP:Ord:HA
C1544657|Fibrin monomer:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Hemagglutination
C1831130|Phosphatidate Ab.IgA:ACnc:Pt:Ser:Qn:EIA
C1831130|Phosphatidate IgA Ser EIA-aCnc
C1831130|Phosphatidate IgA Ab [Units/volume] in Serum by Immunoassay
C1831130|Phosphatidate Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1704393|Deprecated Dilute Russell viper venom time (dRVVT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C1704393|Deprecated dRVV Tme imm NP PPP Qn
C1704393|Coagulation dilute Russell viper venom induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1704393|Coagulation dilute Russell viper venom induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2607830|Fibrinogen [Mass or Molecules/volume] in Platelet poor plasma by Coagulation assay
C2607830|Fibrinogen [Mass or Moles/volume] in Platelet poor plasma by Coagulation assay
C2607830|Fibrinogen PPP-msCnc
C2607830|Fibrinogen:MSCnc:Pt:PPP:Qn:Coag
C2607830|Fibrinogen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2360890|Coagulation surface induced.lupus sensitive.factor substitution^immediately after 4:1 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2360890|Coagulation surface induced.lupus sensitive.factor substitution^immediately after 4:1 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2360890|aPTT-LA imm 4:1 NP PPP
C2360890|aPTT.lupus sensitive.factor substitution in Platelet poor plasma by Coagulation assay --immediately after 4:1 addition of normal plasma
C1978748|Hirudin [Units/volume] in Platelet poor plasma by Chromogenic method
C1978748|Hirudin PPP Chro-aCnc
C1978748|Hirudin:ACnc:Pt:PPP:Qn:Chromo
C1978748|Hirudin:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1954718|Platelet aggregation.adenosine diphosphate induced:ACnc:Pt:PRP:Qn
C1954718|Platelet aggregation ADP induced [Units/volume] in Platelet rich plasma
C1954718|PA ADP PRP-aCnc
C1954718|Platelet aggregation.adenosine diphosphate induced:Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1953452|D dimer FEU PPP EIA-mCnc
C1953452|Fibrin D-dimer FEU:MCnc:Pt:PPP:Qn:EIA
C1953452|Fibrin D-dimer FEU [Mass/volume] in Platelet poor plasma by Immunoassay
C1953452|Fibrin D-dimer FEU:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C2733951|Platelet aggregation ADP induced ATP secretion in Blood --5 umol/L
C2733951|Platelet aggregation.adenosine diphosphate induced ATP secretion^5 umol/L:RelACnc:Pt:Bld:Qn
C2733951|PA ADP ATP secr 5 umol/L Bld
C2733951|Platelet aggregation.adenosine diphosphate induced ATP secretion^5 umol/L:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733736|Platelet aggregation.adenosine diphosphate induced ATP secretion^10 umol/L:RelACnc:Pt:Bld:Qn
C2733736|Platelet aggregation.adenosine diphosphate induced ATP secretion^10 umol/L:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733736|PA ADP ATP secr 10 umol/L Bld
C2733736|Platelet aggregation ADP induced ATP secretion in Blood --10 umol/L
C2598416|PA ADP 20 umol/mL PRP
C2598416|Platelet aggregation ADP induced in Platelet rich plasma --20 umol/mL
C2598416|Platelet aggregation.adenosine diphosphate induced^20 umol/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C2598416|Platelet aggregation.adenosine diphosphate induced^20 umol/mL:RelACnc:Pt:PRP:Qn
C3259769|Clot Lysis 30M p MA LenFr Bld TEG
C3259769|Clot Lysis [Length fraction] in Blood by Thromboelastography --30 minutes post maximum clot amplitude
C3259769|Coagulum lysis^30 minutes post maximum clot amplitude:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C3259769|Coagulum lysis^30M post maximum clot amplitude:LenFr:Pt:Bld:Qn:Thromboelastography
C0365499|PA Serotonin PRP
C0365499|Platelet aggregation.serotonin induced:RelACnc:Pt:PRP:Qn
C0365499|Platelet aggregation.serotonin induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0365499|Platelet aggregation serotonin induced in Platelet rich plasma
C0796781|Activated protein C resistance:TRto:Pt:PPP:Qn:Coag
C0796781|Activated protein C resistance [Time Ratio] in Platelet poor plasma by Coagulation assay
C0796781|aPCR PPP
C0796781|Activated protein C resistance:Time Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0364413|Fibrinopeptide A:MCnc:Pt:Periton fld:Qn
C0364413|Fibrinopeptide A [Mass/volume] in Peritoneal fluid
C0364413|FpA Prt-mCnc
C0364413|Fibrinopeptide A:Mass Concentration:Point in time:Peritoneal fluid /ascites:Quantitative
C0803470|Cardiolipin Ab.IgA:Titr:Pt:Ser:Qn
C0803470|Cardiolipin IgA Ab [Titer] in Serum
C0803470|Cardiolipin IgA Titr Ser
C0803470|Cardiolipin Antibody.immunoglobulin A:Dilution Factor (Titer):Point in time:Serum:Quantitative
C1369549|Coagulation surface induced.factor substitution^immediately after addition of factor IX depleted plasma:Time:Pt:PPP:Qn:Coag
C1369549|Coagulation surface induced.factor substitution^immediately after addition of factor IX depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1369549|aPTT imm FIX DP PPP
C1369549|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor IX depleted plasma
C0365463|Phospholipid Ab.IgG:ACnc:Pt:Ser:Qn:EIA
C0365463|Phospholipid IgG Ab [Units/volume] in Serum by Immunoassay
C0365463|Phospholipid IgG Ser EIA-aCnc
C0365463|Phospholipid Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0482714|Fibrinopeptide A Ag:MCnc:Pt:PPP:Qn:Imm
C0482714|FpA Ag PPP Imm-mCnc
C0482714|Fibrinopeptide A Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482714|Fibrinopeptide A Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0365392|Coagulation surface induced:Time:Pt:Bld:Qn:Coag
C0365392|Coagulation surface induced:Time:Point in time:Whole blood:Quantitative:Coagulation Assay
C0365392|aPTT Bld
C0365392|aPTT in Blood by Coagulation assay
C0482628|Coagulation factor VIII inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482628|Coagulation factor VIII inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482628|Fact VIII Inhib PPP-aCnc
C0482628|Coagulation factor VIII inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1526522|Coagulation factor VIII Ag actual/normal in Platelet poor plasma by Immunologic method
C1526522|Fact VIII Ag Act/Nor PPP Imm
C1526522|Coagulation factor VIII Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C1526522|Coagulation factor VIII Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1544699|Fact Inhib XXX PPP Ql
C1544699|Factor inhibitor XXX [Presence] in Platelet poor plasma by Coagulation assay
C1544699|Factor inhibitor XXX:ACnc:Pt:PPP:Ord:Coag
C1544699|Factor inhibitor XXX:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C0366902|Plasminogen Ag [Mass/volume] in Platelet poor plasma
C0366902|Plasminogen Ag:MCnc:Pt:PPP:Qn
C0366902|PLG Ag PPP-mCnc
C0366902|Plasminogen Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C1624145|Phosphatidylethanolamine Ab.IgG.B2GP1 independent:MoM:Pt:Ser:Qn
C1624145|PE IgG B2GP1 indep MoM Ser
C1624145|Phosphatidylethanolamine IgG Ab B2GP1 independent [Multiple of the median] in Serum
C1624145|Phosphatidylethanolamine Antibody.immunoglobulin G.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1632263|Cardiolipin Ab.IgG.B2GP1 dependent:MoM:Pt:Ser:Qn
C1632263|Cardiolipin IgG Ab B2GP1 dependent [Multiple of the median] in Serum
C1632263|Cardiolipin IgG B2GP1 dep MoM Ser
C1632263|Cardiolipin Antibody.immunoglobulin G.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C0482668|Russell viper venom time in Platelet poor plasma by Coagulation assay
C0482668|Coagulation Russell viper venom induced:Time:Pt:PPP:Qn:Coag
C0482668|Coagulation Russell viper venom induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482668|RVV time PPP
C0482731|Plasmin inhibitor [Units/volume] in Platelet poor plasma by Chromogenic method
C0482731|Plasm Inhib PPP Chro-aCnc
C0482731|Plasmin inhibitor:ACnc:Pt:PPP:Qn:Chromo
C0482731|Plasmin inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3258981|Heparin.unfractionated:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C3258981|Heparin.unfractionated:ACnc:Pt:PPP:Qn
C3258981|UFH PPP-aCnc
C3258981|Heparin unfractionated [Units/volume] in Platelet poor plasma
C3259331|Clot formation^after addition of heparinase:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C3259331|Clot formation^after addition of heparinase:Time:Pt:Bld:Qn:Thromboelastography
C3259331|Clot formation [Time] in Blood by Thromboelastography --after addition of heparinase
C3259331|CFT Heparinase Bld TEG
C0798531|Coagulation surface induced.inhibitor sensitive:Time:Pt:PPP:Qn:Coag
C0798531|Coagulation surface induced.inhibitor sensitive:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0798531|aPTT Inhib Sens PPP
C0798531|aPTT.inhibitor sensitive in Platelet poor plasma by Coagulation assay
C0550587|Coagulation surface induced:Time:Pt:PPP^control:Qn:Coag
C0550587|Coagulation surface induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0550587|aPTT Cont PPP
C0550587|aPTT in control Platelet poor plasma by Coagulation assay
C0364414|Fibrinopeptide B [Mass/volume] in Serum
C0364414|Fibrinopeptide B:MCnc:Pt:Ser:Qn
C0364414|FpB Ser-mCnc
C0364414|Fibrinopeptide B:Mass Concentration:Point in time:Serum:Quantitative
C0803240|Cardiolipin Ab.IgM:Imp:Pt:Ser:Nom
C0803240|Cardiolipin IgM Ser-Imp
C0803240|Cardiolipin Antibody.immunoglobulin M:Impression/interpretation of study:Point in time:Serum:Nominal
C0803240|Cardiolipin IgM Ab [Interpretation] in Serum
C0943518|Pro Frg1+2 Ag SerPl Imm-sCnc
C0943518|Prothrombin Fragment 1.2 Ag [Moles/volume] in Serum or Plasma by Immunologic method
C0943518|Prothrombin fragment 1+2 Ag:SCnc:Pt:Ser/Plas:Qn:Imm
C0943518|Prothrombin fragment 1+2 Antigen:Substance Concentration:Point in time:Serum/Plasma:Quantitative:Imm
C1317051|vWF Cp Inhib PPP Ql
C1317051|von Willebrand factor (vWf) cleaving protease inhibitor [Presence] in Platelet poor plasma
C1317051|von Willebrand factor cleaving protease inhibitor:ACnc:Pt:PPP:Ord
C1317051|von Willebrand factor cleaving protease inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C1369802|Deprecated FpA PPP EIA-mCnc
C1369802|Fibrinopeptide A:MCnc:Pt:PPP:Qn:EIA
C1369802|Fibrinopeptide A:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C1369802|Deprecated Fibrinopeptide A Ag [Mass/volume] in Platelet poor plasma by EIA
C1315778|Phosphatidylinositol Ab:ACnc:Pt:Ser:Ord
C1315778|PI Ab Ser Ql
C1315778|Phosphatidylinositol Ab [Presence] in Serum
C1315778|Phosphatidylinositol Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C2718109|Deprecated Fibrinogen Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C2718109|Deprecated Fibrinogen Ag PPP Imm-mCnc
C2718109|Fibrinogen Ag:MCnc:Pt:PPP:Qn:Imm
C2718109|Fibrinogen Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1316352|Coagulation surface induced.factor substitution^2H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316352|Coagulation surface induced.factor substitution^2 hours post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316352|aPTT 2h p 1:4 NP Cont PPP
C1316352|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --2H post incubation with 1:4 normal plasma
C0365325|Cardiolipin Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative:ENZYME IMMUNOASSAY
C0365325|Cardiolipin Ab.IgG:ACnc:Pt:Ser:Qn:EIA
C0365325|Cardiolipin IgG Ab [Units/volume] in Serum by Immunoassay
C0365325|Cardiolipin IgG Ser EIA-aCnc
C0482624|Coagulation factor VII activity actual/normal [Molar ratio] in Platelet poor plasma by Coagulation assay
C0482624|Fact VII Act/Nor PPP-sRto
C0482624|Coagulation factor VII activity actual/Normal:Substance Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482624|Coagulation factor VII activity actual/Normal:SRto:Pt:PPP:Qn:Coag
C1544094|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --1 hour post XXX challenge
C1544094|Coagulation tissue factor induced^1H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544094|Coagulation tissue factor induced^1 hour post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544094|PT 1h p chal PPP
C1544109|Coagulation surface induced^3H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544109|Coagulation surface induced^3 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544109|aPTT 3h p chal PPP
C1544109|aPTT in Platelet poor plasma by Coagulation assay --3 hours post XXX challenge
C1714867|Coagulation surface induced.factor substitution^1H post incubation after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1714867|Coagulation surface induced.factor substitution^1 hour post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1714867|aPTT 1h NP Cont PPP
C1714867|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --1H post incubation with normal plasma
C1624710|PC IgM B2GP1 dep MoM Ser
C1624710|Phosphatidylcholine IgM Ab B2GP1 dependent [Multiple of the median] in Serum
C1624710|Phosphatidylcholine Ab.IgM.B2GP1 dependent:MoM:Pt:Ser:Qn
C1624710|Phosphatidylcholine Antibody.immunoglobulin M.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C1623609|Phosphatidylserine Ab.IgG.B2GP1 dependent:MoM:Pt:Ser:Qn
C1623609|Phosphatidylserine IgG Ab B2GP1 dependent [Multiple of the median] in Serum
C1623609|PS IgG B2GP1 dep MoM Ser
C1623609|Phosphatidylserine Antibody.immunoglobulin G.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C1715010|Plasminogen activator tissue type:ACnc:Pt:PPP:Ord:Chromo
C1715010|Plasminogen activator tissue type [Presence] in Platelet poor plasma by Chromogenic method
C1715010|tPA PPP Ql Chro
C1715010|Plasminogen activator tissue type:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Chromogenic/Enzymatic Assay
C2360880|Coagulation tissue factor induced.factor substitution^after addition of normal plasma 1H post incubation separate tubes:Time:Pt:PPP:Qn:Coag
C2360880|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --with normal plasma 1H post incubation separate tubes
C2360880|Coagulation tissue factor induced.factor substitution^after addition of normal plasma 1 hour post incubation separate tubes:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2360880|PT NP 1h separate PPP
C2360097|Coagulation surface induced^post heparin adsorption:Time:Pt:PPP:Qn:Coag
C2360097|Coagulation surface induced^post heparin adsorption:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2360097|aPTT p heparin adsorption PPP
C2360097|aPTT in Platelet poor plasma by Coagulation assay --post heparin adsorption
C2361194|Clotting time.intrinsic coagulation system activated.heparin insensitive:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361194|Clotting time.intrinsic coagulation system activated.heparin insensitive:Time:Pt:Bld:Qn:Thromboelastography
C2361194|Clotting time.intrinsic coagulation system activated.heparin insensitive of Blood by Thromboelastography
C2361194|CT.heparin insens Bld TEG
C2361218|Maximum lysis.intrinsic coagulation system activated:LenFr:Pt:Bld:Qn:Thromboelastography
C2361218|Maximum lysis.intrinsic coagulation system activated [Length fraction] in Blood by Thromboelastography
C2361218|Maximum lysis.intrinsic coagulation system activated:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C2361218|ML.intrinsic LenFr Bld TEG
C1977665|Coagulation factor VIII activity actual/normal in Platelet poor plasma by Chromogenic method
C1977665|Coagulation factor VIII activity actual/Normal:RelACnc:Pt:PPP:Qn:Chromo
C1977665|Fact VIII Act/Nor PPP Chro
C1977665|Coagulation factor VIII activity actual/Normal:Relative Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1977547|Mixing studies:Imp:Pt:PPP:Nar
C1977547|Mixing studies PPP-Imp
C1977547|Mixing studies:Impression/interpretation of study:Point in time:Platelet poor plasma:Narrative
C1977547|Mixing studies [Interpretation] in Platelet poor plasma Narrative
C2733953|Platelet aggregation ADP induced ATP secretion [Presence] in Blood --5 umol/L
C2733953|PA ADP ATP secr 5 umol/L Bld Ql
C2733953|Platelet aggregation.adenosine diphosphate induced ATP secretion^5 umol/L:Presence:Point in time:Whole blood:Ordinal
C2733953|Platelet aggregation.adenosine diphosphate induced ATP secretion^5 umol/L:Pr:Pt:Bld:Ord
C2733954|Platelet aggregation.adenosine diphosphate induced^5 umol/L:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733954|Platelet aggregation.adenosine diphosphate induced^5 umol/L:RelACnc:Pt:Bld:Qn
C2733954|PA ADP 5 umol/L Bld
C2733954|Platelet aggregation ADP induced in Blood --5 umol/L
C2598683|Coagulation surface induced.lupus insensitive:Time:Pt:PPP:Qn:Coag
C2598683|Coagulation surface induced.lupus insensitive:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2598683|aPTT-LA insens PPP
C2598683|aPTT.lupus insensitive in Platelet poor plasma by Coagulation assay
C0551329|Phosphatidate Ab.IgM:ACnc:Pt:Ser:Qn
C0551329|Phosphatidate IgM Ser-aCnc
C0551329|Phosphatidate IgM Ab [Units/volume] in Serum
C0551329|Phosphatidate Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0943507|Antithrombin Ag actual/normal in Platelet poor plasma by Immunologic method
C0943507|AT III Ag Act/Nor PPP Imm
C0943507|Antithrombin Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0943507|Antithrombin Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1317033|Coagulation surface induced.lupus sensitive:Time:Pt:PPP^control:Qn:Coag
C1317033|Coagulation surface induced.lupus sensitive:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1317033|aPTT-LA Cont PPP
C1317033|aPTT.lupus sensitive in control Platelet poor plasma by Coagulation assay
C0482656|Coagulation factor XII activity:ACnc:Pt:PPP:Qn:Chromo
C0482656|Fact XII PPP Chro-aCnc
C0482656|Coagulation factor XII activity [Units/volume] in Platelet poor plasma by Chromogenic method
C0482656|Coagulation factor XII activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482728|Coagulation surface induced.hexagonal phase phospholipid:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482728|Coagulation surface induced.hexagonal phase phospholipid:Time:Pt:PPP:Qn:Coag
C0482728|aPTT W excess hexagonal phase phospholipid in Platelet poor plasma by Coagulation assay
C0482728|aPTT Hex PL PPP
C0482771|Prothrombin Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482771|Prothrom Ag PPP Imm-aCnc
C0482771|Prothrombin Ag:ACnc:Pt:PPP:Qn:Imm
C0482771|Prothrombin Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482708|Fibrinogen Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482708|Fibrinogen Ag:MCnc:Pt:PPP:Qn:Imm
C0482708|Fibrinogen Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482708|Fibrinogen Ag PPP Imm-mCnc
C0482712|Fibrinopeptide B beta (15-42) Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482712|Fibrinopeptide B beta (15-42) Ag:MCnc:Pt:PPP:Qn:Imm
C0482712|FpB Beta15-42 Ag PPP Imm-mCnc
C0482712|Fibrinopeptide B beta (15-42) Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0365323|Bleeding time:Time:Point in time:^Patient:Quantitative:Ivy
C0365323|Bleeding time by Ivy method
C0365323|Bleeding time:Time:Pt:^Patient:Qn:Ivy
C0365323|Bleeding time Patient Ivy
C0482652|Fact XI Ag Act/Nor PPP Imm
C0482652|Coagulation factor XI Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482652|Coagulation factor XI Ag actual/normal in Platelet poor plasma by Immunologic method
C0482652|Coagulation factor XI Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482655|Coagulation factor XII activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482655|Coagulation factor XII activity actual/normal in Platelet poor plasma by Coagulation assay
C0482655|Fact XII Act/Nor PPP
C0482655|Coagulation factor XII activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544093|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --30 minutes post XXX challenge
C1544093|Coagulation tissue factor induced^30M post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544093|Coagulation tissue factor induced^30 minutes post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544093|PT 30M p chal PPP
C1544550|PA Epineph 50 umol/L PRP-aCnc
C1544550|Platelet aggregation.epinephrine induced^50 umol/L:ACnc:Pt:PRP:Qn
C1544550|Platelet aggregation.epinephrine induced^50 umol/L:Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1544550|Platelet aggregation epinephrine induced [Units/volume] in Platelet rich plasma --50 umol/L
C2361208|MCF.heparin insens Bld TEG
C2361208|Maximum clot firmness.intrinsic coagulation system activated.heparin insensitive [Length] in Blood by Thromboelastography
C2361208|Maximum clot firmness.intrinsic coagulation system activated.heparin insensitive:Len:Pt:Bld:Qn:Thromboelastography
C2361208|Maximum clot firmness.intrinsic coagulation system activated.heparin insensitive:Length:Point in time:Whole blood:Quantitative:Thromboelastography
C1954800|Coagulation surface induced:Time:Pt:BldCRRT:Qn:Coag
C1954800|Coagulation surface induced:Time:Point in time:BldCRRT:Quantitative:Coagulation Assay
C1954800|aPTT BldCRRT
C1954800|aPTT in Blood drawn from CRRT circuit by Coagulation assay
C0365393|Deprecated Activated partial thrombplastin time (aPTT) in Blood by Coagulation assay
C0365393|Deprecated aPTT Plas Qn
C0365393|Coagulation surface induced:Time:Pt:Plas:Qn:Coag
C0365393|Coagulation surface induced:Time:Point in time:Plasma:Quantitative:Coagulation Assay
C0482673|Coagulation surface induced.factor substitution^20M post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C0482673|Coagulation surface induced.factor substitution^20 minutes post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482673|aPTT 20M NP PPP
C0482673|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --20M post incubation with normal plasma
C3259771|Clot angle:Angle:Pt:Bld:Qn:Thromboelastography
C3259771|Clot angle:Angle:Point in time:Whole blood:Quantitative:Thromboelastography
C3259771|Clot angle in Blood by Thromboelastography
C3259771|Clot angle Bld TEG
C2970621|Prothrombin time (PT) in Platelet poor plasma from Fetus by Coagulation assay
C2970621|Coagulation tissue factor induced:Time:Pt:PPP^fetus:Qn:Coag
C2970621|Coagulation tissue factor induced:Time:Point in time:Platelet poor plasma^Fetus:Quantitative:Coagulation Assay
C2970621|PT PPP Fetus
C2970622|Coagulation surface induced:Time:Pt:PPP^fetus:Qn:Coag
C2970622|Coagulation surface induced:Time:Point in time:Platelet poor plasma^Fetus:Quantitative:Coagulation Assay
C2970622|aPTT PPP Fetus
C2970622|aPTT in Platelet poor plasma from Fetus by Coagulation assay
C0482764|Protein C inhibitor [Mass/volume] in Platelet poor plasma by Immunologic method
C0482764|Protein C inhibitor:MCnc:Pt:PPP:Qn:Imm
C0482764|Prot C Inhib PPP Imm-mCnc
C0482764|Protein C inhibitor:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482763|Prot C CF PPP-aCnc
C0482763|Protein C cofactor:ACnc:Pt:PPP:Qn
C0482763|Protein C cofactor [Units/volume] in Platelet poor plasma
C0482763|Protein C cofactor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0485839|Cardiolipin Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C0485839|Cardiolipin IgM SerPl-aCnc
C0485839|Cardiolipin IgM Ab [Units/volume] in Serum or Plasma
C0485839|Cardiolipin Ab.IgM:ACnc:Pt:Ser/Plas:Qn
C0484862|Coagulation factor VI Ag:ACnc:Pt:Tiss:Ord:Immune stain
C0484862|Fact VI Ag Tiss Ql ImStn
C0484862|Coagulation factor VI Ag [Presence] in Tissue by Immune stain
C0484862|Coagulation factor VI Antigen:Arbitrary Concentration:Point in time:Tissue, unspecified:Ordinal:Immune stain
C0484864|Coagulation factor XIII Ag [Presence] in Tissue by Immune stain
C0484864|Fact XIII Ag Tiss Ql ImStn
C0484864|Coagulation factor XIII Ag:ACnc:Pt:Tiss:Ord:Immune stain
C0484864|Coagulation factor XIII Antigen:Arbitrary Concentration:Point in time:Tissue, unspecified:Ordinal:Immune stain
C0800001|FpB Beta1-42 Ag PPP Imm-aCnc
C0800001|Fibrinopeptide B beta (1-42) Ag:ACnc:Pt:PPP:Qn:Imm
C0800001|Fibrinopeptide B beta (1-42) Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0800001|Fibrinopeptide B beta (1-42) Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0803824|PA PPP-Imp
C0803824|Platelet aggregation:Imp:Pt:PPP:Nom
C0803824|Platelet aggregation:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal
C0803824|Platelet aggregation [Interpretation] in Platelet poor plasma
C0944229|Heparinoid [Units/volume] in Platelet poor plasma by Chromogenic method
C0944229|Heparinoid PPP Chro-aCnc
C0944229|Heparinoid:ACnc:Pt:PPP:Qn:Chromo
C0944229|Heparinoid:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0881644|Platelet aggregation epinephrine induced [Presence] in Platelet rich plasma
C0881644|Platelet aggregation.epinephrine induced:ACnc:Pt:PRP:Ord
C0881644|PA Epineph PRP Ql
C0881644|Platelet aggregation.epinephrine induced:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C1316137|Coagulation thrombin induced.factor substitution^immediately after addition of protamine sulfate:Time:Pt:PPP:Qn:Coag
C1316137|Thrombin time.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of protamine sulfate
C1316137|Coagulation thrombin induced.factor substitution^immediately after addition of protamine sulfate:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1316137|TT imm SO4 PPP
C1317032|Coagulation surface induced.lupus sensitive:Time:Pt:PPP:Qn:Coag
C1317032|Coagulation surface induced.lupus sensitive:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1317032|aPTT.lupus sensitive (LA screen)
C1317032|Screen aPTT
C0482695|Recalcification time in Platelet poor plasma by Coagulation assay
C0482695|Coagulation calcium ion induced:Time:Pt:PPP:Qn:Coag
C0482695|Coagulation calcium ion induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482695|Recal time PPP
C1316001|PA Rist hi dose PRP Cont
C1316001|Platelet aggregation ristocetin induced in control Platelet rich plasma --High dose
C1316001|Platelet aggregation.ristocetin induced^high dose:RelACnc:Pt:PRP^control:Qn
C1316001|Platelet aggregation.ristocetin induced^high dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma^Control:Quantitative
C1316021|PA Rist 900 ug/mL PRP
C1316021|Platelet aggregation ristocetin induced in Platelet rich plasma --900 ug/mL
C1316021|Platelet aggregation.ristocetin induced^900 ug/mL:RelACnc:Pt:PRP:Qn
C1316021|Platelet aggregation.ristocetin induced^900 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1114193|Coagulation surface induced.factor substitution^1H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1114193|Coagulation surface induced.factor substitution^1 hour post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1114193|aPTT 1h NP PPP
C1114193|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --1H post incubation with normal plasma
C0482631|Fact VIII Ab PPP Ql Chro
C0482631|Coagulation factor VIII Ab:ACnc:Pt:PPP:Ord:Chromo
C0482631|Coagulation factor VIII Ab [Presence] in Platelet poor plasma by Chromogenic method
C0482631|Coagulation factor VIII Antibody:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Chromogenic/Enzymatic Assay
C1113787|Cardiolipin Ab:ACnc:Pt:Ser:Ord
C1113787|Cardiolipin Ab Ser Ql
C1113787|Cardiolipin Ab [Presence] in Serum
C1113787|Cardiolipin Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C1544091|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --2 hours pre XXX challenge
C1544091|Coagulation tissue factor induced^2H pre XXX challenge:Time:Pt:PPP:Qn:Coag
C1544091|Coagulation tissue factor induced^2 hours pre XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544091|PT 2h pre chal PPP
C1544551|PA Epineph 100 umol/L PRP-aCnc
C1544551|Platelet aggregation.epinephrine induced^100 umol/L:ACnc:Pt:PRP:Qn
C1544551|Platelet aggregation epinephrine induced [Units/volume] in Platelet rich plasma --100 umol/L
C1544551|Platelet aggregation.epinephrine induced^100 umol/L:Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1717340|Beta 2 glycoprotein 1 IgG Ab [Units/volume] in Serum or Plasma by Immunoassay
C1717340|Beta 2 glycoprotein 1 Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:Enzyme Immunoassay
C1717340|B2 Glycoprot1 IgG SerPl EIA-aCnc
C1717340|Beta 2 glycoprotein 1 Ab.IgG:ACnc:Pt:Ser/Plas:Qn:EIA
C1830791|Coagulation thrombin induced.factor substitution^immediately after addition of bovine thrombin:Time:Pt:PPP:Qn:Coag
C1830791|Thrombin time.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of bovine thrombin
C1830791|Coagulation thrombin induced.factor substitution^immediately after addition of bovine thrombin:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1830791|TT imm Bovine Thrombin PPP
C1623606|PE IgA B2GP1 indep MoM Ser
C1623606|Phosphatidylethanolamine Ab.IgA.B2GP1 independent:MoM:Pt:Ser:Qn
C1623606|Phosphatidylethanolamine IgA Ab B2GP1 independent [Multiple of the median] in Serum
C1623606|Phosphatidylethanolamine Antibody.immunoglobulin A.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1624712|Phosphatidylserine IgM Ab B2GP1 dependent [Multiple of the median] in Serum
C1624712|Phosphatidylserine Ab.IgM.B2GP1 dependent:MoM:Pt:Ser:Qn
C1624712|PS IgM B2GP1 dep MoM Ser
C1624712|Phosphatidylserine Antibody.immunoglobulin M.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C1978233|vWF CBA Act/Nor PPP EIA
C1978233|von Willebrand factor.collagen binding activity actual/Normal:RelRto:Pt:PPP:Qn:EIA
C1978233|von Willebrand factor (vWf).collagen binding activity actual/normal in Platelet poor plasma by Immunoassay
C1978233|von Willebrand factor.collagen binding activity actual/Normal:Relative Ratio:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C1978986|Phosphoserine Ab.IgA:ACnc:Pt:Ser/Plas:Ord
C1978986|Phosphoserine IgA Ab [Presence] in Serum or Plasma
C1978986|Phosphoserine IgA SerPl Ql
C1978986|Phosphoserine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum/Plasma:Ordinal
C1978990|Phosphoethanolamine Ab.IgM:ACnc:Pt:Ser/Plas:Ord
C1978990|Phosphoethanolamine IgM Ab [Presence] in Serum or Plasma
C1978990|PETN IgM SerPl Ql
C1978990|Phosphoethanolamine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum/Plasma:Ordinal
C0482770|Prot S PPP Chro-aCnc
C0482770|Protein S [Units/volume] in Platelet poor plasma by Chromogenic method
C0482770|Protein S:ACnc:Pt:PPP:Qn:Chromo
C0482770|Protein S:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482767|Protein S.free:ACnc:Pt:PPP:Qn:Coag
C0482767|Prot S Free PPP-aCnc
C0482767|Protein S Free [Units/volume] in Platelet poor plasma by Coagulation assay
C0482767|Protein S.free:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482737|tPA Ag 20M PPP Imm-mCnc
C0482737|Plasminogen activator tissue type Ag^20M post venistasis:MCnc:Pt:PPP:Qn:Imm
C0482737|Plasminogen activator tissue type Ag [Mass/volume] in Platelet poor plasma by Immunologic method --20 minutes post venistasis
C0482737|Plasminogen activator tissue type Antigen^20 minutes post venistasis:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0486261|Deprecated tPA 20M PPP-mCnc
C0486261|Plasminogen activator tissue type^20M post venistasis:MCnc:Pt:PPP:Qn:Enzy
C0486261|Deprecated Plasminogen activator tissue type [Units/volume] in Platelet poor plasma by Chromogenic method --20 minutes post venistasis
C0486261|Plasminogen activator tissue type^20 minutes post venistasis:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Enzy
C2733741|PA Coll ATP secr 5 ug/mL Bld
C2733741|Platelet aggregation.collagen induced ATP secretion^5 ug/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733741|Platelet aggregation collagen induced ATP secretion in Blood --5 ug/mL
C2733741|Platelet aggregation.collagen induced ATP secretion^5 ug/mL:RelACnc:Pt:Bld:Qn
C0484866|Coagulation reptilase induced:Time:Pt:PPP:Qn:Tilt tube
C0484866|Deprecated Reptilase PPP Qn
C0484866|Deprecated Reptilase time in Platelet poor plasma by Coagulation assay
C0484866|Coagulation reptilase induced:Time:Point in time:Platelet poor plasma:Quantitative:Tilt tube
C3172627|Coagulation surface induced actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3172627|Coagulation surface induced actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3172627|aPTT Act/Nor PPP
C3172627|aPTT actual/normal in Platelet poor plasma by Coagulation assay
C0482755|Platelet factor 4 [Units/volume] in Platelet poor plasma
C0482755|Platelet factor 4:ACnc:Pt:PPP:Qn
C0482755|PF4 PPP-aCnc
C0482755|Platelet factor 4:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C3481505|Coagulation thrombin induced actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3481505|Coagulation thrombin induced actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3481505|Thrombin time/normal
C3481505|Thrombin time actual/Normal
C0800000|Fibrinopeptide B beta (1-14) Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0800000|Fibrinopeptide B beta (1-14) Ag:ACnc:Pt:PPP:Qn:Imm
C0800000|FpB Beta1-14 Ag PPP Imm-aCnc
C0800000|Fibrinopeptide B beta (1-14) Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0800002|Fibrinopeptide B beta (15-42) Ag:ACnc:Pt:PPP:Qn:Imm
C0800002|Fibrinopeptide B beta (15-42) Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0800002|FpB Beta15-42 Ag PPP Imm-aCnc
C0800002|Fibrinopeptide B beta (15-42) Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0798529|Coagulation dilute Russell viper venom induced actual/Normal:ACnc:Pt:PPP:Ord:Coag
C0798529|Coagulation dilute Russell viper venom induced actual/Normal:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C0798529|dRVVT Act/Nor PPP Ql
C0798529|dRVVT actual/normal [Presence] in Platelet poor plasma by Coagulation assay
C0550841|Heparin [Units/volume] in Platelet poor plasma
C0550841|Heparin:ACnc:Pt:PPP:Qn
C0550841|Heparin PPP-aCnc
C0550841|Heparin:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0482657|Coagulation factor XII Ag:ACnc:Pt:PPP:Qn:Imm
C0482657|Fact XII Ag PPP Imm-aCnc
C0482657|Coagulation factor XII Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482657|Coagulation factor XII Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1316348|Coagulation tissue factor induced.factor substitution^2H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1316348|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --2H post incubation with 1:4 normal plasma
C1316348|Coagulation tissue factor induced.factor substitution^2 hours post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1316348|PT 2h p 1:4 NP PPP
C0482713|FpB Beta43-47 Ag PPP Imm-mCnc
C0482713|Fibrinopeptide B beta (43-47) Ag:MCnc:Pt:PPP:Qn:Imm
C0482713|Fibrinopeptide B beta (43-47) Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482713|Fibrinopeptide B beta (43-47) Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482638|Coagulation factor VIII Ag:MCnc:Pt:PPP:Qn:Imm
C0482638|Fact VIII Ag PPP Imm-mCnc
C0482638|Coagulation factor VIII Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482638|Coagulation factor VIII Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1526524|Fibrinopeptide A:MCnc:Pt:Urine:Qn
C1526524|Fibrinopeptide A [Mass/volume] in Urine
C1526524|FpA Ur-mCnc
C1526524|Fibrinopeptide A:Mass Concentration:Point in time:Urine:Quantitative
C1717468|Cardiolipin Ab [Presence] in Serum by Immunoassay
C1717468|Cardiolipin Ab Ser Ql EIA
C1717468|Cardiolipin Ab:ACnc:Pt:Ser:Ord:EIA
C1717468|Cardiolipin Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal:Enzyme Immunoassay
C1624148|Fibrinogen Ag:MCnc:Pt:PPP:Qn:Nephelometry
C1624148|Fibrinogen Ag [Mass/volume] in Platelet poor plasma by Nephlometry
C1624148|Fibrinogen Ag PPP Neph-mCnc
C1624148|Fibrinogen Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Nephelometry
C1624695|Heparin [Units/volume] in Platelet poor plasma by Chromogenic method
C1624695|Heparin PPP Chro-aCnc
C1624695|Heparin:ACnc:Pt:PPP:Qn:Chromo
C1624695|Heparin:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C2359912|PS IgM Titr Ser IF
C2359912|Phosphatidylserine Ab.IgM:Titr:Pt:Ser:Qn:IF
C2359912|Phosphatidylserine IgM Ab [Titer] in Serum by Immunofluorescence
C2359912|Phosphatidylserine Antibody.immunoglobulin M:Dilution Factor (Titer):Point in time:Serum:Quantitative:Immune Fluorescence
C0367396|Cardiolipin IgA Ser EIA-aCnc
C0367396|Cardiolipin Ab.IgA:ACnc:Pt:Ser:Qn:EIA
C0367396|Cardiolipin IgA Ab [Units/volume] in Serum by Immunoassay
C0367396|Cardiolipin Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1954167|von Willebrand evaluation:Imp:Pt:PPP:Nom
C1954167|von Willebrand eval PPP-Imp
C1954167|von Willebrand evaluation:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal
C1954167|von Willebrand evaluation [Interpretation] in Platelet poor plasma
C2713266|Deprecated Dilute Russell viper venom time (dRVVT) in Platelet poor plasma by Coagulation assay
C2713266|Deprecated dRVV Tme Plas Qn
C2713266|Coagulation dilute Russell viper venom induced:Time:Pt:Plas:Qn:Coag
C2713266|Coagulation dilute Russell viper venom induced:Time:Point in time:Plasma:Quantitative:Coagulation Assay
C0482688|Deprecated PT imm NP PPP Cont Qn
C0482688|Deprecated Prothrombin time (PT) factor substitution in Platelet poor plasma from control by Coagulation assay --immediately after addition of normal plasma
C0482688|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP^control:Qn:Tilt tube
C0482688|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Tilt tube
C3481475|Coagulation surface induced.lupus sensitive.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3481475|Coagulation surface induced.lupus sensitive.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C3481475|aPTT-LA imm NP PPP
C3481475|aPTT.lupus sensitive.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C3262763|Coagulation dilute Russell viper venom induced.excess phospholipid actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3262763|Coagulation dilute Russell viper venom induced.excess phospholipid actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3262763|Confirm dRVVT/normal
C3262763|dRVVT W excess phospholipid actual/normal (normalized LA confirm)
C0550589|Coagulation surface induced^3rd specimen:Time:Pt:PPP:Qn:Coag
C0550589|Coagulation surface induced^3rd specimen:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0550589|aPTT sp3 PPP
C0550589|aPTT in Platelet poor plasma by Coagulation assay --3rd specimen
C0551335|Phosphatidylethanolamine IgM Ab [Units/volume] in Serum
C0551335|Phosphatidylethanolamine Ab.IgM:ACnc:Pt:Ser:Qn
C0551335|PE IgM Ser-aCnc
C0551335|Phosphatidylethanolamine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0803789|Antithrombin:Imp:Pt:PPP:Nom
C0803789|AT III PPP-Imp
C0803789|Antithrombin:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal
C0803789|Antithrombin [Interpretation] in Platelet poor plasma
C0803828|TT Bld-Imp
C0803828|Coagulation thrombin induced:Imp:Pt:Bld:Nom
C0803828|Coagulation thrombin induced:Impression/interpretation of study:Point in time:Whole blood:Nominal
C0803828|Thrombin time [Interpretation] in Blood
C0364116|Bradykinin SerPl-mCnc
C0364116|Bradykinin:MCnc:Pt:Ser/Plas:Qn
C0364116|Bradykinin [Mass/volume] in Serum or Plasma
C0364116|Bradykinin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0800569|Phosphatidylethanolamine Ab.IgM:ACnc:Pt:Ser:Ord
C0800569|Phosphatidylethanolamine IgM Ab [Presence] in Serum
C0800569|PE IgM Ser Ql
C0800569|Phosphatidylethanolamine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal
C0944744|Fibrin degradation products [Presence] in Blood by Agglutination
C0944744|Fibrin degradation products:ACnc:Pt:Bld:Ord:Aggl
C0944744|FDP Bld Ql Aggl
C0944744|Fibrin degradation products:Arbitrary Concentration:Point in time:Whole blood:Ordinal:Agglutination
C1317031|Lupus anticoagulant neutralization.high phospholipid.factor substitution^immediately after 1:2 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1317031|Lupus anticoagulant neutralization high phospholipid.factor substitution [Time] in Platelet poor plasma by Coagulation assay --immediately after 1:2 addition of normal plasma
C1317031|Lupus anticoagulant neutralization.high phospholipid.factor substitution^immediately after 1:2 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1317031|LA Nt HPL imm 1:2 NP PPP
C1316357|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --1H post incubation with 1:4 normal plasma
C1316357|Coagulation tissue factor induced.factor substitution^1H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1316357|Coagulation tissue factor induced.factor substitution^1 hour post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1316357|PT 1h p 1:4 NP PPP
C1542959|Fibrin D-dimer:Titr:Pt:PPP:Qn
C1542959|D Dimer Titr PPP
C1542959|Fibrin D-dimer [Titer] in Platelet poor plasma
C1542959|Fibrin D-dimer:Dilution Factor (Titer):Point in time:Platelet poor plasma:Quantitative
C1508152|Coagulation surface induced^1H post incubation:Time:Pt:PPP^pool:Qn:Coag
C1508152|Coagulation surface induced^1 hour post incubation:Time:Point in time:Platelet poor plasma^Pool specimen:Quantitative:Coagulation Assay
C1508152|aPTT 1h p Inc Pool PPP
C1508152|aPTT in Pooled Platelet poor plasma by Coagulation assay --1 hour post incubation
C1625223|PE IgA B2GP1 dep MoM Ser
C1625223|Phosphatidylethanolamine IgA Ab B2GP1 dependent [Multiple of the median] in Serum
C1625223|Phosphatidylethanolamine Ab.IgA.B2GP1 dependent:MoM:Pt:Ser:Qn
C1625223|Phosphatidylethanolamine Antibody.immunoglobulin A.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C2359872|Thrombin time.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of XXX
C2359872|Coagulation thrombin induced.factor substitution^immediately after addition of XXX:Time:Pt:PPP:Qn:Coag
C2359872|Coagulation thrombin induced.factor substitution^immediately after addition of XXX:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2359872|TT imm XXX PPP
C2361166|PK activity Act/Nor PPP
C2361166|Prekallikrein (Fletcher Factor) activity actual/normal in Platelet poor plasma by Coagulation assay
C2361166|Prekallikrein activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C2361166|Prekallikrein activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2361180|Coagulation surface induced^after addition of protein C activator/Coagulation surface induced:Time Ratio:Point in time:Platelet poor plasma:Quantitative:COAGULATION ASSAY
C2361180|Coagulation surface induced^after addition of protein C activator/Coagulation surface induced:TRto:Pt:PPP:Qn:Coag
C2361180|aPTTprotein C activator/aPTT PPP
C2361180|Activated partial thromboplastin time (aPTT) in Platelet poor plasma by Coagulation assay -- after addition of protein C activator/Activated partial thromboplastin time (aPTT)
C2361186|Clot formation.intrinsic coagulation system activated:Time:Pt:Bld:Qn:Thromboelastography
C2361186|Clot formation.intrinsic coagulation system activated [Time] in Blood by Thromboelastography
C2361186|Clot formation.intrinsic coagulation system activated:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361186|CFT.intrinsic Bld TEG
C2359886|Coagulation tissue factor induced.factor substitution^after addition of 1:4 normal plasma 1H post incubation separate tubes:Time:Pt:PPP:Qn:Coag
C2359886|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --with 1:4 normal plasma 1H post incubation separate tubes
C2359886|Coagulation tissue factor induced.factor substitution^after addition of 1:4 normal plasma 1 hour post incubation separate tubes:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2359886|PT 1:4 NP 1h separate PPP
C1978984|PETN IgA SerPl Ql
C1978984|Phosphoethanolamine IgA Ab [Presence] in Serum or Plasma
C1978984|Phosphoethanolamine Ab.IgA:ACnc:Pt:Ser/Plas:Ord
C1978984|Phosphoethanolamine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum/Plasma:Ordinal
C0482690|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Tilt tube
C0482690|Deprecated PT imm NP PPP Qn
C0482690|Deprecated Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C0482690|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Tilt tube
C0365405|Prothrombin time (PT) in Blood by Coagulation assay
C0365405|Coagulation tissue factor induced:Time:Pt:Bld:Qn:Coag
C0365405|Coagulation tissue factor induced:Time:Point in time:Whole blood:Quantitative:Coagulation Assay
C0365405|PT Bld
C0482739|Plasminogen activator inhibitor 1 Ag:ACnc:Pt:PPP:Qn:Imm
C0482739|PAI1 Ag PPP Imm-aCnc
C0482739|Plasminogen activator inhibitor 1 Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482739|Plasminogen activator inhibitor 1 Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482741|PAI2 Ag PPP Imm-aCnc
C0482741|Plasminogen activator inhibitor 2 Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482741|Plasminogen activator inhibitor 2 Ag:ACnc:Pt:PPP:Qn:Imm
C0482741|Plasminogen activator inhibitor 2 Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C2733964|PA Thromb ATP secr 5 U/mL Bld
C2733964|Platelet aggregation.thrombin induced ATP secretion^5 U/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733964|Platelet aggregation.thrombin induced ATP secretion^5 U/mL:RelACnc:Pt:Bld:Qn
C2733964|Platelet aggregation thrombin induced ATP secretion in Blood --5 U/mL
C2733965|PA Thromb ATP secr 1 U/mL Bld Ql
C2733965|Platelet aggregation thrombin induced ATP secretion [Presence] in Blood --1 U/mL
C2733965|Platelet aggregation.thrombin induced ATP secretion^1 U/mL:ACnc:Pt:Bld:Ord
C2733965|Platelet aggregation.thrombin induced ATP secretion^1 U/mL:Arbitrary Concentration:Point in time:Whole blood:Ordinal
C2598679|PA Coll 8.0 ug/mL PRP
C2598679|Platelet aggregation collagen induced in Platelet rich plasma --8.0 ug/mL
C2598679|Platelet aggregation.collagen induced^8.0 ug/mL:RelACnc:Pt:PRP:Qn
C2598679|Platelet aggregation.collagen induced^8.0 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C3259334|MCF Heparinase Bld TEG
C3259334|Maximum clot firmness^after addition of heparinase:Len:Pt:Bld:Qn:Thromboelastography
C3259334|Maximum clot firmness [Length] in Blood by Thromboelastography --after addition of heparinase
C3259334|Maximum clot firmness^after addition of heparinase:Length:Point in time:Whole blood:Quantitative:Thromboelastography
C0365494|PA Ca Ionoph PRP
C0365494|Platelet aggregation.calcium ionophore induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0365494|Platelet aggregation calcium ionophore induced in Platelet rich plasma
C0365494|Platelet aggregation.calcium ionophore induced:RelACnc:Pt:PRP:Qn
C3699643|Apixaban PPP Chro-mCnc
C3699643|Apixaban [Mass/volume] in Platelet poor plasma by Chromogenic method
C3699643|Apixaban:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3699643|Apixaban:MCnc:Pt:PPP:Qn:Chromo
C3262207|von Willebrand factor.activity actual/Normal:RelRto:Pt:PPP:Qn:Imm
C3262207|von Willebrand factor (vWf).activity actual/normal in Platelet poor plasma by Immunologic method
C3262207|von Willebrand factor.activity actual/Normal:Relative Ratio:Point in time:Platelet poor plasma:Quantitative:Imm
C3262207|vWf:Ac Act/Nor PPP Imm
C1973915|Streptokinase Ab &#x7C; bld-ser-plas
C0798528|Coagulation dilute Russell viper venom induced actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0798528|Coagulation dilute Russell viper venom induced actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0798528|Screen dRVVT/normal
C0798528|dRVVT actual/normal (normalized LA screen)
C0796782|Factor inhibitor XXX [Units/volume] in Platelet poor plasma by Coagulation assay
C0796782|Fact Inhib XXX PPP-aCnc
C0796782|Factor inhibitor XXX:ACnc:Pt:PPP:Qn:Coag
C0796782|Factor inhibitor XXX:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0803799|Fibrinogen PPP-Imp
C0803799|Fibrinogen:Imp:Pt:PPP:Nom
C0803799|Fibrinogen:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal
C0803799|Fibrinogen [Interpretation] in Platelet poor plasma
C0943509|Coagulation factor VII+Coagulation factor X activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0943509|Coagulation factor VII+Coagulation factor X actual/normal in Platelet poor plasma by Coagulation assay
C0943509|Fact VII+Fact X Act/Nor PPP
C0943509|Coagulation factor VII+Coagulation factor X activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0944233|Coagulation factor X activated actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C0944233|Coagulation factor X activated actual/normal in Platelet poor plasma by Chromogenic method
C0944233|Fact Xa Act/Nor PPP Chro
C0944233|Coagulation factor X activated actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0881646|PA Rist PRP Ql
C0881646|Platelet aggregation ristocetin induced [Presence] in Platelet rich plasma
C0881646|Platelet aggregation.ristocetin induced:ACnc:Pt:PRP:Ord
C0881646|Platelet aggregation.ristocetin induced:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C0482658|Coagulation factor XII Ag actual/normal in Platelet poor plasma by Immunologic method
C0482658|Coagulation factor XII Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482658|Fact XII Ag Act/Nor PPP Imm
C0482658|Coagulation factor XII Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482724|Kininogen.high molecular weight:MCnc:Pt:PPP:Qn:Imm
C0482724|HMWK PPP Imm-mCnc
C0482724|Kininogen HMW [Mass/volume] in Platelet poor plasma by Immunologic method
C0482724|Kininogen.high molecular weight:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482701|Fibrin Frg PPP IEP
C0482701|Fibrin fragments [Identifier] in Platelet poor plasma by Immunoelectrophoresis
C0482701|Fibrin fragments:Prid:Pt:PPP:Nom:Immunoelectrophoresis
C0482701|Fibrin fragments:Presence or Identity:Point in time:Platelet poor plasma:Nominal:Immunoelectrophoresis
C1316349|Coagulation tissue factor induced.factor substitution^2H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316349|Coagulation tissue factor induced.factor substitution^2 hours post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316349|Prothrombin time (PT) factor substitution in control Platelet poor plasma by Coagulation assay --2H post incubation with 1:4 normal plasma
C1316349|PT 2h p 1:4 NP Cont PPP
C1316393|aPTT W excess hexagonal phospholipid (StaClot LA confirm)
C1316393|Confirm aPTT StaClot
C1316393|Coagulation surface induced.hexagonal phase phospholipid:ACnc:Pt:PPP:Ord
C1316393|Coagulation surface induced.hexagonal phase phospholipid:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C0365324|Cardiolipin Ab:ACnc:Pt:Ser:Qn:EIA
C0365324|Cardiolipin Ab Ser EIA-aCnc
C0365324|Cardiolipin Ab [Units/volume] in Serum by Immunoassay
C0365324|Cardiolipin Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0482608|Coagulation activated:Time:Pt:Bld:Qn:Coag
C0482608|Activated clotting time in Blood by Coagulation assay
C0482608|Coagulation activated:Time:Point in time:Whole blood:Quantitative:Coagulation Assay
C0482608|ACT Bld
C0482611|Fact IX Act/Nor PPP
C0482611|Coagulation factor IX activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482611|Coagulation factor IX activity actual/normal in Platelet poor plasma by Coagulation assay
C0482611|Coagulation factor IX activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482625|Fact VII Ag PPP Imm-aCnc
C0482625|Coagulation factor VII Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482625|Coagulation factor VII Ag:ACnc:Pt:PPP:Qn:Imm
C0482625|Coagulation factor VII Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1526521|Capillary fragility:ACnc:Pt:^Patient:Ord
C1526521|Capillary fragility [Presence]
C1526521|Capillary Fragility Patient Ql
C1526521|Capillary fragility:Arbitrary Concentration:Point in time:^Patient:Ordinal
C1544096|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --2 hours post XXX challenge
C1544096|Coagulation tissue factor induced^2H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544096|Coagulation tissue factor induced^2 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544096|PT 2h p chal PPP
C1544602|Lupus anticoagulant neutralization.platelet:ACnc:Pt:PPP:Ord:Coag
C1544602|Lupus anticoagulant neutralization platelet [Presence] in Platelet poor plasma by Coagulation assay
C1544602|Lupus anticoagulant neutralization.platelet:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C1544602|LA Nt Platelet PPP Ql
C1646771|Phosphatidylcholine IgA Ab B2GP1 independent [Multiple of the median] in Serum
C1646771|PC IgA B2GP1 indep MoM Ser
C1646771|Phosphatidylcholine Ab.IgA.B2GP1 independent:MoM:Pt:Ser:Qn
C1646771|Phosphatidylcholine Antibody.immunoglobulin A.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1624711|Phosphatidylserine Ab.IgG.B2GP1 independent:MoM:Pt:Ser:Qn
C1624711|Phosphatidylserine IgG Ab B2GP1 independent [Multiple of the median] in Serum
C1624711|PS IgG B2GP1 indep MoM Ser
C1624711|Phosphatidylserine Antibody.immunoglobulin G.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1704394|Coagulation dilute Russell viper venom induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:COAGULATION ASSAY
C1704394|Coagulation dilute Russell viper venom induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1704394|dRVVT factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C1704394|dRVVT imm NP PPP
C1715216|Beta 2 glycoprotein 1 Ab.IgA:ACnc:Pt:Ser:Ord
C1715216|Beta 2 glycoprotein 1 IgA Ab [Presence] in Serum
C1715216|B2 Glycoprot1 IgA Ser Ql
C1715216|Beta 2 glycoprotein 1 Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Ordinal
C2361741|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after 1:4 addition of normal plasma
C2361741|Coagulation tissue factor induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2361741|Coagulation tissue factor induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2361741|PT imm 1:4 NP PPP
C1953434|Coagulation kaolin induced:ACnc:Pt:Bld:Qn
C1953434|Kaolin activated time [Units/volume] in Blood
C1953434|Coagulation kaolin induced:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C1953434|KCT Bld-aCnc
C2924051|Coagulation dilute Russell viper venom induced.factor substitution^2H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2924051|Coagulation dilute Russell viper venom induced.factor substitution^2 hours post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2924051|dRVVT factor substitution in Platelet poor plasma by Coagulation assay --2H post incubation with normal plasma
C2924051|dRVVT 2h NP PPP
C2733955|Platelet aggregation.adenosine diphosphate induced^10 umol/L:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733955|Platelet aggregation ADP induced in Blood --10 umol/L
C2733955|Platelet aggregation.adenosine diphosphate induced^10 umol/L:RelACnc:Pt:Bld:Qn
C2733955|PA ADP 10 umol/L Bld
C0482750|Plasminogen activator tissue type^10M post venistasis:ACnc:Pt:PPP:Qn:Chromo
C0482750|Plasminogen activator tissue type [Units/volume] in Platelet poor plasma by Chromogenic method --10 minutes post venistasis
C0482750|tPA 10M PPP Chro-aCnc
C0482750|Plasminogen activator tissue type^10 minutes post venistasis:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0005789|Blood Coagulation Factor
C0005789|Blood Coagulation Factors
C0005789|Factor, Blood Coagulation
C0005789|Factors, Blood Coagulation
C0005789|clotting factor
C0005789|COAG FACTORS
C0005789|BLOOD COAG FACTOR
C0005789|COAG FACTOR
C0005789|COAG FACTORS BLOOD
C0005789|BLOOD COAG FACTORS
C0005789|FACTORS COAG
C0005789|FACTOR COAG
C0005789|COAG FACTOR BLOOD
C0005789|Coagulation Factors
C0005789|Factors, Coagulation
C0005789|Coagulation Factor
C0005789|Blood Coagulation Factors [Chemical/Ingredient]
C0005789|Coagulation Factor, Blood
C0005789|Factor, Coagulation
C0005789|Coagulation Factors, Blood
C0005789|Clotting factors
C0005789|Coagulation factor (substance)
C0005789|Blood clotting factor
C0005789|Blood clotting factor (product)
C0005789|Coagulation factor, NOS
C0005789|Blood clotting factor (substance)
C0799301|B2 Glycoprot1 IgM Ser-aCnc
C0799301|Beta 2 glycoprotein 1 IgM Ab [Units/volume] in Serum
C0799301|Beta 2 glycoprotein 1 Ab.IgM:ACnc:Pt:Ser:Qn
C0799301|Beta 2 glycoprotein 1 Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0797429|PC IgM Ser Ql
C0797429|Phosphatidylcholine Ab.IgM:ACnc:Pt:Ser:Ord
C0797429|Phosphatidylcholine IgM Ab [Presence] in Serum
C0797429|Phosphatidylcholine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal
C0551333|PE IgA Ser-aCnc
C0551333|Phosphatidylethanolamine Ab.IgA:ACnc:Pt:Ser:Qn
C0551333|Phosphatidylethanolamine IgA Ab [Units/volume] in Serum
C0551333|Phosphatidylethanolamine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C0943514|Protein C actual/normal in Platelet poor plasma by Coagulation assay
C0943514|Prot C Act/Nor PPP
C0943514|Protein C actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0943514|Protein C actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0943661|Fibrinogen fragments [Mass/volume] in Urine by Latex agglutination
C0943661|Fibrinogen Frg Ur LA-mCnc
C0943661|Fibrinogen fragments:MCnc:Pt:Urine:Qn:LA
C0943661|Fibrinogen fragments:Mass Concentration:Point in time:Urine:Quantitative:Latex Agglutination
C0941530|Coagulation calcium ion induced:Time:Pt:PPP^control:Qn:Coag
C0941530|Coagulation calcium ion induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0941530|Recalcification time in control Platelet poor plasma by Coagulation assay
C0941530|Recal time Cont PPP
C1316135|Platelet aggregation.collagen induced lag^high dose:Time:Pt:PRP^control:Qn
C1316135|Platelet aggregation.collagen induced lag^high dose:Time:Point in time:Platelet rich plasma^Control:Quantitative
C1316135|Platelet aggregation collagen induced lag [Time] in control Platelet rich plasma --High dose
C1316135|PA Coll Lag time hi dose Cont PRP
C0482726|LMWK PPP Imm-mCnc
C0482726|Kininogen.low molecular weight:MCnc:Pt:PPP:Qn:Imm
C0482726|Kininogen LMW [Mass/volume] in Platelet poor plasma by Immunologic method
C0482726|Kininogen.low molecular weight:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1315995|Coagulation reptilase induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1315995|Reptilase time.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C1315995|Coagulation reptilase induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1315995|Reptilase time imm NP PPP
C1316020|PA Rist 1200 ug/mL PRP
C1316020|Platelet aggregation.ristocetin induced^1200 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1316020|Platelet aggregation.ristocetin induced^1200 ug/mL:RelACnc:Pt:PRP:Qn
C1316020|Platelet aggregation ristocetin induced in Platelet rich plasma --1200 ug/mL
C2363272|Coagulation factor VIII Ag [Units/volume] in Platelet poor plasma by Immunologic method
C2363272|Fact VIII Ag PPP Imm-aCnc
C2363272|Coagulation factor VIII Ag:ACnc:Pt:PPP:Qn:Imm
C2363272|Coagulation factor VIII Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482639|Coagulation factor X inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482639|Fact X Inhib PPP-aCnc
C0482639|Coagulation factor X inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482639|Coagulation factor X inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1114118|Deprecated Fibrin D-dimer:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C1114118|Fibrin D-dimer:MCnc:Pt:PPP:Qn
C1114118|Deprecated D Dimer PPP-mCnc
C1114118|Deprecated Fibrin D-dimer
C1114118|Fibrin D-dimer:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C1544097|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --3 hours post XXX challenge
C1544097|Coagulation tissue factor induced^3H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544097|Coagulation tissue factor induced^3 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544097|PT 3h p chal PPP
C1625224|PE IgM B2GP1 dep MoM Ser
C1625224|Phosphatidylethanolamine Ab.IgM.B2GP1 dependent:MoM:Pt:Ser:Qn
C1625224|Phosphatidylethanolamine IgM Ab B2GP1 dependent [Multiple of the median] in Serum
C1625224|Phosphatidylethanolamine Antibody.immunoglobulin M.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C1624706|Fibrin D-dimer DDU [Mass/volume] in Cerebral spinal fluid by Latex agglutination
C1624706|D dimer DDU CSF LA-mCnc
C1624706|Fibrin D-dimer DDU:MCnc:Pt:CSF:Qn:LA
C1624706|Fibrin D-dimer DDU:Mass Concentration:Point in time:Cerebral spinal fluid:Quantitative:Latex Agglutination
C2361168|Prothrombin time (PT) PIVKA sensitive actual/normal in Capillary blood by Coagulation assay
C2361168|PT PIVKA sensitive Act/Nor BldC
C2361168|Coagulation tissue factor induced.PIVKA sensitive actual/Normal:RelTime:Pt:BldC:Qn:Coag
C2361168|Coagulation tissue factor induced.PIVKA sensitive actual/Normal:Relative Time:Point in time:Blood capillary:Quantitative:Coagulation Assay
C2361212|Maximum lysis:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C2361212|ML LenFr Bld TEG
C2361212|Maximum lysis:LenFr:Pt:Bld:Qn:Thromboelastography
C2361212|Maximum lysis [Length fraction] in Blood by Thromboelastography
C1978758|Coagulation surface induced:Time:Pt:PPP^pool:Qn:Coag
C1978758|Coagulation surface induced:Time:Point in time:Platelet poor plasma^Pool specimen:Quantitative:Coagulation Assay
C1978758|aPTT Pool PPP
C1978758|aPTT in Pooled Platelet poor plasma by Coagulation assay
C1954262|Fibrinogen:MCnc:Pt:PPP:Qn:Coag.derived
C1954262|Fibrinogen PPP Coag.derived-mCnc
C1954262|Fibrinogen [Mass/volume] in Platelet poor plasma by Coagulation.derived
C1954262|Fibrinogen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay.derived
C0482686|Deprecated PT PPP Qn
C0482686|Deprecated Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --20M post incubation with normal plasma
C0482686|Coagulation tissue factor induced.factor substitution^20 minutes post incubation.37 deg c after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Tilt tube
C0482686|Coagulation tissue factor induced.factor substitution^20M post incubation.37 deg c after addition of normal plasma:Time:Pt:PPP:Qn:Tilt tube
C2599018|Platelet aggregation ADP induced [Units/volume] in Blood
C2599018|PA ADP Bld-aCnc
C2599018|Platelet aggregation.adenosine diphosphate induced:ACnc:Pt:Bld:Qn
C2599018|Platelet aggregation.adenosine diphosphate induced:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2923557|Coagulation surface induced.lupus sensitive.factor substitution^2 hours post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2923557|Coagulation surface induced.lupus sensitive.factor substitution^2H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2923557|aPTT-LA 2h NP PPP
C2923557|aPTT.lupus sensitive.factor substitution in Platelet poor plasma by Coagulation assay --2H post incubation with normal plasma
C2970085|Coagulation ecarin induced:Time:Pt:PPP:Qn:Coag
C2970085|Ecarin clotting time (ECT) [Time] in Platelet poor plasma by Coagulation assay
C2970085|Coagulation ecarin induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2970085|ECT PPP
C0482759|Protein C [Units/volume] in Platelet poor plasma by Coagulation assay
C0482759|Protein C:ACnc:Pt:PPP:Qn:Coag
C0482759|Prot C PPP-aCnc
C0482759|Protein C:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0797367|Thrombin antithrombin complex Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0797367|TAT Ag PPP Imm-mCnc
C0797367|Thrombin antithrombin complex Ag:MCnc:Pt:PPP:Qn:Imm
C0797367|Thrombin antithrombin complex Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0551328|Phosphatidate Ab.IgG:ACnc:Pt:Ser:Qn
C0551328|Phosphatidate IgG Ser-aCnc
C0551328|Phosphatidate IgG Ab [Units/volume] in Serum
C0551328|Phosphatidate Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0551338|PG IgM Ser-aCnc
C0551338|Phosphatidylglycerol Ab.IgM:ACnc:Pt:Ser:Qn
C0551338|Phosphatidylglycerol IgM Ab [Units/volume] in Serum
C0551338|Phosphatidylglycerol Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0801387|Protein S Ag/Coagulation factor VII Ag:MRto:Pt:PPP:Qn:Coag
C0801387|Protein S Ag/Coagulation factor VII Ag Ag [Mass Ratio] in Platelet poor plasma by Coagulation assay
C0801387|Prot S Ag/Fact VII Ag PPP
C0801387|Protein S Antigen/Coagulation factor VII Antigen:Mass Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0881645|PA Coll PRP Ql
C0881645|Platelet aggregation.collagen induced:ACnc:Pt:PRP:Ord
C0881645|Platelet aggregation collagen induced [Presence] in Platelet rich plasma
C0881645|Platelet aggregation.collagen induced:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C1316136|PA Rist + Cont PPP PRP
C1316136|Platelet aggregation.ristocetin+Control PPP induced in Platelet rich plasma
C1316136|Platelet aggregation.ristocetin+Control PPP induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1316136|Platelet aggregation.ristocetin+Control PPP induced:RelACnc:Pt:PRP:Qn
C1369551|Coagulation tissue factor induced.factor substitution^immediately after addition of factor X depleted plasma:Time:Pt:PPP:Qn:Coag
C1369551|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor X depleted plasma
C1369551|Coagulation tissue factor induced.factor substitution^immediately after addition of factor X depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1369551|PT imm FX DP PPP
C0482659|Coagulation factor XIII inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482659|Coagulation factor XIII inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482659|Fact XIII Inhib PPP-aCnc
C0482659|Coagulation factor XIII inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1114343|Phosphatidylserine Ab.IgA:ACnc:Pt:Ser:Ord
C1114343|PS IgA Ser Ql
C1114343|Phosphatidylserine IgA Ab [Presence] in Serum
C1114343|Phosphatidylserine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Ordinal
C1544431|Beta 2 glycoprotein 1 Ab [Units/volume] in Serum
C1544431|B2 Glycoprot1 Ab Ser-aCnc
C1544431|Beta 2 glycoprotein 1 Ab:ACnc:Pt:Ser:Qn
C1544431|Beta 2 glycoprotein 1 Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative
C1831353|Heparin cofactor II Ag:ACnc:Pt:PPP:Qn
C1831353|Heparin CF II Ag PPP-aCnc
C1831353|Heparin cofactor II Ag [Units/volume] in Platelet poor plasma
C1831353|Heparin cofactor II Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C1623605|Phosphatidylcholine IgA Ab B2GP1 dependent [Multiple of the median] in Serum
C1623605|PC IgA B2GP1 dep MoM Ser
C1623605|Phosphatidylcholine Ab.IgA.B2GP1 dependent:MoM:Pt:Ser:Qn
C1623605|Phosphatidylcholine Antibody.immunoglobulin A.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C2361154|Coagulation surface induced.factor sensitive:Time:Pt:PPP:Qn:Coag
C2361154|Coagulation surface induced.factor sensitive:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2361154|aPTT-FS PPP
C2361154|aPTT.factor sensitive in Platelet poor plasma by Coagulation assay
C0486260|Deprecated reverse INR in Platelet poor plasma by Coagulation assay
C0486260|Coagulation tissue factor induced.normal/Actual:TRto:Pt:Plas:Qn:Coag-inverse ratio
C0486260|Deprecated PT Inv Ratio Plas
C0486260|Coagulation tissue factor induced.normal/Actual:Time Ratio:Point in time:Plasma:Quantitative:Coagulation Assay-inverse ratio
C0482733|Plasm Inhib Ag PPP Imm-mCnc
C0482733|Plasmin inhibitor Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482733|Plasmin inhibitor Ag:MCnc:Pt:PPP:Qn:Imm
C0482733|Plasmin inhibitor Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482744|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex:MCnc:Pt:PPP:Qn:Imm
C0482744|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex [Mass/volume] in Platelet poor plasma by Immunologic method
C0482744|tPA-PAI1 PPP Imm-mCnc
C0482744|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0365485|Plasminogen activator urokinase type [Units/volume] in Urine
C0365485|Plasminogen activator urokinase type:ACnc:Pt:Urine:Qn
C0365485|uPA Ur-aCnc
C0365485|Plasminogen activator urokinase type:Arbitrary Concentration:Point in time:Urine:Quantitative
C2970122|Fibrinogen Antigen:Arbitrary Concentration:Point in time:Tissue, unspecified:Ordinal:Immune Fluorescence
C2970122|Fibrinogen Ag Tiss Ql IF
C2970122|Fibrinogen Ag:ACnc:Pt:Tiss:Ord:IF
C2970122|Fibrinogen Ag [Presence] in Tissue by Immunofluorescence
C0797430|Phosphatidylserine Ab.IgG:ACnc:Pt:Ser:Qn
C0797430|PS IgG Ser-aCnc
C0797430|Phosphatidylserine IgG Ab [Units/volume] in Serum
C0797430|Phosphatidylserine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0551339|Phosphatidylinositol IgA Ab [Units/volume] in Serum
C0551339|PI IgA Ser-aCnc
C0551339|Phosphatidylinositol Ab.IgA:ACnc:Pt:Ser:Qn
C0551339|Phosphatidylinositol Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C0800573|Phosphatidylinositol IgA Ab [Presence] in Serum
C0800573|PI IgA Ser Ql
C0800573|Phosphatidylinositol Ab.IgA:ACnc:Pt:Ser:Ord
C0800573|Phosphatidylinositol Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Ordinal
C0944235|Prekallikrein actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C0944235|Prekallikrein (Fletcher Factor) actual/normal in Platelet poor plasma by Chromogenic method
C0944235|PK Act/Nor PPP Chro
C0944235|Prekallikrein actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1315779|Phosphatidylserine Ab [Presence] in Serum
C1315779|PS Ab Ser Ql
C1315779|Phosphatidylserine Ab:ACnc:Pt:Ser:Ord
C1315779|Phosphatidylserine Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C0365462|Phospholipid Ab [Units/volume] in Serum by Immunoassay
C0365462|Phospholipid Ab:ACnc:Pt:Ser:Qn:EIA
C0365462|Phospholipid Ab Ser EIA-aCnc
C0365462|Phospholipid Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1147245|Phospholipid IgA Ser-aCnc
C1147245|Phospholipid IgA Ab [Units/volume] in Serum
C1147245|Phospholipid Ab.IgA:ACnc:Pt:Ser:Qn
C1147245|Phospholipid Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C1113902|Fibrin+Fibrinogen fragments [Mass/volume] in Serum by Latex agglutination
C1113902|Fibrin+Fibrinogen fragments:MCnc:Pt:Ser:Qn:LA
C1113902|FSP Ser LA-mCnc
C1113902|Fibrin+Fibrinogen fragments:Mass Concentration:Point in time:Serum:Quantitative:Latex Agglutination
C1624143|Phosphatidylcholine Ab.IgG.B2GP1 independent:MoM:Pt:Ser:Qn
C1624143|PC IgG B2GP1 indep MoM Ser
C1624143|Phosphatidylcholine IgG Ab B2GP1 independent [Multiple of the median] in Serum
C1624143|Phosphatidylcholine Antibody.immunoglobulin G.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1644652|von Willebrand factor Antigen actual/Normal:Relative Ratio:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C1644652|Deprecated vWF Ag Act/Nor PPP EIA
C1644652|von Willebrand factor Ag actual/Normal:RelRto:Pt:PPP:Qn:EIA
C1644652|Deprecated von Willebrand factor (vWf) Ag actual/normal in Platelet poor plasma by EIA
C1715215|B2 Glycoprot1 IgG Ser Ql
C1715215|Beta 2 glycoprotein 1 Ab.IgG:ACnc:Pt:Ser:Ord
C1715215|Beta 2 glycoprotein 1 IgG Ab [Presence] in Serum
C1715215|Beta 2 glycoprotein 1 Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C2361160|Coagulation surface induced.lupus sensitive:ACnc:Pt:PPP:Ord:Coag
C2361160|aPTT-LA PPP Ql
C2361160|Coagulation surface induced.lupus sensitive:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C2361160|aPTT.lupus sensitive [Presence] in Platelet poor plasma by Coagulation assay
C1978980|PA Coll 190 ug/mL PRP Ql
C1978980|Platelet aggregation.collagen induced^190 ug/mL:ACnc:Pt:PRP:Ord
C1978980|Platelet aggregation collagen induced [Presence] in Platelet rich plasma --190 ug/mL
C1978980|Platelet aggregation.collagen induced^190 ug/mL:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C1978988|Phosphoserine IgG Ab [Presence] in Serum or Plasma
C1978988|Phosphoserine Ab.IgG:ACnc:Pt:Ser/Plas:Ord
C1978988|Phosphoserine IgG SerPl Ql
C1978988|Phosphoserine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum/Plasma:Ordinal
C1977529|Coagulation factor VII Ag actual/Normal:RelACnc:Pt:PPP:Qn:Imm
C1977529|Coagulation factor VII Ag actual/normal in Platelet poor plasma by Immunologic method
C1977529|Fact VII Ag Act/Nor PPP Imm
C1977529|Coagulation factor VII Antigen actual/Normal:Relative Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482765|Protein S+Acarboxy Ag:ACnc:Pt:PPP:Qn:Imm
C0482765|Protein S+Acarboxy Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482765|Prot S+ACA Ag PPP Imm-aCnc
C0482765|Protein S+Acarboxy Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482685|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --20M post incubation with normal plasma
C0482685|Coagulation tissue factor induced.factor substitution^20M post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C0482685|Coagulation tissue factor induced.factor substitution^20 minutes post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482685|PT 20M NP PPP
C2706782|Thrombin time.factor substitution in Platelet poor plasma by Coagulation assay --immediately after 1:4 addition of normal plasma
C2706782|Coagulation thrombin induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2706782|Coagulation thrombin induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2706782|TT imm 1:4 NP PPP
C2733690|Phosphatidylserine Ab.IgM:MoM:Pt:Ser:Qn
C2733690|Phosphatidylserine IgM Ab [Multiple of the median] in Serum
C2733690|PS IgM MoM Ser
C2733690|Phosphatidylserine Antibody.immunoglobulin M:Multiple of the median:Point in time:Serum:Quantitative
C2598682|PA Rist 800 ug/mL PRP
C2598682|Platelet aggregation ristocetin induced in Platelet rich plasma --800 ug/mL
C2598682|Platelet aggregation.ristocetin induced^800 ug/mL:RelACnc:Pt:PRP:Qn
C2598682|Platelet aggregation.ristocetin induced^800 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0365492|PA ADP PRP
C0365492|Platelet aggregation.adenosine diphosphate induced:RelACnc:Pt:PRP:Qn
C0365492|Platelet aggregation ADP induced in Platelet rich plasma
C0365492|Platelet aggregation.adenosine diphosphate induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C2970620|Coagulation tissue factor induced.INR:RelTime:Pt:PPP^fetus:Qn:Coag
C2970620|INR in Platelet poor plasma from Fetus by Coagulation assay
C2970620|Coagulation tissue factor induced.INR:Relative Time:Point in time:Platelet poor plasma^Fetus:Quantitative:Coagulation Assay
C2970620|INR PPP Fetus
C3481967|Thrombin time.high dose in Platelet poor plasma by Coagulation assay
C3481967|Coagulation thrombin induced.high dose:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3481967|Coagulation thrombin induced.high dose:Time:Pt:PPP:Qn:Coag
C3481967|HiTT PPP
C0798331|Coag Fact Intrinsic PPP-Imp
C0798331|Coagulation factor.intrinsic factor:Imp:Pt:PPP:Nar
C0798331|Coagulation factor.intrinsic factor:Impression/interpretation of study:Point in time:Platelet poor plasma:Narrative
C0798331|Coagulation factor Intrinsic Factor [Interpretation] in Platelet poor plasma Narrative
C0551334|Phosphatidylethanolamine Ab.IgG:ACnc:Pt:Ser:Qn
C0551334|Phosphatidylethanolamine IgG Ab [Units/volume] in Serum
C0551334|PE IgG Ser-aCnc
C0551334|Phosphatidylethanolamine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0796783|PA XXX PRP
C0796783|Platelet aggregation XXX induced in Platelet rich plasma
C0796783|Platelet aggregation.XXX induced:RelACnc:Pt:PRP:Qn
C0796783|Platelet aggregation.XXX induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0800585|Plasminogen activator inhibitor 1 Ag:ACnc:Pt:PPP:Qn:EIA
C0800585|Deprecated Plasminogen activator inhibitor 1 Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0800585|Deprecated PAI1 Ag PPP EIA-aCnc
C0800585|Plasminogen activator inhibitor 1 Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C1315158|LMWH PPP-aCnc
C1315158|LMW Heparin [Units/volume] in Platelet poor plasma
C1315158|Heparin.low molecular weight:ACnc:Pt:PPP:Qn
C1315158|Heparin.low molecular weight:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0482723|Kininogen HMW [Units/volume] in Platelet poor plasma by Coagulation assay
C0482723|Kininogen.high molecular weight:ACnc:Pt:PPP:Qn:Coag
C0482723|HMWK PPP-aCnc
C0482723|Kininogen.high molecular weight:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482729|Lupus anticoagulant neutralization.high phospholipid:Time:Pt:PPP:Qn:Coag
C0482729|Lupus anticoagulant neutralization high phospholipid [Time] in Platelet poor plasma by Coagulation assay
C0482729|Lupus anticoagulant neutralization.high phospholipid:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482729|LA Nt HPL PPP
C0365422|Clot Retraction [Time] in Blood Qualitative by Coagulation assay
C0365422|Clot Retract Bld Ql
C0365422|Coagulum retraction:Time:Pt:Bld:Ord:Coag
C0365422|Coagulum retraction:Time:Point in time:Whole blood:Ordinal:Coagulation Assay
C1315993|Coagulum lysis:Time:Pt:PPP^control:Qn:Coag
C1315993|Coagulum lysis:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1315993|Clot Lysis [Time] in control Platelet poor plasma by Coagulation assay
C1315993|Clot Lysis Cont PPP
C0482604|Antithrombin [Units/volume] in Platelet poor plasma by Chromogenic method
C0482604|Antithrombin:ACnc:Pt:PPP:Qn:Chromo
C0482604|AT III PPP Chro-aCnc
C0482604|Antithrombin:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482627|Coagulation factor VII+Acarboxy Ag activity actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482627|Fact VII+ACA Ag Act/Nor PPP Imm
C0482627|Coagulation factor VII+Acarboxy Ag activity actual/normal in Platelet poor plasma by Immunologic method
C0482627|Coagulation factor VII+Acarboxy Antigen activity actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482645|Coagulation factor X+Acarboxy Ag:ACnc:Pt:PPP:Qn:Imm
C0482645|Fact X+AAC Ag PPP Imm-aCnc
C0482645|Coagulation factor X+Acarboxy Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482645|Coagulation factor X+Acarboxy Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482654|Coagulation factor XII activated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482654|Fact XIIa PPP-aCnc
C0482654|Coagulation factor XII activated activity:ACnc:Pt:PPP:Qn:Coag
C0482654|Coagulation factor XII activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544101|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --12 hours post XXX challenge
C1544101|Coagulation tissue factor induced^12H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544101|Coagulation tissue factor induced^12 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544101|PT 12h p chal PPP
C1715672|B2 Glycoprot1 IgA SerPl EIA-aCnc
C1715672|Beta 2 glycoprotein 1 Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:Enzyme Immunoassay
C1715672|Beta 2 glycoprotein 1 IgA Ab [Units/volume] in Serum or Plasma by Immunoassay
C1715672|Beta 2 glycoprotein 1 Ab.IgA:ACnc:Pt:Ser/Plas:Qn:EIA
C0365516|Deprecated Protein S:Arbitrary Concentration:Point in time:Plasma:Quantitative:COAGULATION ASSAY
C0365516|Protein S:ACnc:Pt:Plas:Qn:Coag
C0365516|Deprecated Prot S Plas-aCnc
C0365516|Deprecated Protein S [Units/volume] in Platelet poor plasma by Coagulation assay
C0365516|Protein S:Arbitrary Concentration:Point in time:Plasma:Quantitative:Coagulation Assay
C1625221|Cardiolipin IgM B2GP1 dep MoM Ser
C1625221|Cardiolipin Ab.IgM.B2GP1 dependent:MoM:Pt:Ser:Qn
C1625221|Cardiolipin IgM Ab B2GP1 dependent [Multiple of the median] in Serum
C1625221|Cardiolipin Antibody.immunoglobulin M.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C2361179|Coagulation surface induced^after addition of protein C activator+factor V depleted plasma/Coagulation surface induced:Time Ratio:Point in time:Platelet poor plasma:Quantitative:COAGULATION ASSAY
C2361179|Coagulation surface induced^after addition of protein C activator+Factor V depleted plasma/Coagulation surface induced:TRto:Pt:PPP:Qn:Coag
C2361179|aPTT protein C activator+FV DP/aPTT PPP
C2361179|aPTT in Platelet poor plasma by Coagulation assay -- after addition of protein C activator + Factor V depleted plasma/aPTT
C2361190|Clotting time.extrinsic coagulation system activated of Blood by Thromboelastography
C2361190|Clotting time.extrinsic coagulation system activated:Time:Pt:Bld:Qn:Thromboelastography
C2361190|Clotting time.extrinsic coagulation system activated:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361190|CT.extrinsic Bld TEG
C2361196|Clotting time.intrinsic coagulation system activated of Blood by Thromboelastography
C2361196|Clotting time.intrinsic coagulation system activated:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361196|Clotting time.intrinsic coagulation system activated:Time:Pt:Bld:Qn:Thromboelastography
C2361196|CT.intrinsic Bld TEG
C1954719|PA AA PRP-aCnc
C1954719|Platelet aggregation.arachidonate induced:ACnc:Pt:PRP:Qn
C1954719|Platelet aggregation arachidonate induced [Units/volume] in Platelet rich plasma
C1954719|Platelet aggregation.arachidonate induced:Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0486259|Deprecated INR in Platelet poor plasma by Coagulation assay
C0486259|Coagulation tissue factor induced.INR:TRto:Pt:Plas:Qn:Coag
C0486259|Deprecated INR Plas
C0486259|Coagulation tissue factor induced.INR:Time Ratio:Point in time:Plasma:Quantitative:Coagulation Assay
C0482674|Deprecated aPTT PPP Qn
C0482674|Deprecated Activated partial thrombplastin time (aPTT).factor substitution in Platelet poor plasma by Coagulation assay --20M post incubation with normal plasma
C0482674|Coagulation surface induced.factor substitution^20M post incubation.37 deg c after addition of normal plasma:Time:Pt:PPP:Qn:Tilt tube
C0482674|Coagulation surface induced.factor substitution^20 minutes post incubation.37 deg c after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Tilt tube
C0482683|Coagulation tissue factor induced.factor substitution^20M post incubation after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C0482683|Coagulation tissue factor induced.factor substitution^20 minutes post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482683|Prothrombin time (PT) factor substitution in control Platelet poor plasma by Coagulation assay --20M post incubation with normal plasma
C0482683|PT 20M NP Cont PPP
C0482684|Deprecated Prothrombin time (PT) factor substitution in Platelet poor plasma from control by Coagulation assay --20M post incubation with normal plasma
C0482684|Deprecated PT PPP Cont Qn
C0482684|Coagulation tissue factor induced.factor substitution^20 minutes post incubation.37 deg c after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Tilt tube
C0482684|Coagulation tissue factor induced.factor substitution^20M post incubation.37 deg c after addition of normal plasma:Time:Pt:PPP^control:Qn:Tilt tube
C2736181|Fact XIII Inhib PPP Ql
C2736181|Coagulation factor XIII inhibitor:ACnc:Pt:PPP:Ord:Coag
C2736181|Coagulation factor XIII inhibitor [Presence] in Platelet poor plasma by Coagulation assay
C2736181|Coagulation factor XIII inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C2736185|Coagulation surface induced.factor substitution^immediately after addition of normal plasma/Coagulation surface induced:TRto:Pt:PPP:Qn:Coag
C2736185|aPTT imm NP/pre NP PPP
C2736185|Coagulation surface induced.factor substitution^immediately after addition of normal plasma/Coagulation surface induced:Time Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2736185|Activated partial thromboplastin time (aPTT).factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma/pre addition of normal plasma
C2733956|Platelet aggregation arachidonate induced in Blood --500 umol/L
C2733956|Platelet aggregation.arachidonate induced^500 umol/L:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733956|Platelet aggregation.arachidonate induced^500 umol/L:RelACnc:Pt:Bld:Qn
C2733956|PA AA 500 umol/L Bld
C2733960|Platelet aggregation collagen induced ATP secretion [Presence] in Blood --5 ug/mL
C2733960|Platelet aggregation.collagen induced ATP secretion^5 ug/mL:ACnc:Pt:Bld:Ord
C2733960|PA Coll ATP secr 5 ug/mL Bld Ql
C2733960|Platelet aggregation.collagen induced ATP secretion^5 ug/mL:Arbitrary Concentration:Point in time:Whole blood:Ordinal
C2598677|PA ADP 50 umol/mL PRP
C2598677|Platelet aggregation.adenosine diphosphate induced^50 umol/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C2598677|Platelet aggregation.adenosine diphosphate induced^50 umol/mL:RelACnc:Pt:PRP:Qn
C2598677|Platelet aggregation ADP induced in Platelet rich plasma --50 umol/mL
C3259773|Circ assist status Patient
C3259773|Circulatory assist status:Prid:Pt:^Patient:Nom
C3259773|Circulatory assist status [Identifier]
C3259773|Circulatory assist status:Presence or Identity:Point in time:^Patient:Nominal
C3259778|Clot strength in Blood by Thromboelastography --after addition of heparinase
C3259778|Clot strength^after addition of heparinase:ArEnrg:Pt:Bld:Qn:Thromboelastography
C3259778|Clot strength^after addition of heparinase:Energy/Area:Point in time:Whole blood:Quantitative:Thromboelastography
C3259778|Clot strength Heparinase Bld TEG
C3259336|Clot lysis estimate Prctl Bld TEG
C3259336|Clot lysis estimate [Percentile] by Thromboelastography
C3259336|Clot lysis estimate:Percentile:Point in time:Whole blood:Quantitative:Thromboelastography
C3259336|Clot lysis estimate:Prctl:Pt:Bld:Qn:Thromboelastography
C0482746|tPA-PAI1 20M PPP Imm-mCnc
C0482746|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex [Mass/volume] in Platelet poor plasma by Immunologic method --20 minutes post venistasis
C0482746|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex^20M post venistasis:MCnc:Pt:PPP:Qn:Imm
C0482746|Plasminogen activator tissue type-Plasminogen activator inhibitor 1 complex^20 minutes post venistasis:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482748|Plasminogen activator tissue type:ACnc:Pt:PPP:Qn:Chromo
C0482748|tPA PPP Chro-aCnc
C0482748|Plasminogen activator tissue type [Units/volume] in Platelet poor plasma by Chromogenic method
C0482748|Plasminogen activator tissue type:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0550594|Deprecated Protein S:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0550594|Protein S:ACnc:Pt:PPP:Qn
C0550594|Deprecated Prot S PPP-aCnc
C0550594|Protein S:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0550594|Deprecated Protein S [Units/volume] in Platelet poor plasma
C0796785|Prekallikrein:ACnc:Pt:PPP:Ord
C0796785|Prekallikrein (Fletcher Factor) [Presence] in Platelet poor plasma
C0796785|PK PPP Ql
C0796785|Prekallikrein:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C0803296|Cardiolipin IgG Titr Ser
C0803296|Cardiolipin Ab.IgG:Titr:Pt:Ser:Qn
C0803296|Cardiolipin IgG Ab [Titer] in Serum
C0803296|Cardiolipin Antibody.immunoglobulin G:Dilution Factor (Titer):Point in time:Serum:Quantitative
C0881721|Platelet function (closure time) collagen+Epinephrine induced [Time] in Blood
C0881721|Platelet function.collagen+Epinephrine induced:Time:Pt:Bld:Qn
C0881721|Platelet function.collagen+Epinephrine induced:Time:Point in time:Whole blood:Quantitative
C0881721|Closure Tme Coll+Epinep Bld
C1369550|Coagulation surface induced.factor substitution^immediately after addition of factor XIII depleted plasma:Time:Pt:PPP:Qn:Coag
C1369550|Coagulation surface induced.factor substitution^immediately after addition of factor XIII depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1369550|aPTT imm FXIII DP PPP
C1369550|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor XIII depleted plasma
C1369552|Coagulation tissue factor induced.factor substitution^immediately after addition of factor II depleted plasma:Time:Pt:PPP:Qn:Coag
C1369552|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor II depleted plasma
C1369552|Coagulation tissue factor induced.factor substitution^immediately after addition of factor II depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1369552|PT imm FII DP PPP
C0482696|Coagulation thrombin induced:Time:Pt:PPP:Qn:Coag
C0482696|Coagulation thrombin induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482696|Thrombin time
C0365464|Phospholipid Ab.IgM:ACnc:Pt:Ser:Qn:EIA
C0365464|Phospholipid IgM Ser EIA-aCnc
C0365464|Phospholipid IgM Ab [Units/volume] in Serum by Immunoassay
C0365464|Phospholipid Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0482772|Prothrombin.activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482772|Prothrom Act/Nor PPP
C0482772|Prothrombin activity actual/normal in Platelet poor plasma by Coagulation assay
C0482772|Prothrombin.activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1315997|PA ADP hi dose PRP Cont
C1315997|Platelet aggregation ADP induced in control Platelet rich plasma --High dose
C1315997|Platelet aggregation.adenosine diphosphate induced^high dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma^Control:Quantitative
C1315997|Platelet aggregation.adenosine diphosphate induced^high dose:RelACnc:Pt:PRP^control:Qn
C1315109|Coagulation factor II inhibitor:ACnc:Pt:PPP:Qn:Coag
C1315109|Coagulation factor II inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C1315109|Fact II Inhib PPP-aCnc
C1315109|Coagulation factor II inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482715|Fibrinopeptide B Ag:MCnc:Pt:PPP:Qn:Imm
C0482715|FpB Ag PPP Imm-mCnc
C0482715|Fibrinopeptide B Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482715|Fibrinopeptide B Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1316056|Phosphatidylinositol Ab:ACnc:Pt:Ser:Qn:EIA
C1316056|PI Ab Ser EIA-aCnc
C1316056|Phosphatidylinositol Ab [Units/volume] in Serum by Immunoassay
C1316056|Phosphatidylinositol Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1114697|Fibrinogen PPP Heat Denat-mCnc
C1114697|Fibrinogen:MCnc:Pt:PPP:Qn:Heat denaturation
C1114697|Fibrinogen [Mass/volume] in Platelet poor plasma by Heat denaturation
C1114697|Fibrinogen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Heat denaturation
C1544110|Coagulation surface induced^4H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544110|Coagulation surface induced^4 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544110|aPTT 4h p chal PPP
C1544110|aPTT in Platelet poor plasma by Coagulation assay --4 hours post XXX challenge
C1544111|Coagulation surface induced^6H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544111|Coagulation surface induced^6 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544111|aPTT 6h p chal PPP
C1544111|aPTT in Platelet poor plasma by Coagulation assay --6 hours post XXX challenge
C1544553|Prothrom IgM SerPl-aCnc
C1544553|Prothrombin IgM Ab [Units/volume] in Serum or Plasma
C1544553|Prothrombin Ab.IgM:ACnc:Pt:Ser/Plas:Qn
C1544553|Prothrombin Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C1644653|von Willebrand factor Ag:ACnc:Pt:PPP:Qn
C1644653|von Willebrand factor (vWf) Ag [Units/volume] in Platelet poor plasma
C1644653|vWF Ag PPP-aCnc
C1644653|von Willebrand factor Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C1978994|Phosphoserine IgM SerPl Ql
C1978994|Phosphoserine Ab.IgM:ACnc:Pt:Ser/Plas:Ord
C1978994|Phosphoserine IgM Ab [Presence] in Serum or Plasma
C1978994|Phosphoserine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum/Plasma:Ordinal
C1953440|D dimer DDU PPP EIA-mCnc
C1953440|Fibrin D-dimer DDU [Mass/volume] in Platelet poor plasma by Immunoassay
C1953440|Fibrin D-dimer DDU:MCnc:Pt:PPP:Qn:EIA
C1953440|Fibrin D-dimer DDU:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C2926242|Protein S Ag/Coagulation factor IX Ag:MRto:Pt:PPP:Qn:Imm
C2926242|Protein S Antigen/Coagulation factor IX Antigen:Mass Ratio:Point in time:Platelet poor plasma:Quantitative:Imm
C2926242|Prot S Ag/Fact IX Ag PPP Imm
C2926242|Protein S Ag/Coagulation factor IX Ag [Mass Ratio] in Platelet poor plasma by Immunologic method
C0365475|Plasminogen activator inhibitor 1:MCnc:Pt:PPP:Qn:Chromo
C0365475|Plasminogen activator inhibitor 1 [Mass/volume] in Platelet poor plasma by Chromogenic method
C0365475|PAI1 PPP Chro-mCnc
C0365475|Plasminogen activator inhibitor 1:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C2713204|Deprecated Cardiolipin IgM Ab [Units/volume] in Serum by Immunoassay
C2713204|Cardiolipin Ab.IgM:ACnc:Pt:Ser:Qn:EIA
C2713204|Deprecated Cardiolipin IgM Ser EIA-aCnc
C2713204|Cardiolipin Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C2713204|Deprecated Cardiolipin IgM Ab [Units/volume] in Serum by Immunoassay.
C3260553|Coagulation surface induced.factor substitution^after addition of normal plasma 2 hours post incubation separate tubes:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3260553|Coagulation surface induced.factor substitution^after addition of normal plasma 2H post incubation separate tubes:Time:Pt:PPP:Qn:Coag
C3260553|aPTT NP 2h separate PPP
C3260553|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --with normal plasma 2H post incubation separate tubes
C0482743|Plasminogen activator inhibitor Ag:MCnc:Pt:PPP:Qn:Imm
C0482743|Plasminogen activator inhibitor Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482743|PAI Ag PPP Imm-mCnc
C0482743|Plasminogen activator inhibitor Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482747|Plasminogen activator urokinase type:ACnc:Pt:PPP:Qn
C0482747|uPA PPP-aCnc
C0482747|Plasminogen activator urokinase type [Units/volume] in Platelet poor plasma
C0482747|Plasminogen activator urokinase type:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0482760|Protein C:ACnc:Pt:PPP:Qn:Chromo
C0482760|Protein C [Units/volume] in Platelet poor plasma by Chromogenic method
C0482760|Prot C PPP Chro-aCnc
C0482760|Protein C:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3481609|Argatroban:ACnc:Pt:PPP:Qn:Chromo
C3481609|Argatroban:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3481609|Argatroban [Units/volume] in Platelet poor plasma by Chromogenic method
C3481609|Argatroban PPP Chro-aCnc
C0799997|FpA Ag Prt Imm-aCnc
C0799997|Fibrinopeptide A Ag:ACnc:Pt:Periton fld:Qn:Imm
C0799997|Fibrinopeptide A Ag [Units/volume] in Peritoneal fluid by Immunologic method
C0799997|Fibrinopeptide A Antigen:Arbitrary Concentration:Point in time:Peritoneal fluid /ascites:Quantitative:Imm
C2713202|Deprecated von Willebrand factor (vWf) Ag [Units/volume] in Platelet poor plasma by Immunologic method
C2713202|Deprecated vWF:Ag PPP Imm-aCnc
C2713202|von Willebrand factor Ag:ACnc:Pt:PPP:Qn:Imm
C2713202|von Willebrand factor Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0796780|Activated protein C resistance:ACnc:Pt:Bld:Ord:Probe.amp.tar
C0796780|aPCR Bld Ql PCR
C0796780|Activated protein C resistance:Arbitrary Concentration:Point in time:Whole blood:Ordinal:DNA Nucleic Acid Probe.amp.tar
C0796780|Activated protein C resistance [Presence] in Blood by Probe and target amplification method
C0551343|Phosphatidylserine IgG Ab [Presence] in Serum
C0551343|Phosphatidylserine Ab.IgG:ACnc:Pt:Ser:Ord
C0551343|PS IgG Ser Ql
C0551343|Phosphatidylserine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C0364003|Antithrombin Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0364003|AT III Ag PPP Imm-mCnc
C0364003|Antithrombin Ag:MCnc:Pt:PPP:Qn:Imm
C0364003|Antithrombin Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0943508|Prothrombin Ag actual/normal in Platelet poor plasma by Immunologic method
C0943508|Prothrom Ag Act/Nor PPP Imm
C0943508|Prothrombin Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0943508|Prothrombin Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0943511|von Willebrand factor Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0943511|vWF Ag Act/Nor PPP Imm
C0943511|von Willebrand factor (vWf) Ag actual/normal in Platelet poor plasma by Immunologic method
C0943511|von Willebrand factor Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1316138|PA Rist + Cont PRP PPP
C1316138|Platelet aggregation.ristocetin+Control PRP induced in Platelet poor plasma
C1316138|Platelet aggregation.ristocetin+Control PRP induced:RelACnc:Pt:PPP:Qn
C1316138|Platelet aggregation.ristocetin+Control PRP induced:Relative Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C1369554|Coagulation surface induced.factor substitution^immediately after addition of factor XII depleted plasma:Time:Pt:PPP:Qn:Coag
C1369554|Coagulation surface induced.factor substitution^immediately after addition of factor XII depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1369554|aPTT imm FXII DP PPP
C1369554|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor XII depleted plasma
C0482710|Fibrinopeptide B beta (1-14) Ag:MCnc:Pt:PPP:Qn:Imm
C0482710|Fibrinopeptide B beta (1-14) Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482710|FpB Beta1-14 Ag PPP Imm-mCnc
C0482710|Fibrinopeptide B beta (1-14) Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1316022|PA Rist 600 ug/mL PRP
C1316022|Platelet aggregation ristocetin induced in Platelet rich plasma --600 ug/mL
C1316022|Platelet aggregation.ristocetin induced^600 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1316022|Platelet aggregation.ristocetin induced^600 ug/mL:RelACnc:Pt:PRP:Qn
C0482609|Coagulation factor IX inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482609|Coagulation factor IX inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482609|Fact IX Inhib PPP-aCnc
C0482609|Coagulation factor IX inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482617|Coagulation factor V activity actual/normal in Platelet poor plasma by Coagulation assay
C0482617|Fact V Act/Nor PPP
C0482617|Coagulation factor V activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482617|Coagulation factor V activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482630|Coagulation factor VIII inhibitor:ACnc:Pt:PPP:Ord:Coag
C0482630|Coagulation factor VIII inhibitor [Presence] in Platelet poor plasma by Coagulation assay
C0482630|Fact VIII Inhib PPP Ql
C0482630|Coagulation factor VIII inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C1147901|von Willebrand factor (vWf) multimers [Presence] in Platelet poor plasma
C1147901|von Willebrand factor multimers:ACnc:Pt:PPP:Ord
C1147901|vWF multimers PPP Ql
C1147901|von Willebrand factor multimers:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C1113984|Coagulation factor IX inhibitor [Presence] in Platelet poor plasma by Coagulation assay
C1113984|Fact IX Inhib PPP Ql
C1113984|Coagulation factor IX inhibitor:ACnc:Pt:PPP:Ord:Coag
C1113984|Coagulation factor IX inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C1544099|Coagulation tissue factor induced^6H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544099|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --6 hours post XXX challenge
C1544099|Coagulation tissue factor induced^6 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544099|PT 6h p chal PPP
C1830125|Coagulation thrombin induced^after addition of heparinase:Time:Pt:PPP:Qn:Coag
C1830125|Thrombin time in Platelet poor plasma by Coagulation assay --after addition of heparinase
C1830125|Coagulation thrombin induced^after addition of heparinase:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1830125|TT Heparinase PPP
C1623607|PE IgG B2GP1 dep MoM Ser
C1623607|Phosphatidylethanolamine Ab.IgG.B2GP1 dependent:MoM:Pt:Ser:Qn
C1623607|Phosphatidylethanolamine IgG Ab B2GP1 dependent [Multiple of the median] in Serum
C1623607|Phosphatidylethanolamine Antibody.immunoglobulin G.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C1646206|Phosphatidylserine IgA Ab B2GP1 dependent [Multiple of the median] in Serum
C1646206|PS IgA B2GP1 dep MoM Ser
C1646206|Phosphatidylserine Ab.IgA.B2GP1 dependent:MoM:Pt:Ser:Qn
C1646206|Phosphatidylserine Antibody.immunoglobulin A.B2GP1 dependent:Multiple of the median:Point in time:Serum:Quantitative
C1643196|Prothrombin time (PT) in Platelet poor plasma by Coagulation 1:1 saline
C1643196|Coagulation tissue factor induced:Time:Pt:PPP:Qn:Coag.saline 1:1
C1643196|Coagulation tissue factor induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay.saline 1:1
C1643196|PT PPP 1:1 saline
C2361170|Prothrombin time (PT) PIVKA sensitive actual/normal in Platelet poor plasma by Coagulation assay
C2361170|PT PIVKA sensitive Act/Nor PPP
C2361170|Coagulation tissue factor induced.PIVKA sensitive actual/Normal:RelTime:Pt:PPP:Qn:Coag
C2361170|Coagulation tissue factor induced.PIVKA sensitive actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2361206|MCF.intrinsic Bld TEG
C2361206|Maximum clot firmness.intrinsic coagulation system activated [Length] in Blood by Thromboelastography
C2361206|Maximum clot firmness.intrinsic coagulation system activated:Length:Point in time:Whole blood:Quantitative:Thromboelastography
C2361206|Maximum clot firmness.intrinsic coagulation system activated:Len:Pt:Bld:Qn:Thromboelastography
C0482734|Plasmin-plasmin inhibitor complex:MCnc:Pt:PPP:Qn:Imm
C0482734|PAP PPP Imm-mCnc
C0482734|Plasmin-plasmin inhibitor complex [Mass/volume] in Platelet poor plasma by Immunologic method
C0482734|Plasmin-plasmin inhibitor complex:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C2924050|Coagulation dilute Russell viper venom induced.factor substitution^1H post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2924050|Coagulation dilute Russell viper venom induced.factor substitution^1 hour post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2924050|dRVVT 1h NP PPP
C2924050|dRVVT factor substitution in Platelet poor plasma by Coagulation assay --1H post incubation with normal plasma
C2598678|PA ADP 100 umol/mL PRP
C2598678|Platelet aggregation ADP induced in Platelet rich plasma --100 umol/mL
C2598678|Platelet aggregation.adenosine diphosphate induced^100 umol/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C2598678|Platelet aggregation.adenosine diphosphate induced^100 umol/mL:RelACnc:Pt:PRP:Qn
C0484865|Coagulation reptilase induced:Time:Pt:PPP:Qn:Coag
C0484865|Coagulation reptilase induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0484865|Reptilase time
C0484868|Fibrinogen Ag [Presence] in Tissue by Immune stain
C0484868|Fibrinogen Ag:ACnc:Pt:Tiss:Ord:Immune stain
C0484868|Fibrinogen Ag Tiss Ql ImStn
C0484868|Fibrinogen Antigen:Arbitrary Concentration:Point in time:Tissue, unspecified:Ordinal:Immune stain
C2603365|Deprecated Activated partial thrombplastin time (aPTT) in Blood from control by Coagulation assay
C2603365|Coagulation surface induced:Time:Pt:Bld^control:Qn:Coag
C2603365|Deprecated aPTT Bld Cont Qn
C2603365|Coagulation surface induced:Time:Point in time:Whole blood^Control:Quantitative:Coagulation Assay
C0551342|PS IgA Ser-aCnc
C0551342|Phosphatidylserine IgA Ab [Units/volume] in Serum
C0551342|Phosphatidylserine Ab.IgA:ACnc:Pt:Ser:Qn
C0551342|Phosphatidylserine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C0880259|Plasminogen activator inhibitor 1 Ag:MCnc:Pt:PPP:Qn:Imm
C0880259|Plasminogen activator inhibitor 1 Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0880259|PAI1 Ag PPP Imm-mCnc
C0880259|Plasminogen activator inhibitor 1 Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0803244|Phospholipid IgM Ser Ql
C0803244|Phospholipid IgM Ab [Presence] in Serum
C0803244|Phospholipid Ab.IgM:ACnc:Pt:Ser:Ord
C0803244|Phospholipid Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482730|Lupus anticoagulant neutralization platelet [Time] in Platelet poor plasma by Coagulation assay
C0482730|Lupus anticoagulant neutralization.platelet:Time:Pt:PPP:Qn:Coag
C0482730|Lupus anticoagulant neutralization.platelet:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482730|LA Nt Platelet PPP
C0365429|Fibrin+Fibrinogen fragments [Units/volume] in Serum by Latex agglutination
C0365429|Fibrin+Fibrinogen fragments:ACnc:Pt:Ser:Qn:LA
C0365429|FSP Ser LA-aCnc
C0365429|Fibrin+Fibrinogen fragments:Arbitrary Concentration:Point in time:Serum:Quantitative:Latex Agglutination
C0482641|Coagulation factor X activity actual/normal in Platelet poor plasma by Coagulation assay
C0482641|Coagulation factor X activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C0482641|Fact X Act/Nor PPP
C0482641|Coagulation factor X activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482643|Fact X Ag PPP Imm-aCnc
C0482643|Coagulation factor X Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482643|Coagulation factor X Ag:ACnc:Pt:PPP:Qn:Imm
C0482643|Coagulation factor X Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1544103|Coagulation surface induced^2H pre XXX challenge:Time:Pt:PPP:Qn:Coag
C1544103|Coagulation surface induced^2 hours pre XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544103|aPTT 2h pre chal PPP
C1544103|aPTT in Platelet poor plasma by Coagulation assay --2 hours pre XXX challenge
C1542937|Coagulation surface induced^18H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1542937|Coagulation surface induced^18H post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1542937|aPTT 18h p chal PPP
C1542937|aPTT in Platelet poor plasma by Coagulation assay --18 hours post XXX challenge
C1624713|PS IgM B2GP1 indep MoM Ser
C1624713|Phosphatidylserine Ab.IgM.B2GP1 independent:MoM:Pt:Ser:Qn
C1624713|Phosphatidylserine IgM Ab B2GP1 independent [Multiple of the median] in Serum
C1624713|Phosphatidylserine Antibody.immunoglobulin M.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C2360889|Coagulation dilute Russell viper venom induced.factor substitution^immediately after 4:1 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2360889|Coagulation dilute Russell viper venom induced.factor substitution^immediately after 4:1 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2360889|dRVVT factor substitution in Platelet poor plasma by Coagulation assay --immediately after 4:1 addition of normal plasma
C2360889|dRVVT imm 4:1 NP PPP
C1954161|Coagulation surface induced^after addition of APC:Time:Pt:PPP:Qn:Coag
C1954161|Coagulation surface induced^after addition of APC:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1954161|aPTT after addition of APC PPP
C1954161|aPTT in Platelet poor plasma by Coagulation assay --after addition of APC
C1953449|Fibrin D-dimer FEU [Mass/volume] in Platelet poor plasma
C1953449|Fibrin D-dimer FEU:MCnc:Pt:PPP:Qn
C1953449|D dimer FEU PPP-mCnc
C1953449|Fibrin D-dimer FEU:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C2735810|Platelet Ab:ACnc:Pt:Ser:Ord:IF
C2735810|Platelet Ab [Presence] in Serum by Immunofluorescence
C2735810|Platelet Ab Ser Ql IF
C2735810|Platelet Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal:Immune Fluorescence
C2598681|PA AA 500 ug/mL PRP
C2598681|Platelet aggregation.arachidonate induced^500 ug/mL:RelACnc:Pt:PRP:Qn
C2598681|Platelet aggregation arachidonate induced in Platelet rich plasma --500 ug/mL
C2598681|Platelet aggregation.arachidonate induced^500 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0482775|von Willebrand factor.ristocetin cofactor activity actual/Normal:RelTime:Pt:PPP:Qn:Aggr
C0482775|von Willebrand factor (vWf) ristocetin cofactor actual/normal in Platelet poor plasma by Aggregation
C0482775|vWf:RCo Act/Nor PPP Aggr
C0482775|von Willebrand factor.ristocetin cofactor activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Aggr
C0484870|Phospholipid IgG Ser-aCnc
C0484870|Phospholipid IgG Ab [Units/volume] in Serum
C0484870|Phospholipid Ab.IgG:ACnc:Pt:Ser:Qn
C0484870|Phospholipid Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative
C0483194|Coagulation thrombin induced
C0483194|Coagulation reptilase induced
C0550585|Bleeding time:Time:Point in time:^Patient:Quantitative
C0550585|Bleeding time
C0550585|Bleeding time:Time:Pt:^Patient:Qn
C0550585|Bleeding time Patient
C0947259|Plasm Inhib Act/Nor PPP Chro
C0947259|Plasmin inhibitor actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C0947259|Plasmin inhibitor actual/normal in Platelet poor plasma by Chromogenic method
C0947259|Plasmin inhibitor actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0881642|vWF multimers PPP EIA-aCnc
C0881642|von Willebrand factor multimers:ACnc:Pt:PPP:Qn:EIA
C0881642|von Willebrand factor (vWf) multimers in Platelet poor plasma by Immunoassay
C0881642|von Willebrand factor multimers:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C1317030|Coagulation dilute Russell viper venom induced.factor substitution^immediately after 1:2 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1317030|Coagulation dilute Russell viper venom induced.factor substitution^immediately after 1:2 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1317030|dRVVT factor substitution in Platelet poor plasma by Coagulation assay --immediately after 1:2 addition of normal plasma
C1317030|dRVVT imm 1:2 NP PPP
C0482707|Fibrinogen:MCnc:Pt:PPP:Ord:Turbidimetry
C0482707|Deprecated Fibrinogen
C0482707|Deprecated Fibrinogen PPP Ql
C0482707|Fibrinogen:Mass Concentration:Point in time:Platelet poor plasma:Ordinal:Turbidimetry
C1315989|PA Coll hi dose PRP
C1315989|Platelet aggregation.collagen induced^high dose:RelACnc:Pt:PRP:Qn
C1315989|Platelet aggregation.collagen induced^high dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1315989|Platelet aggregation collagen induced in Platelet rich plasma --High dose
C0365322|Bleeding time:Time:Point in time:^Patient:Quantitative:Duke
C0365322|Bleeding time by Duke method
C0365322|Bleeding time:Time:Pt:^Patient:Qn:Duke
C0365322|Bleeding time Patient Duke
C0482615|Fact V Inhib PPP-aCnc
C0482615|Coagulation factor V inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482615|Coagulation factor V inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482615|Coagulation factor V inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482635|Coagulation factor VIII activity actual/Normal:RelTime:Pt:PPP:Qn:Coag.two stage
C0482635|Coagulation factor VIII activity actual/normal in Platelet poor plasma by Coagulation.2 stage
C0482635|Fact VIII Act/Nor PPP 2Stg
C0482635|Coagulation factor VIII activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay.two stage
C0482640|Coagulation factor X activated activity:ACnc:Pt:PPP:Qn:Coag
C0482640|Coagulation factor X activated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482640|Fact Xa PPP-aCnc
C0482640|Coagulation factor X activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482646|Fact X+AAC Ag Act/Nor PPP Imm
C0482646|Coagulation factor X+Acarboxy Ag actual/normal in Platelet poor plasma by Immunologic method
C0482646|Coagulation factor X+Acarboxy Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482646|Coagulation factor X+Acarboxy Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482647|Fact XI Inhib PPP-aCnc
C0482647|Coagulation factor XI inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482647|Coagulation factor XI inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482647|Coagulation factor XI inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1715082|Coagulation surface induced:Time:Pt:PPP:Qn:Coag.saline 1:1
C1715082|Coagulation surface induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay.saline 1:1
C1715082|aPTT PPP 1:1 saline
C1715082|aPTT in Platelet poor plasma by Coagulation 1:1 saline
C2361153|Activated protein C resistance [Presence] in Platelet poor plasma by Coagulation assay
C2361153|aPCR PPP Ql
C2361153|Activated protein C resistance:Threshold:Pt:PPP:Ord:Coag
C2361153|Activated protein C resistance:Threshold:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C2361157|Prothrombin time (PT) PIVKA insensitive actual/normal in Platelet poor plasma by Coagulation assay
C2361157|PT PIVKA insensitive Act/Nor PPP
C2361157|Coagulation tissue factor induced.PIVKA insensitive actual/Normal:RelTime:Pt:PPP:Qn:Coag
C2361157|Coagulation tissue factor induced.PIVKA insensitive actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2361204|MCF.platelet inhib Bld TEG
C2361204|Maximum clot firmness.extrinsic coagulation system activated.platelets inhibited:Len:Pt:Bld:Qn:Thromboelastography
C2361204|Maximum clot firmness.extrinsic coagulation system activated.platelets inhibited [Length] in Blood by Thromboelastography
C2361204|Maximum clot firmness.extrinsic coagulation system activated.platelets inhibited:Length:Point in time:Whole blood:Quantitative:Thromboelastography
C1954163|Fibrin+Fibrinogen fragments [Titer] in Platelet poor plasma by Latex agglutination
C1954163|FSP Titr PPP LA
C1954163|Fibrin+Fibrinogen fragments:Titr:Pt:PPP:Qn:LA
C1954163|Fibrin+Fibrinogen fragments:Dilution Factor (Titer):Point in time:Platelet poor plasma:Quantitative:Latex Agglutination
C2926240|Protein C Ag/Coagulation factor IX Ag:MRto:Pt:PPP:Qn:Imm
C2926240|Protein C Ag/Coagulation factor IX Ag [Mass Ratio] in Platelet poor plasma by Immunologic method
C2926240|Prot C Ag/Fact IX Ag PPP Imm
C2926240|Protein C Antigen/Coagulation factor IX Antigen:Mass Ratio:Point in time:Platelet poor plasma:Quantitative:Imm
C2735574|Lupus anticoagulant neutralization dilute phospholipid/Lupus anticoagulant neutralization.high phospholipid [Ratio] in Platelet poor plasma by Coagulation assay
C2735574|Lupus anticoagulant neutralization.dilute phospholipid/Lupus anticoagulant neutralization.high phospholipid:Ratio:Pt:PPP:Qn:Coag
C2735574|Lupus anticoagulant neutralization.dilute phospholipid/Lupus anticoagulant neutralization.high phospholipid:Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2735574|LA Nt dPL/LA Nt HPL PPP-Rto
C3259780|Coagulation index:ACnc:Pt:Bld:Qn:Thromboelastography
C3259780|CI Bld TEG-aCnc
C3259780|Coagulation index:Arbitrary Concentration:Point in time:Whole blood:Quantitative:Thromboelastography
C3259780|Coagulation index in Blood by Thromboelastography
C0482754|PF3 PPP-aCnc
C0482754|Platelet factor 3:ACnc:Pt:PPP:Qn
C0482754|Platelet factor 3 [Units/volume] in Platelet poor plasma
C0482754|Platelet factor 3:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0482773|von Willebrand factor Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482773|vWF Ag PPP Imm-aCnc
C0482773|von Willebrand factor Ag:ACnc:Pt:PPP:Qn:Imm
C0482773|von Willebrand factor (vWf) Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0485837|Cardiolipin IgA SerPl-aCnc
C0485837|Cardiolipin IgA Ab [Units/volume] in Serum or Plasma
C0485837|Cardiolipin Ab.IgA:ACnc:Pt:Ser/Plas:Qn
C0485837|Cardiolipin Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C3481608|Dabigatran:ACnc:Pt:PPP:Qn:Chromo
C3481608|Dabigatran:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3481608|Dabigatran PPP Chro-aCnc
C3481608|Dabigatran [Units/volume] in Platelet poor plasma by Chromogenic method
C0033706|Factor, Differentiation Reversal
C0033706|Prothrombin
C0033706|Blood-coagulation factor II
C0033706|Factor II, Coagulation
C0033706|II, Coagulation Factor
C0033706|COAG FACTOR II
C0033706|BLOOD COAG FACTOR II
C0033706|Coagulation Factor II
C0033706|EC 3.4.21.5
C0033706|Factor II
C0033706|Blood Coagulation Factor II
C0033706|Prothrombin [Chemical/Ingredient]
C0033706|Differentiation Reversal Factor
C0033706|Coagulation factor II (substance)
C0550590|Coagulation surface induced^4th specimen:Time:Pt:PPP:Qn:Coag
C0550590|Coagulation surface induced^4th specimen:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0550590|aPTT sp4 PPP
C0550590|aPTT in Platelet poor plasma by Coagulation assay --4th specimen
C0551344|Phosphatidylserine IgM Ab [Presence] in Serum
C0551344|PS IgM Ser Ql
C0551344|Phosphatidylserine Ab.IgM:ACnc:Pt:Ser:Ord
C0551344|Phosphatidylserine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482721|Heparin.unfractionated:ACnc:Pt:PPP:Qn:Coag
C0482721|Heparin unfractionated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482721|Heparin.unfractionated:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482721|UFH PPP clot-aCnc
C0482660|Coagulation factor XIII activated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482660|Fact XIIIa PPP-aCnc
C0482660|Coagulation factor XIII activated activity:ACnc:Pt:PPP:Qn:Coag
C0482660|Coagulation factor XIII activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482727|Lupus anticoagulant:Imp:Pt:PPP:Nom
C0482727|Lupus anticoagulant:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal
C0482727|LA PPP-Imp
C0482727|Lupus anticoagulant [Interpretation] in Platelet poor plasma
C1315999|PA Epineph PRP Cont
C1315999|Platelet aggregation epinephrine induced in control Platelet rich plasma
C1315999|Platelet aggregation.epinephrine induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma^Control:Quantitative
C1315999|Platelet aggregation.epinephrine induced:RelACnc:Pt:PRP^control:Qn
C1316002|PA Rist lo dose PRP Cont
C1316002|Platelet aggregation ristocetin induced in control Platelet rich plasma --Low dose
C1316002|Platelet aggregation.ristocetin induced^low dose:RelACnc:Pt:PRP^control:Qn
C1316002|Platelet aggregation.ristocetin induced^low dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma^Control:Quantitative
C1146787|Protein S actual/normal in Platelet poor plasma by Chromogenic method
C1146787|Protein S actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C1146787|Prot S Act/Nor PPP Chro
C1146787|Protein S actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482612|Coagulation factor IX activity:ACnc:Pt:PPP:Qn:Chromo
C0482612|Fact IX PPP Chro-aCnc
C0482612|Coagulation factor IX activity [Units/volume] in Platelet poor plasma by Chromogenic method
C0482612|Coagulation factor IX activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C0482619|Coagulation factor V Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0482619|Fact V Ag Act/Nor PPP Imm
C0482619|Coagulation factor V Ag actual/normal in Platelet poor plasma by Immunologic method
C0482619|Coagulation factor V Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482620|Fact VII Inhib PPP-aCnc
C0482620|Coagulation factor VII inhibitor:ACnc:Pt:PPP:Qn:Coag
C0482620|Coagulation factor VII inhibitor [Units/volume] in Platelet poor plasma by Coagulation assay
C0482620|Coagulation factor VII inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544104|Coagulation surface induced^baseline:Time:Pt:PPP:Qn:Coag
C1544104|Coagulation surface induced^baseline:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544104|aPTT BS PPP
C1544104|aPTT in Platelet poor plasma by Coagulation assay --baseline
C1544433|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --immediately after addition of factor VIII depleted plasma
C1544433|Coagulation tissue factor induced.factor substitution^immediately after addition of factor VIII depleted plasma:Time:Pt:PPP:Qn:Coag
C1544433|Coagulation tissue factor induced.factor substitution^immediately after addition of factor VIII depleted plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544433|PT imm FVIII DP PPP
C1507507|PA XXX PRP Donr
C1507507|Platelet aggregation XXX induced in Platelet rich plasma from donor
C1507507|Platelet aggregation.XXX induced:RelACnc:Pt:PRP^donor:Qn
C1507507|Platelet aggregation.XXX induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma^Donor:Quantitative
C1830307|INR BldC
C1830307|INR in Capillary blood by Coagulation assay
C1830307|Coagulation tissue factor induced.INR:RelTime:Pt:BldC:Qn:Coag
C1830307|Coagulation tissue factor induced.INR:Relative Time:Point in time:Blood capillary:Quantitative:Coagulation Assay
C2361158|Kininogen HMW activity actual/normal in Platelet poor plasma by Coagulation assay
C2361158|HMWK activity Act/Nor PPP
C2361158|Kininogen.high molecular weight activity actual/Normal:RelTime:Pt:PPP:Qn:Coag
C2361158|Kininogen.high molecular weight activity actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2361188|Clot formation.intrinsic coagulation system activated.heparin insensitive [Time] in Blood by Thromboelastography
C2361188|Clot formation.intrinsic coagulation system activated.heparin insensitive:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361188|Clot formation.intrinsic coagulation system activated.heparin insensitive:Time:Pt:Bld:Qn:Thromboelastography
C2361188|CFT.heparin insens Bld TEG
C1978254|aPTT circulating inhib PPP Ql
C1978254|Coagulation surface induced circulating inhibitor:ACnc:Pt:PPP:Ord
C1978254|Coagulation surface induced circulating inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C1978254|aPTT circulating inhibitor [Presence] in Platelet poor plasma
C1978283|Coagulation dilute Russell viper venom induced/Coagulation dilute Russell viper venom induced.excess phospholipid:Ratio:Pt:PPP:Qn:Coag
C1978283|Coagulation dilute Russell viper venom induced/Coagulation dilute Russell viper venom induced.excess phospholipid:Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1978283|dRVVT screen to confirm ratio
C1978283|dRVVT/dRVVT W excess phospholipid (screen to confirm ratio)
C1978992|Phosphoethanolamine Ab.IgG:ACnc:Pt:Ser/Plas:Ord
C1978992|PETN IgG SerPl Ql
C1978992|Phosphoethanolamine IgG Ab [Presence] in Serum or Plasma
C1978992|Phosphoethanolamine Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum/Plasma:Ordinal
C1976975|Coagulation surface induced.factor substitution^2H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1976975|Coagulation surface induced.factor substitution^2 hours post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1976975|aPTT 2h p 1:4 NP PPP
C1976975|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --2H post incubation with 1:4 normal plasma
C1976977|Coagulation surface induced.factor substitution^after addition of normal plasma 1H post incubation separate tubes:Time:Pt:PPP:Qn:Coag
C1976977|Coagulation surface induced.factor substitution^after addition of normal plasma 1 hour post incubation separate tubes:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1976977|aPTT NP 1h separate PPP
C1976977|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --with normal plasma 1H post incubation separate tubes
C2733680|Lupus anticoagulant neutralization high phospholipid.factor substitution [Time] in Platelet poor plasma by Coagulation assay --immediately after 1:2 addition of platelet lysate
C2733680|Lupus anticoagulant neutralization.high phospholipid.factor substitution^immediately after 1:2 addition of platelet lysate:Time:Pt:PPP:Qn:Coag
C2733680|Lupus anticoagulant neutralization.high phospholipid.factor substitution^immediately after 1:2 addition of platelet lysate:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2733680|LA Nt HPL imm 1:2 Plat lysate PPP
C2733957|PA Coll 1 ug/mL Bld
C2733957|Platelet aggregation collagen induced in Blood --1 ug/mL
C2733957|Platelet aggregation.collagen induced^1 ug/mL:RelACnc:Pt:Bld:Qn
C2733957|Platelet aggregation.collagen induced^1 ug/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733738|Platelet aggregation.arachidonate induced ATP secretion^500 umol/L:Presence:Point in time:Whole blood:Ordinal
C2733738|Platelet aggregation arachidonate induced ATP secretion [Presence] in Blood --500 umol/L
C2733738|Platelet aggregation.arachidonate induced ATP secretion^500 umol/L:Pr:Pt:Bld:Ord
C2733738|PA AA ATP secr 500 umol/L Bld Ql
C2733959|Platelet aggregation.collagen induced ATP secretion^1 ug/mL:ACnc:Pt:Bld:Ord
C2733959|Platelet aggregation collagen induced ATP secretion [Presence] in Blood --1 ug/mL
C2733959|PA Coll ATP secr 1 ug/mL Bld Ql
C2733959|Platelet aggregation.collagen induced ATP secretion^1 ug/mL:Arbitrary Concentration:Point in time:Whole blood:Ordinal
C3259752|Normalized silica clotting time:Ratio:Pt:PPP:Qn
C3259752|Normalized silica clotting time of Platelet poor plasma
C3259752|Normalized silica clotting time:Ratio:Point in time:Platelet poor plasma:Quantitative
C3259752|Normalized SCT PPP-Rto
C3259779|Heparin Nt Bld Ql TEG
C3259779|Heparin neutralization:ACnc:Pt:Bld:Ord:Thromboelastography
C3259779|Heparin neutralization [Presence] in Blood by Thromboelastography
C3259779|Heparin neutralization:Arbitrary Concentration:Point in time:Whole blood:Ordinal:Thromboelastography
C0482692|Coagulation tissue factor induced.normal/Actual:RelTime:Pt:PPP:Qn:Coag inverse ratio
C0482692|Coagulation tissue factor induced.normal/Actual:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay inverse ratio
C0482692|Prothrombin index in Platelet poor plasma by Coagulation assay
C0482692|PT index PPP
C0365495|PA Coll PRP
C0365495|Platelet aggregation.collagen induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0365495|Platelet aggregation collagen induced in Platelet rich plasma
C0365495|Platelet aggregation.collagen induced:RelACnc:Pt:PRP:Qn
C0482758|Prekallikrein (Fletcher Factor) [Mass/volume] in Platelet poor plasma by Chromogenic method
C0482758|PK PPP Chro-mCnc
C0482758|Prekallikrein:MCnc:Pt:PPP:Qn:Chromo
C0482758|Prekallikrein:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3481501|Coagulation kaolin induced actual/Normal:RelTime:Pt:PPP:Qn
C3481501|Kaolin activated time actual/normal in Platelet poor plasma
C3481501|Coagulation kaolin induced actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative
C3481501|KCT Act/Nor PPP
C0368981|Coagulation calcium ion induced
C0032139|Inhibitor, Plasmin
C0032139|PLASMIN INHIB
C0032139|plasmin inhibitor
C0032139|Inhibitors, Plasmin
C0032139|Antiplasmins
C0032139|Plasmin Inhibitors
C0032139|Plasmin inhibitor (substance)
C0032139|Plasmin inhibitor, NOS
C0485827|Phosphatidylserine Ab.IgM:ACnc:Pt:Ser:Ord:EIA
C0485827|Phosphatidylserine IgM Ab [Presence] in Serum by Immunoassay
C0485827|PS IgM Ser Ql EIA
C0485827|Phosphatidylserine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Ordinal:Enzyme Immunoassay
C0797431|Phosphatidylserine IgM Ab [Units/volume] in Serum
C0797431|Phosphatidylserine Ab.IgM:ACnc:Pt:Ser:Qn
C0797431|PS IgM Ser-aCnc
C0797431|Phosphatidylserine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0797197|PC IgM Ser EIA-aCnc
C0797197|Phosphatidylcholine IgM Ab [Units/volume] in Serum by Immunoassay
C0797197|Phosphatidylcholine Ab.IgM:ACnc:Pt:Ser:Qn:EIA
C0797197|Phosphatidylcholine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0803239|Cardiolipin Ab.IgG:Imp:Pt:Ser:Nom
C0803239|Cardiolipin IgG Ser-Imp
C0803239|Cardiolipin Antibody.immunoglobulin G:Impression/interpretation of study:Point in time:Serum:Nominal
C0803239|Cardiolipin IgG Ab [Interpretation] in Serum
C0800571|Phosphatidylglycerol Ab.IgG:ACnc:Pt:Ser:Ord
C0800571|PG IgG Ser Ql
C0800571|Phosphatidylglycerol IgG Ab [Presence] in Serum
C0800571|Phosphatidylglycerol Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C0943515|Protein C Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0943515|Protein C Ag actual/normal in Platelet poor plasma by Immunologic method
C0943515|Prot C Ag Act/Nor PPP Imm
C0943515|Protein C Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0943660|Fibrinogen fragments [Mass/volume] in Platelet poor plasma by Latex agglutination
C0943660|Fibrinogen Frg PPP LA-mCnc
C0943660|Fibrinogen fragments:MCnc:Pt:PPP:Qn:LA
C0943660|Fibrinogen fragments:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Latex Agglutination
C0482719|LMWH PPP Coag-aCnc
C0482719|Heparin.low molecular weight:ACnc:Pt:PPP:Qn:Coag
C0482719|LMW Heparin [Units/volume] in Platelet poor plasma by Coagulation assay
C0482719|Heparin.low molecular weight:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1317034|Coagulation surface induced.lupus sensitive.factor substitution^immediately after 1:2 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1317034|Coagulation surface induced.lupus sensitive.factor substitution^immediately after 1:2 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1317034|aPTT-LA imm 1:2 NP PPP
C1317034|aPTT.lupus sensitive.factor substitution in Platelet poor plasma by Coagulation assay --immediately after 1:2 addition of normal plasma
C0482661|Coagulation factor XIII Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482661|Fact XIII Ag PPP Imm-aCnc
C0482661|Coagulation factor XIII Ag:ACnc:Pt:PPP:Qn:Imm
C0482661|Coagulation factor XIII Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1114106|Fibrin+Fibrinogen fragments:MCnc:Pt:PPP:Qn
C1114106|Fibrin+Fibrinogen fragments [Mass/volume] in Platelet poor plasma
C1114106|FSP PPP-mCnc
C1114106|Fibrin+Fibrinogen fragments:Mass Concentration:Point in time:Platelet poor plasma:Quantitative
C1543007|INR in Platelet poor plasma or blood by Coagulation assay
C1543007|Coagulation tissue factor induced.INR:RelTime:Pt:PPP/Bld:Qn:Coag
C1543007|Coagulation tissue factor induced.INR:Relative Time:Point in time:Platelet poor plasma/Whole blood:Quantitative:Coagulation Assay
C1543007|INR PPP/Bld
C1544113|Coagulation surface induced^12H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544113|Coagulation surface induced^12 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544113|aPTT 12h p chal PPP
C1544113|aPTT in Platelet poor plasma by Coagulation assay --12 hours post XXX challenge
C0366909|vWf:RCo PPP-aCnc
C0366909|von Willebrand factor.ristocetin cofactor:ACnc:Pt:PPP:Qn
C0366909|von Willebrand factor (vWf) ristocetin cofactor [Units/volume] in Platelet poor plasma
C0366909|von Willebrand factor.ristocetin cofactor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C1714660|Lupus anticoagulant neutralization.buffer:Time:Pt:PPP:Qn:Coag
C1714660|Lupus anticoagulant neutralization buffer [Time] in Platelet poor plasma by Coagulation assay
C1714660|Lupus anticoagulant neutralization.buffer:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1714660|LA Nt Buffer PPP
C2361220|Maximum lysis.intrinsic coagulation system activated.heparin insensitive:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C2361220|ML.heparin insens LenFr Bld TEG
C2361220|Maximum lysis.intrinsic coagulation system activated.heparin insensitive:LenFr:Pt:Bld:Qn:Thromboelastography
C2361220|Maximum lysis.intrinsic coagulation system activated.heparin insensitive [Length fraction] in Blood by Thromboelastography
C2361222|Clotting time:Time:Pt:Bld:Qn:Thromboelastography
C2361222|Clotting time:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361222|Clotting time of Blood by Thromboelastography
C2361222|Clotting time Bld TEG
C1976976|Coagulation surface induced.factor substitution^1H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP:Qn:Coag
C1976976|Coagulation surface induced.factor substitution^1 hour post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1976976|aPTT 1h p 1:4 NP PPP
C1976976|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --1H post incubation with 1:4 normal plasma
C0482693|Coagulation tissue factor induced:Time:Pt:PPP^control:Qn:Coag
C0482693|Coagulation tissue factor induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482693|Prothrombin time (PT) in control Platelet poor plasma by Coagulation assay
C0482693|PT Cont PPP
C0482670|Deprecated Russell viper venom time in Platelet poor plasma by Coagulation assay
C0482670|Deprecated Coag RVV Ind PPP Qn
C0482670|Coagulation Russell viper venom induced:Time:Pt:PPP:Qn:Tilt tube
C0482670|Coagulation Russell viper venom induced:Time:Point in time:Platelet poor plasma:Quantitative:Tilt tube
C2733689|Phosphatidylserine Ab.IgG:MoM:Pt:Ser:Qn
C2733689|PS IgG MoM Ser
C2733689|Phosphatidylserine IgG Ab [Multiple of the median] in Serum
C2733689|Phosphatidylserine Antibody.immunoglobulin G:Multiple of the median:Point in time:Serum:Quantitative
C2733692|PA ADP 5 umol/L PRP Ql
C2733692|Platelet aggregation.adenosine diphosphate induced^5 umol/L:Pr:Pt:PRP:Ord
C2733692|Platelet aggregation.adenosine diphosphate induced^5 umol/L:Presence:Point in time:Platelet rich plasma:Ordinal
C2733692|Platelet aggregation ADP induced [Presence] in Platelet rich plasma --5 umol/L
C2733952|PA ADP ATP secr 10 umol/L Bld Ql
C2733952|Platelet aggregation ADP induced ATP secretion [Presence] in Blood --10 umol/L
C2733952|Platelet aggregation.adenosine diphosphate induced ATP secretion^10 umol/L:Pr:Pt:Bld:Ord
C2733952|Platelet aggregation.adenosine diphosphate induced ATP secretion^10 umol/L:Presence:Point in time:Whole blood:Ordinal
C2733740|Platelet aggregation arachidonate induced ATP secretion in Blood --500 umol/L
C2733740|PA AA ATP secr 500 umol/L Bld
C2733740|Platelet aggregation.arachidonate induced ATP secretion^500 umol/L:RelACnc:Pt:Bld:Qn
C2733740|Platelet aggregation.arachidonate induced ATP secretion^500 umol/L:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733963|PA Thromb ATP secr 1 U/mL Bld
C2733963|Platelet aggregation.thrombin induced ATP secretion^1 U/mL:Relative Arbitrary Concentration:Point in time:Whole blood:Quantitative
C2733963|Platelet aggregation thrombin induced ATP secretion in Blood --1 U/mL
C2733963|Platelet aggregation.thrombin induced ATP secretion^1 U/mL:RelACnc:Pt:Bld:Qn
C2708404|Coagulation surface induced.factor substitution^5M post incubation after addition of normal plasma:Time:Pt:PPP:Qn:Coag
C2708404|Coagulation surface induced.factor substitution^5 minutes post incubation after addition of normal plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2708404|aPTT 5M p NP PPP
C2708404|aPTT.factor substitution in Platelet poor plasma by Coagulation assay --5 minutes post incubation after addition of normal plasma
C3259775|Clot angle^after addition of heparinase:Angle:Pt:Bld:Qn:Thromboelastography
C3259775|Clot angle^after addition of heparinase:Angle:Point in time:Whole blood:Quantitative:Thromboelastography
C3259775|Clot angle in Blood by Thromboelastography --after addition of heparinase
C3259775|Clot angle Heparinase Bld TEG
C0365329|Coagulation dilute Russell viper venom induced:Time:Point in time:Platelet poor plasma:Quantitative:COAGULATION ASSAY
C0365329|Coagulation dilute Russell viper venom induced:Time:Pt:PPP:Qn:Coag
C0365329|dRVVT (LA screen)
C0365329|Screen dRVVT
C3654079|von Willebrand factor.activity:ACnc:Pt:PPP:Qn:Imm
C3654079|vWf:Ac PPP Imm-aCnc
C3654079|von Willebrand factor.activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C3654079|von Willebrand factor (vWf).activity [Units/volume] in Platelet poor plasma by Immunologic method
C2713203|Deprecated Cardiolipin IgG Ab [Units/volume] in Serum by Immunoassay
C2713203|Cardiolipin Ab.IgG:ACnc:Pt:Ser:Qn:EIA
C2713203|Deprecated Cardiolipin IgG Ser EIA-aCnc
C2713203|Cardiolipin Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C2713203|Deprecated Cardiolipin IgG Ab [Units/volume] in Serum by Immunoassay.
C0085278|Anti Phospholipid Syndrome
C0085278|Antiphospholipid Syndrome
C0085278|Syndrome, Anti-Phospholipid
C0085278|Syndrome, Antiphospholipid
C0085278|Anti Phospholipid Antibody Syndrome
C0085278|Antibody Syndrome, Anti-Phospholipid
C0085278|Antibody Syndrome, Antiphospholipid
C0085278|Antiphospholipid Antibody Syndromes
C0085278|Syndrome, Anti-Phospholipid Antibody
C0085278|Syndrome, Antiphospholipid Antibody
C0085278|antiphospholipid syndrome (diagnosis)
C0085278|Antiphospholipid Antibody Syndrome
C0085278|Anti-Phospholipid Syndrome
C0085278|Antiphospholipid Syndrome [Disease/Finding]
C0085278|Anti-Phospholipid Antibody Syndrome
C0085278|Anticardiolipin syndrome
C0085278|Antiphospholipid syndrome (disorder)
C0085278|Syndrome, Hughes
C0085278|Hughes Syndrome
C0085278|APL - Antiphospholipid syndrome
C0085278|APS - Antiphospholipid syndrome
C0085278|syndrome; anticardiolipin
C0085278|syndrome; antiphospholipid
C0085278|anticardiolipin; syndrome
C0085278|antiphospholipid; syndrome
C0799998|Fibrinopeptide A Ag:ACnc:Pt:PPP:Qn:Imm
C0799998|Fibrinopeptide A Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0799998|FpA Ag PPP Imm-aCnc
C0799998|Fibrinopeptide A Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0803902|Beta 2 glycoprotein 1 IgA Ab [Units/volume] in Serum
C0803902|Beta 2 glycoprotein 1 Ab.IgA:ACnc:Pt:Ser:Qn
C0803902|B2 Glycoprot1 IgA Ser-aCnc
C0803902|Beta 2 glycoprotein 1 Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Quantitative
C0803798|Coagulation factor VIII:Imp:Pt:XXX:Nom
C0803798|Fact VIII XXX-Imp
C0803798|Coagulation factor VIII:Impression/interpretation of study:Point in time:To be specified in another part of the message:Nominal
C0803798|Coagulation factor VIII [Interpretation] in Unspecified specimen
C0800586|PAI2 Ag PPP EIA-aCnc
C0800586|Plasminogen activator inhibitor 2 Ag:ACnc:Pt:PPP:Qn:EIA
C0800586|Plasminogen activator inhibitor 2 Ag [Units/volume] in Platelet poor plasma by Immunoassay
C0800586|Plasminogen activator inhibitor 2 Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C0881722|Platelet function (closure time) collagen+ADP induced [Time] in Blood
C0881722|Platelet function.collagen+Adenosine diphosphate induced:Time:Pt:Bld:Qn
C0881722|Platelet function.collagen+Adenosine diphosphate induced:Time:Point in time:Whole blood:Quantitative
C0881722|Closure Tme Coll+ADP Bld
C1316837|Streptokinase Ab [Titer] in Serum
C1316837|Streptokinase Ab Titr Ser
C1316837|Streptokinase Ab:Titr:Pt:Ser:Qn
C1316837|Streptokinase Antibody:Dilution Factor (Titer):Point in time:Serum:Quantitative
C0482704|Fibrin.soluble:ACnc:Pt:PPP:Qn:Chromo
C0482704|Fibrin Sol PPP Chro-aCnc
C0482704|Fibrin.soluble [Units/volume] in Platelet poor plasma by Chromogenic method
C0482704|Fibrin.soluble:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1316358|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --2 hours post incubation
C1316358|Coagulation tissue factor induced.factor substitution^2H post incubation:Time:Pt:PPP:Qn:Coag
C1316358|Coagulation tissue factor induced.factor substitution^2 hours post incubation:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1316358|PT 2h p Inc PPP
C1544098|Coagulation tissue factor induced^4H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544098|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --4 hours post XXX challenge
C1544098|Coagulation tissue factor induced^4 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544098|PT 4h p chal PPP
C1544641|Platelet factor 3:ACnc:Pt:PRP:Qn
C1544641|PF3 PRP-aCnc
C1544641|Platelet factor 3 [Units/volume] in Platelet rich plasma
C1544641|Platelet factor 3:Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1715673|B2 Glycoprot1 IgM SerPl EIA-aCnc
C1715673|Beta 2 glycoprotein 1 Ab.IgM:ACnc:Pt:Ser/Plas:Qn:EIA
C1715673|Beta 2 glycoprotein 1 IgM Ab [Units/volume] in Serum or Plasma by Immunoassay
C1715673|Beta 2 glycoprotein 1 Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:Enzyme Immunoassay
C2361161|dRVVT confirm PPP Ql
C2361161|Coagulation dilute Russell viper venom induced.excess phospholipid:ACnc:Pt:PPP:Ord:Coag
C2361161|Coagulation dilute Russell viper venom induced.excess phospholipid:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Coagulation Assay
C2361161|dRVVT excess phospholipid [Presence] in Platelet poor plasma by Coagulation assay
C2361184|Clot formation.extrinsic coagulation system activated:Time:Pt:Bld:Qn:Thromboelastography
C2361184|Clot formation.extrinsic coagulation system activated [Time] in Blood by Thromboelastography
C2361184|Clot formation.extrinsic coagulation system activated:Time:Point in time:Whole blood:Quantitative:Thromboelastography
C2361184|CFT.extrinsic Bld TEG
C1978979|Platelet aggregation.adenosine diphosphate induced^4 umol/L:Pr:Pt:PRP:Ord
C1978979|Platelet aggregation ADP induced [Presence] in Platelet rich plasma --4 umol/L
C1978979|PA ADP 4 umol/L PRP Ql
C1978979|Platelet aggregation.adenosine diphosphate induced^4 umol/L:Presence:Point in time:Platelet rich plasma:Ordinal
C1977231|PA Rist 1800 ug/mL PRP
C1977231|Platelet aggregation.ristocetin induced^1800 ug/mL:RelACnc:Pt:PRP:Qn
C1977231|Platelet aggregation.ristocetin induced^1800 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C1977231|Platelet aggregation ristocetin induced in Platelet rich plasma --1800 ug/mL
C1977082|Prot S Ag/Fact X Ag PPP
C1977082|Protein S Ag/Coagulation factor X Ag Ag [Mass Ratio] in Platelet poor plasma by Coagulation assay
C1977082|Protein S Ag/Coagulation factor X Ag:MRto:Pt:PPP:Qn:Coag
C1977082|Protein S Antigen/Coagulation factor X Antigen:Mass Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1977872|Platelet aggregation collagen induced [Identifier] in Platelet rich plasma
C1977872|Platelet aggregation.collagen induced:Prid:Pt:PRP:Nom
C1977872|Platelet aggregation.collagen induced:Presence or Identity:Point in time:Platelet rich plasma:Nominal
C1977872|PA Coll PRP Nom
C0482680|Coagulation thrombin induced:Time:Pt:PPP^control:Qn:Coag
C0482680|Coagulation thrombin induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482680|Thrombin time in control Platelet poor plasma by Coagulation assay
C0482680|TT Cont PPP
C2733664|Cardiolipin IgM Ab [Multiple of the median] in Serum
C2733664|Cardiolipin Ab.IgM:MoM:Pt:Ser:Qn
C2733664|Cardiolipin IgM MoM Ser
C2733664|Cardiolipin Antibody.immunoglobulin M:Multiple of the median:Point in time:Serum:Quantitative
C2733679|Lupus anticoagulant neutralization.high phospholipid.factor substitution^immediately after 1:2 addition of saline:Time:Pt:PPP:Qn:Coag
C2733679|Lupus anticoagulant neutralization high phospholipid.factor substitution [Time] in Platelet poor plasma by Coagulation assay --immediately after 1:2 addition of saline
C2733679|Lupus anticoagulant neutralization.high phospholipid.factor substitution^immediately after 1:2 addition of saline:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C2733679|LA Nt HPL imm 1:2 saline PPP
C2734631|B2 Glycoprot1 Ab Ser EIA-aCnc
C2734631|Beta 2 glycoprotein 1 Ab [Units/volume] in Serum by Immunoassay
C2734631|Beta 2 glycoprotein 1 Ab:ACnc:Pt:Ser:Qn:EIA
C2734631|Beta 2 glycoprotein 1 Antibody:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C0799996|Fibrinogen PPP Ql
C0799996|Fibrinogen:ACnc:Pt:PPP:Ord
C0799996|Fibrinogen [Presence] in Platelet poor plasma
C0799996|Fibrinogen:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C0797427|Phosphatidylcholine IgA Ab [Presence] in Serum
C0797427|Phosphatidylcholine Ab.IgA:ACnc:Pt:Ser:Ord
C0797427|PC IgA Ser Ql
C0797427|Phosphatidylcholine Antibody.immunoglobulin A:Arbitrary Concentration:Point in time:Serum:Ordinal
C0550591|Coagulation kaolin induced:ACnc:Pt:PPP:Qn
C0550591|Kaolin activated time [Units/volume] in Platelet poor plasma
C0550591|Coagulation kaolin induced:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0550591|KCT PPP-aCnc
C0550592|Fibrin+Fibrinogen fragments:ACnc:Pt:Urine:Qn
C0550592|FSP Ur-aCnc
C0550592|Fibrin+Fibrinogen fragments [Units/volume] in Urine
C0550592|Fibrin+Fibrinogen fragments:Arbitrary Concentration:Point in time:Urine:Quantitative
C0551332|PC IgM Ser-aCnc
C0551332|Phosphatidylcholine Ab.IgM:ACnc:Pt:Ser:Qn
C0551332|Phosphatidylcholine IgM Ab [Units/volume] in Serum
C0551332|Phosphatidylcholine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative
C0796784|PA PG PRP
C0796784|Platelet aggregation prostaglandin induced in Platelet rich plasma
C0796784|Platelet aggregation.prostaglandin induced:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0796784|Platelet aggregation.prostaglandin induced:RelACnc:Pt:PRP:Qn
C0943517|Prot S Ag Act/Nor PPP Imm
C0943517|Protein S Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0943517|Protein S Ag actual/normal in Platelet poor plasma by Immunologic method
C0943517|Protein S Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0943022|Cardiolipin Ab.IgG:ACnc:Pt:Ser:Ord
C0943022|Cardiolipin IgG Ser Ql
C0943022|Cardiolipin IgG Ab [Presence] in Serum
C0943022|Cardiolipin Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C0482718|Heparin neutralization:ACnc:Pt:PPP:Ord
C0482718|Heparin neutralization [Presence] in Platelet poor plasma
C0482718|Heparin Nt PPP Ql
C0482718|Heparin neutralization:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C1316355|Coagulation surface induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316355|Coagulation surface induced.factor substitution^immediately after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316355|aPTT imm 1:4 NP Cont PPP
C1316355|aPTT.factor substitution in control Platelet poor plasma by Coagulation assay --immediately after 1:4 addition of normal plasma
C0365326|Cardiolipin Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative:ENZYME IMMUNOASSAY
C0365326|Cardiolipin IgM Ser EIA-aCnc
C0365326|Cardiolipin IgM Ab [Units/volume] in Serum by Immunoassay
C0365326|Cardiolipin Ab.IgM:ACnc:Pt:Ser:Qn:EIA
C0482616|Fact Va PPP-aCnc
C0482616|Coagulation factor V activated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482616|Coagulation factor V activated activity:ACnc:Pt:PPP:Qn:Coag
C0482616|Coagulation factor V activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1147717|PS IgM Ser EIA-aCnc
C1147717|Phosphatidylserine Ab.IgM:ACnc:Pt:Ser:Qn:EIA
C1147717|Phosphatidylserine IgM Ab [Units/volume] in Serum by Immunoassay
C1147717|Phosphatidylserine Antibody.immunoglobulin M:Arbitrary Concentration:Point in time:Serum:Quantitative:Enzyme Immunoassay
C1544095|Coagulation tissue factor induced^1.5H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544095|Prothrombin time (PT) in Platelet poor plasma by Coagulation assay --1.5 hours post XXX challenge
C1544095|Coagulation tissue factor induced^1 1/2 hour post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544095|PT 1.5h p chal PPP
C1544106|Coagulation surface induced^1H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544106|Coagulation surface induced^1 hour post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544106|aPTT 1h p chal PPP
C1544106|aPTT in Platelet poor plasma by Coagulation assay --1 hour post XXX challenge
C1544114|Coagulation surface induced^1D post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544114|Coagulation surface induced^1 day post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544114|aPTT 1D p chal PPP
C1544114|aPTT in Platelet poor plasma by Coagulation assay --1 day post XXX challenge
C2361200|MCF Bld TEG
C2361200|Maximum clot firmness:Len:Pt:Bld:Qn:Thromboelastography
C2361200|Maximum clot firmness:Length:Point in time:Whole blood:Quantitative:Thromboelastography
C2361200|Maximum clot firmness [Length] in Blood by Thromboelastography
C2361732|Coagulation dilute Russell viper venom induced:Time:Pt:PPP^control:Qn:Coag
C2361732|Coagulation dilute Russell viper venom induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C2361732|dRVVT Cont PPP
C2361732|dRVVT in control Platelet poor plasma by Coagulation assay
C1953856|Kaolin activated time in Platelet poor plasma
C1953856|Coagulation kaolin induced:Time:Pt:PPP:Qn
C1953856|Coagulation kaolin induced:Time:Point in time:Platelet poor plasma:Quantitative
C1953856|KCT PPP
C2599019|PA AA Bld-aCnc
C2599019|Platelet aggregation.arachidonate induced:ACnc:Pt:Bld:Qn
C2599019|Platelet aggregation arachidonate induced [Units/volume] in Blood
C2599019|Platelet aggregation.arachidonate induced:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C3482455|Fibrin D-dimer FEU:MCnc:Pt:Bld:Qn:EIA
C3482455|Fibrin D-dimer FEU:Mass Concentration:Point in time:Whole blood:Quantitative:Enzyme Immunoassay
C3482455|Fibrin D-dimer FEU [Mass/volume] in Blood by Immunoassay
C3482455|D dimer FEU Bld EIA-mCnc
C0482717|Heparin cofactor II Ag:MCnc:Pt:PPP:Qn:Imm
C0482717|Heparin CF II Ag PPP Imm-mCnc
C0482717|Heparin cofactor II Ag [Mass/volume] in Platelet poor plasma by Immunologic method
C0482717|Heparin cofactor II Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1316439|Deprecated PAI1 Ag PPP EIA-mCnc
C1316439|Plasminogen activator inhibitor 1 Ag:MCnc:Pt:PPP:Qn:EIA
C1316439|Plasminogen activator inhibitor 1 Antigen:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Enzyme Immunoassay
C1316439|Deprecated Plasminogen activator inhibitor 1 Ag [Mass/volume] in Platelet poor plasma by EIA
C1316447|Coagulation factor X activity actual/Normal:RelCCnc:Pt:PPP:Qn:Chromo
C1316447|Coagulation factor X activity actual/normal in Platelet poor plasma by Chromogenic method
C1316447|Fact X Act/Nor PPP Chro
C1316447|Coagulation factor X activity actual/Normal:Relative Catalytic Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C1369580|INR Bld
C1369580|INR in Blood by Coagulation assay
C1369580|Coagulation tissue factor induced.INR:RelTime:Pt:Bld:Qn:Coag
C1369580|Coagulation tissue factor induced.INR:Relative Time:Point in time:Whole blood:Quantitative:Coagulation Assay
C0482663|Coagulation factor XIII coagulum dissolution:ACnc:Pt:PPP:Qn:Coag
C0482663|Fact XIII Clot Dis PPP-aCnc
C0482663|Coagulation factor XIII coagulum dissolution [Units/volume] in Platelet poor plasma by Coagulation assay
C0482663|Coagulation factor XIII coagulum dissolution:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1316346|Coagulation tissue factor induced.factor substitution^1H post incubation after 1:4 addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C1316346|Coagulation tissue factor induced.factor substitution^1 hour post incubation after 1:4 addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C1316346|Prothrombin time (PT) factor substitution in control Platelet poor plasma by Coagulation assay --1H post incubation with 1:4 normal plasma
C1316346|PT 1h p 1:4 NP Cont PPP
C0482626|Coagulation factor VII+Acarboxy Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482626|Fact VII+ACA Ag PPP Imm-aCnc
C0482626|Coagulation factor VII+Acarboxy Ag:ACnc:Pt:PPP:Qn:Imm
C0482626|Coagulation factor VII+Acarboxy Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0482648|Deprecated Fact Xia Fr PPP
C0482648|Coagulation factor XI activated activity:CFr:Pt:PPP:Qn:Coag
C0482648|Deprecated Coagulation factor XI activated activity
C0482648|Coagulation factor XI activated activity:Catalytic Fraction:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544108|Coagulation surface induced^2H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544108|Coagulation surface induced^2 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544108|aPTT 2h p chal PPP
C1544108|aPTT in Platelet poor plasma by Coagulation assay --2 hours post XXX challenge
C1716406|Low molecular weight heparin induced platelet Ab:ACnc:Pt:Ser:Ord
C1716406|Low molecular weight heparin induced platelet Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal
C1716406|LMW heparin (plat) Ab Ser Ql
C1716406|Low molecular weight heparin induced platelet Ab [Presence] in Serum
C0482768|Protein S.free Ag:ACnc:Pt:PPP:Qn:Imm
C0482768|Protein S Free Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482768|Prot S Free Ag PPP Imm-aCnc
C0482768|Protein S.free Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1714710|Cardiolipin IgM Ab [Mass/volume] in Serum
C1714710|Cardiolipin Ab.IgM:MCnc:Pt:Ser:Qn
C1714710|Cardiolipin IgM Ser-mCnc
C1714710|Cardiolipin Antibody.immunoglobulin M:Mass Concentration:Point in time:Serum:Quantitative
C1715177|AT III Ag PPP Ql Imm
C1715177|Antithrombin Ag:ACnc:Pt:PPP:Ord:Imm
C1715177|Antithrombin Ag [Presence] in Platelet poor plasma by Immunologic method
C1715177|Antithrombin Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Imm
C2361155|Prothrombin time (PT) PIVKA insensitive actual/normal in Capillary blood by Coagulation assay
C2361155|Coagulation tissue factor induced.PIVKA insensitive actual/Normal:RelTime:Pt:BldC:Qn:Coag
C2361155|PT PIVKA insensitive Act/Nor BldC
C2361155|Coagulation tissue factor induced.PIVKA insensitive actual/Normal:Relative Time:Point in time:Blood capillary:Quantitative:Coagulation Assay
C1978974|Deprecated Acarboxyprothrombin [Mass/volume] in Serum
C1978974|Acarboxyprothrombin:MCnc:Pt:Ser:Qn
C1978974|Deprecated Acarboxyprothrombin Ser-mCnc
C1978974|Acarboxyprothrombin:Mass Concentration:Point in time:Serum:Quantitative
C1954162|aPCR PPP-Imp
C1954162|Activated protein C resistance:Imp:Pt:PPP:Nom
C1954162|Activated protein C resistance:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal
C1954162|Activated protein C resistance [Interpretation] in Platelet poor plasma
C0482672|Deprecated Activated partial thrombplastin time (aPTT).factor substitution in Platelet poor plasma from control by Coagulation assay --20M post incubation with normal plasma
C0482672|Deprecated aPTT PPP Cont Qn
C0482672|Coagulation surface induced.factor substitution^20M post incubation.37 deg c after addition of normal plasma:Time:Pt:PPP^control:Qn:Tilt tube
C0482672|Coagulation surface induced.factor substitution^20 minutes post incubation.37 deg c after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Tilt tube
C0482732|Plasm Inhib Ag PPP Imm-aCnc
C0482732|Plasmin inhibitor Ag:ACnc:Pt:PPP:Qn:Imm
C0482732|Plasmin inhibitor Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482732|Plasmin inhibitor Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C2598477|Lupus anticoagulant neutralization.dilute phospholipid:Time:Pt:PPP:Qn
C2598477|Lupus anticoagulant neutralization dilute phospholipid [Time] in Platelet poor plasma
C2598477|Lupus anticoagulant neutralization.dilute phospholipid:Time:Point in time:Platelet poor plasma:Quantitative
C2598477|LA Nt dPL PPP
C2733691|PA ADP 2.5 umol/L PRP Ql
C2733691|Platelet aggregation ADP induced [Presence] in Platelet rich plasma --2.5 umol/L
C2733691|Platelet aggregation.adenosine diphosphate induced^2.5 umol/L:Pr:Pt:PRP:Ord
C2733691|Platelet aggregation.adenosine diphosphate induced^2.5 umol/L:Presence:Point in time:Platelet rich plasma:Ordinal
C2733695|PA Rist 500 mg/L PRP Ql
C2733695|Platelet aggregation.ristocetin induced^500 mg/L:ACnc:Pt:PRP:Ord
C2733695|Platelet aggregation ristocetin induced [Presence] in Platelet rich plasma --500 mg/L
C2733695|Platelet aggregation.ristocetin induced^500 mg/L:Arbitrary Concentration:Point in time:Platelet rich plasma:Ordinal
C2733961|PA Thromb ATP secr 5 U/mL Bld Ql
C2733961|Platelet aggregation thrombin induced ATP secretion [Presence] in Blood --5 U/mL
C2733961|Platelet aggregation.thrombin induced ATP secretion^5 U/mL:ACnc:Pt:Bld:Ord
C2733961|Platelet aggregation.thrombin induced ATP secretion^5 U/mL:Arbitrary Concentration:Point in time:Whole blood:Ordinal
C0482761|Protein C Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0482761|Protein C Ag:ACnc:Pt:PPP:Qn:Imm
C0482761|Prot C Ag PPP Imm-aCnc
C0482761|Protein C Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0484867|Fibrin D-dimer [Units/volume] in Platelet poor plasma
C0484867|D Dimer PPP-aCnc
C0484867|Fibrin D-dimer:ACnc:Pt:PPP:Qn
C0484867|Fibrin D-dimer:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative
C0799778|Coagulation surface induced:Time:Pt:Bld:Qn:Coag.saline 1:1
C0799778|Coagulation surface induced:Time:Point in time:Whole blood:Quantitative:Coagulation Assay.saline 1:1
C0799778|aPTT Bld 1:1 saline
C0799778|aPTT in Blood by Coagulation 1:1 saline
C0799999|Fibrinopeptide B Ag [Units/volume] in Platelet poor plasma by Immunologic method
C0799999|FpB Ag PPP Imm-aCnc
C0799999|Fibrinopeptide B Ag:ACnc:Pt:PPP:Qn:Imm
C0799999|Fibrinopeptide B Antigen:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0799776|Coagulation surface induced:Time:Point in time:Whole blood^Control:Quantitative:COAGULATION ASSAY
C0799776|Coagulation surface induced:Time:Pt:Bld^control:Qn:Coag
C0799776|aPTT Cont Bld
C0799776|aPTT in control Blood by Coagulation assay
C0803243|Phospholipid IgG Ser Ql
C0803243|Phospholipid Ab.IgG:ACnc:Pt:Ser:Ord
C0803243|Phospholipid IgG Ab [Presence] in Serum
C0803243|Phospholipid Antibody.immunoglobulin G:Arbitrary Concentration:Point in time:Serum:Ordinal
C0943516|Protein S Free Ag actual/normal in Platelet poor plasma by Immunologic method
C0943516|Prot S Free Ag Act/Nor PPP Imm
C0943516|Protein S.free Ag actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0943516|Protein S.free Antigen actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C0944234|Plasmin inhibitor actual/Normal:RelMCnc:Pt:PPP:Qn:Imm
C0944234|Plasmin inhibitor actual/normal in Platelet poor plasma by Immunologic method
C0944234|Plasm Inhib Act/Nor PPP Imm
C0944234|Plasmin inhibitor actual/Normal:Relative Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Imm
C1317050|von Willebrand factor cleaving protease:ACnc:Pt:PPP:Ord
C1317050|von Willebrand factor (vWf) cleaving protease [Presence] in Platelet poor plasma
C1317050|vWF Cp PPP Ql
C1317050|von Willebrand factor cleaving protease:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal
C0482699|Deprecated Fibrin D-dimer:Mass Concentration:Point in time:Platelet poor plasma:Ordinal:LATEX AGGLUTINATION
C0482699|Deprecated D Dimer PPP Ql LA
C0482699|Fibrin D-dimer:MCnc:Pt:PPP:Ord:LA
C0482699|Fibrin D-dimer:Mass Concentration:Point in time:Platelet poor plasma:Ordinal:Latex Agglutination
C0482699|Deprecated Fibrin D-dimer by agglutination
C0482702|Fibrin monomer:ACnc:Pt:PPP:Qn:LA
C0482702|Fibrin monomer [Units/volume] in Platelet poor plasma by Latex agglutination
C0482702|Fibrin Monomer PPP LA-aCnc
C0482702|Fibrin monomer:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Latex Agglutination
C1315826|Prothrombin time (PT) factor substitution in Platelet poor plasma by Coagulation assay --1 hour post incubation
C1315826|Coagulation tissue factor induced.factor substitution^1H post incubation:Time:Pt:PPP:Qn:Coag
C1315826|Coagulation tissue factor induced.factor substitution^1 hour post incubation:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1315826|PT 1h p Inc PPP
C1315992|PA Rist lo dose PRP
C1315992|Platelet aggregation.ristocetin induced^low dose:RelACnc:Pt:PRP:Qn
C1315992|Platelet aggregation ristocetin induced in Platelet rich plasma --Low dose
C1315992|Platelet aggregation.ristocetin induced^low dose:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C0365444|Heparin Ab:Threshold:Pt:Ser:Qn:Platelet aggr
C0365444|Heparin Ab Ser Qn Pl Agg
C0365444|Heparin Ab [Threshold] in Serum by Platelet aggregation
C0365444|Heparin Antibody:Threshold:Point in time:Serum:Quantitative:Platelet aggr
C0482610|Coagulation factor IX activated [Units/volume] in Platelet poor plasma by Coagulation assay
C0482610|Fact IXa PPP-aCnc
C0482610|Coagulation factor IX activated activity:ACnc:Pt:PPP:Qn:Coag
C0482610|Coagulation factor IX activated activity:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544112|Coagulation surface induced^8H post XXX challenge:Time:Pt:PPP:Qn:Coag
C1544112|Coagulation surface induced^8 hours post XXX challenge:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C1544112|aPTT 8h p chal PPP
C1544112|aPTT in Platelet poor plasma by Coagulation assay --8 hours post XXX challenge
C1544432|Prothrom Ab SerPl-aCnc
C1544432|Prothrombin Ab [Units/volume] in Serum or Plasma
C1544432|Prothrombin Ab:ACnc:Pt:Ser/Plas:Qn
C1544432|Prothrombin Antibody:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C1623603|Cardiolipin Ab.IgG.B2GP1 independent:MoM:Pt:Ser:Qn
C1623603|Cardiolipin IgG B2GP1 indep MoM Ser
C1623603|Cardiolipin IgG Ab B2GP1 independent [Multiple of the median] in Serum
C1623603|Cardiolipin Antibody.immunoglobulin G.B2GP1 independent:Multiple of the median:Point in time:Serum:Quantitative
C1978603|Fact XIII Inhib PPP Ql Chro
C1978603|Coagulation factor XIII inhibitor:ACnc:Pt:PPP:Ord:Chromo
C1978603|Coagulation factor XIII inhibitor [Presence] in Platelet poor plasma by Chromogenic method
C1978603|Coagulation factor XIII inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Ordinal:Chromogenic/Enzymatic Assay
C1978977|PA ADP 20 umol/L PRP Ql
C1978977|Platelet aggregation.adenosine diphosphate induced^20 umol/L:Pr:Pt:PRP:Ord
C1978977|Platelet aggregation ADP induced [Presence] in Platelet rich plasma --20 umol/L
C1978977|Platelet aggregation.adenosine diphosphate induced^20 umol/L:Presence:Point in time:Platelet rich plasma:Ordinal
C0482666|Deprecated Reptilase PPP Cont Qn
C0482666|Deprecated Reptilase time in Platelet poor plasma from control by Coagulation assay
C0482666|Coagulation reptilase induced:Time:Pt:PPP^control:Qn:Tilt tube
C0482666|Coagulation reptilase induced:Time:Point in time:Platelet poor plasma^Control:Quantitative:Tilt tube
C0482687|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Pt:PPP^control:Qn:Coag
C0482687|Coagulation tissue factor induced.factor substitution^immediately after addition of normal plasma:Time:Point in time:Platelet poor plasma^Control:Quantitative:Coagulation Assay
C0482687|Prothrombin time (PT) factor substitution in control Platelet poor plasma by Coagulation assay --immediately after addition of normal plasma
C0482687|PT imm NP Cont PPP
C3259332|Clot firmness^30 minutes after maximum clot amplitude after addition of heparinase:Length Fraction:Point in time:Whole blood:Quantitative:Thromboelastography
C3259332|CF 30M p MA after hepase LenFr Bld TEG
C3259332|Clot firmness^30M after maximum clot amplitude after addition of heparinase:LenFr:Pt:Bld:Qn:Thromboelastography
C3259332|Clot firmness [Length fraction] in Blood by Thromboelastography --30 minutes after maximum clot amplitude after addition of heparinase
C0482749|Plasminogen activator tissue type:MCnc:Pt:PPP:Qn:Chromo
C0482749|tPA PPP Chro-mCnc
C0482749|Plasminogen activator tissue type [Mass/volume] in Platelet poor plasma by Chromogenic method
C0482749|Plasminogen activator tissue type:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3699650|Dabigatran:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3699650|Dabigatran PPP-mCnc
C3699650|Dabigatran:MCnc:Pt:PPP:Qn:Coag
C3699650|Dabigatran [Mass/volume] in Platelet poor plasma by Coagulation assay
C3481607|Rivaroxaban [Units/volume] in Platelet poor plasma by Chromogenic method
C3481607|Rivaroxaban:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3481607|Rivaroxaban:ACnc:Pt:PPP:Qn:Chromo
C3481607|Rivaroxaban PPP Chro-aCnc
C0373776|Clotting; factor VIII, VW factor antigen
C0373776|Clotting; factor VIII, VW factor antigen (procedure)
C0373776|CLOTTING FACTOR VIII VW FACTOR ANTIGEN
C0373776|CLOT FACTOR VIII VW ANTIGEN
C0373776|Clotting factor VIII (VW factor) antigen
C0200411|Clotting factor XII assay
C0200411|factor XII assay (lab test)
C0200411|factor XII assay
C0200411|factor XII level
C0200411|Clotting; factor XII (Hageman)
C0200411|CLOTTING FACTOR XII HAGEMAN
C0200411|Assay for clotting factor XII (Hageman)
C0200411|CLOT FACTOR XII HAGEMAN
C0200411|Clotting factor XII (Hageman) measurement
C0200411|Hageman factor assay
C0200411|Clotting factor XII assay (procedure)
C0200398|factor VII assay
C0200398|factor VII assay (lab test)
C0200398|factor VII level
C0200398|Clotting; factor VII (proconvertin, stable factor)
C0200398|CLOTTING FACTOR VII PROCONVERTIN STABLE FACTOR
C0200398|Assay for clotting factor VII
C0200398|Clotting factor VII (proconvertin, stable factor)
C0200398|CLOT FACTOR VII PROCONVERTIN
C0200398|Plasma factor VII level (procedure)
C0200398|Plasma factor VII level
C0200398|Clotting factor VII assay
C0200398|Stable factor assay
C0200398|Proconvertin assay
C0200398|Autoprothrombin I assay
C0200398|Clotting factor VII assay (procedure)
C0200398|Plasma factor VII level assay
C0200405|Factor VIII assay, one stage (procedure)
C0200405|Clotting; factor VIII (AHG), 1-stage
C0200405|CLOTTING FACTOR VIII AHG 1 STAGE
C0200405|Clotting factor VIII (AHG) measurement
C0200405|1-stage assay for clotting factor VIII (AHG)
C0200405|CLOT FACTOR VIII AHG 1 STAGE
C0200405|Factor VIII assay, one stage
C0373775|Clotting; factor VIII, VW factor, ristocetin cofactor
C0373775|Clotting; factor VIII, VW factor, ristocetin cofactor (procedure)
C0373775|CLOTTING FACTOR VIII VW FACTOR RISTOCETIN COFACT
C0373775|CLOT FACTOR VIII VW RISTOCTN
C0373778|Clotting; factor XIII (fibrin stabilizing), screen solubility
C0373778|CLOTTING FACTOR XIII FIBRN STABILIZ SCREEN SOLUB
C0373778|Clotting factor XIII (fibrin stabilizing) screening test
C0373778|CLOT FACTOR XIII FIBRIN SCRN
C0373778|Solubility screening for clotting factor XIII (fibrin stabilizing)
C0200396|Clotting factor II assay
C0200396|Clotting; factor II, prothrombin, specific
C0200396|Prothrombin level
C0200396|factor II assay
C0200396|factor II assay (lab test)
C0200396|factor II level
C0200396|Prothrombin.activity
C0200396|Prothrombin Measurement
C0200396|Assay for clotting factor II
C0200396|CLOTTING FACTOR II PROTHROMBIN SPECIFIC
C0200396|Clotting factor II prothrombin, measurement
C0200396|CLOT FACTOR II PROTHROM SPEC
C0200396|Factor II level (procedure)
C0200396|Factor II
C0200396|Prothrombin
C0200396|FACTII
C0200396|Coagulation factor II level
C0200396|Prothrombin activity
C0200396|Prothrombin assay
C0200396|Clotting factor II assay (procedure)
C0200409|Clotting factor X assay
C0200409|factor X assay
C0200409|factor X assay (lab test)
C0200409|factor X level
C0200409|Clotting; factor X (Stuart-Prower)
C0200409|CLOTTING FACTOR X STUART-PROWER
C0200409|CLOT FACTOR X STUART-POWER
C0200409|Clotting factor X (Stuart-Prower) measurement
C0200409|Assay for clotting factor X (Stuart-Prower)
C0200409|Plasma factor X level (procedure)
C0200409|Plasma factor X level
C0200409|Stuart factor assay
C0200409|Stuart-Prower factor assay
C0200409|Clotting factor X assay (procedure)
C0200410|Clotting factor XI assay
C0200410|factor XI assay
C0200410|factor XI assay (lab test)
C0200410|factor XI level
C0200410|Clotting; factor XI (PTA)
C0200410|CLOTTING FACTOR XI PTA
C0200410|Clotting factor XI (PTA) measurement
C0200410|CLOT FACTOR XI PTA
C0200410|Assay for clotting factor XI (PTA)
C0200410|Plasma factor XI level (procedure)
C0200410|Plasma factor XI level
C0200410|Plasma thromboplastin antecedent assay
C0200410|PTA assay
C0200410|Clotting factor XI assay (procedure)
C0200415|Fletcher factor assay (procedure)
C0200415|Fletcher's factor assay (lab test)
C0200415|prekallikrein Assay
C0200415|Fletcher's factor assay
C0200415|Fletcher's factor level
C0200415|Clotting; prekallikrein assay (Fletcher factor assay)
C0200415|CLOTTING PREKALLIKREIN ASSAY FLETCHER FACT ASSAY
C0200415|Assay for prekallikrein (Fletcher factor)
C0200415|Fletcher factor (clotting factor) measurement
C0200415|CLOT FACTOR FLETCHER FACT
C0200415|Fletcher factor assay
C0427597|factor XIII assay (lab test)
C0427597|factor XIII assay
C0427597|Clotting; factor XIII (fibrin stabilizing)
C0427597|CLOTTING FACTOR XIII FIBRIN STABILIZING
C0427597|CLOT FACTOR XIII FIBRIN STAB
C0427597|Clotting factor XIII (fibrin stabilizing) measurement
C0427597|Assay for clotting factor XIII (fibrin stabilizing)
C0427597|Clotting factor XIII assay
C0427597|Fibrinoligase assay
C0427597|Laki-Lorand factor assay
C0427597|Fibrin stabilizing factor assay
C0427597|Factor XIII activity
C0427597|Factor XIII level
C0427597|Clotting factor XIII assay (procedure)
C0427597|Fibrin stabilising factor assay
C0373777|Clotting; factor VIII, von Willebrand factor, multimetric analysis
C0373777|CLOTTING FACTOR VIII MULTIMETRIC ANALYSIS
C0373777|CLOT FACTOR VIII MULTIMETRIC
C0427584|Clotting; factor VIII related antigen
C0427584|CLOTTING FACTOR VIII RELATED ANTIGEN
C0427584|Clotting factor VIII related antigen measurement
C0427584|CLOT FACTOR VIII RELTD ANTGN
C0427584|Assay for clotting factor VIII-related antigen
C0427584|Clotting factor VIII (VW factor) measurement
C0427584|Factor VIII R: Ag assay
C0427584|Factor VIII related antigen assay
C0427584|RAg - Factor VIII related antigen level
C0427584|Factor VIII R: Ag assay (procedure)
C0427584|Blood clot factor VIII test
C0427592|Clotting; factor V (AcG or proaccelerin), labile factor
C0427592|factor V assay (lab test)
C0427592|factor V assay
C0427592|factor V level
C0427592|CLOTTING FACTOR V ACG/PROACCELERIN LABILE FACTOR
C0427592|Clotting factor V (ACP or proaccelerin) measurement
C0427592|Assay for clotting factor V (AcG or proaccelerin)
C0427592|BLOOC CLOT FACTOR V TEST
C0427592|Clotting factor V assay
C0427592|Labile factor assay
C0427592|Proaccelerin assay
C0427592|Ac-Globulin assay
C0427592|Clotting factor V assay (procedure)
C0427592|Plasma factor V level
C0200414|Fitzgerald factor assay (procedure)
C0200414|Fitzgerald's factor assay
C0200414|Fitzgerald's factor assay (lab test)
C0200414|Fitzgerald's factor level
C0200414|Clotting; high molecular weight kininogen assay (Fitzgerald factor assay)
C0200414|CLOTTING HI MOLEC WEIGHT KININOGEN ASSAY
C0200414|Assay for high molecular weight kininogen (Fitzgerald factor)
C0200414|CLOT FACTOR WGHT KININOGEN
C0200414|Fitzgerald factor (clotting factor) measurement
C0200414|Fitzgerald factor assay
C0200414|High molecular weight kininogen assay
C0200414|HMW kininogen assay
C0200414|Williams-Fitzgerald Flaujeac factor assay
C3813128|FACTXIII
C3813128|Factor XIII
C3813128|Factor XIII Measurement
C3813128|Fibrin Stablizing Factor
C3827252|Clot Detection
C3259781|Coagulation Index
C3259781|CI
C3259781|COAGIDX
C3259781|Coagulation Index Measurement
C3274476|Activated PTT/Standard Ratio Measurement
C3274476|Activated Partial Thromboplastin Time/Standard Thromboplastin Time
C3274476|APTTSTND
C3274476|Activated PTT/Standard
C3274476|Activated PTT/Standard PTT
C3274476|Activated PTT to Standard PTT Ratio Measurement
C3820394|Thrombin/Antithrombin
C3820394|Thrombin to Antithrombin Ratio Measurement
C3820394|Thrombin/Antithrombin III
C3820394|TAT
C3847087|Rivaroxaban:MCnc:Pt:PPP:Qn:Chromo
C3847087|Rivaroxaban [Mass/volume] in Platelet poor plasma by Chromogenic method
C3847087|Rivaroxaban PPP Chro-mCnc
C3847087|Rivaroxaban:Mass Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C3847420|von Willebrand factor.activity actual/Normal^immediately after 1:1 addition of normal plasma:Relative Ratio:Point in time:Platelet poor plasma:Quantitative:Imm
C3847420|vWf:Ac Act/Nor imm 1:1 NP PPP Imm
C3847420|von Willebrand factor.activity actual/Normal^immediately after 1:1 addition of normal plasma:RelRto:Pt:PPP:Qn:Imm
C3847420|von Willebrand factor (vWf).activity actual/normal in Platelet poor plasma by Immunologic method --immediately after 1:1 addition of normal plasma
C3847419|vWf:Ac Act/Nor PPP Cont Imm
C3847419|von Willebrand factor.activity actual/Normal:Relative Ratio:Point in time:Platelet poor plasma^Control:Quantitative:Imm
C3847419|von Willebrand factor.activity actual/Normal:RelRto:Pt:PPP^control:Qn:Imm
C3847419|von Willebrand factor (vWf).activity actual/normal in control Platelet poor plasma by Immunologic method
C3870346|Coagulation surface induced.lupus sensitive percent correction:PctDiff:Pt:PPP:Qn:Coag
C3870346|aPTT.lupus sensitive W excess phospholipid percent correction
C3870346|Coagulation surface induced.lupus sensitive percent correction:Percent difference:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870346|aPTT % correction
C3870036|aPTT screen to confirm ratio
C3870036|Coagulation surface induced.lupus sensitive/Coagulation surface induced.lupus sensitive.excess phospholipid:Ratio:Pt:PPP:Qn:Coag
C3870036|Coagulation surface induced.lupus sensitive/Coagulation surface induced.lupus sensitive.excess phospholipid:Ratio:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870036|aPTT.lupus sensitive/aPTT.lupus sensitive W excess phospholipid (screen to confirm ratio)
C3870347|Coagulation surface induced.lupus sensitive.excess phospholipid:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870347|Coagulation surface induced.lupus sensitive.excess phospholipid:Time:Pt:PPP:Qn:Coag
C3870347|Confirm aPTT
C3870347|aPTT.lupus sensitive W excess phospholipid (LA confirm)
C3870344|Coagulation surface induced.lupus sensitive with 1:1 Pooled Normal Plasma actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3870344|aPTT.lupus sensitive with 1:1 PNP actual/Normal (normalized LA mix)
C3870344|Mixing aPTT/normal
C3870344|Coagulation surface induced.lupus sensitive with 1:1 Pooled Normal Plasma actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870339|Lupus anticoagulant two screening tests W Reflex [interpretation]
C3870339|Lupus anticoagulant two screening tests W Reflex:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal:Coagulation Assay
C3870339|Lupus anticoagulant two screening tests W Reflex:Imp:Pt:PPP:Nom:Coag
C3870339|LA 2 screen W Reflex-Imp
C3870038|LA 3 screen W Reflex-Imp
C3870038|Lupus anticoagulant three screening tests W Reflex:Imp:Pt:PPP:Nom:Coag
C3870038|Lupus anticoagulant three screening tests W Reflex [interpretation]
C3870038|Lupus anticoagulant three screening tests W Reflex:Impression/interpretation of study:Point in time:Platelet poor plasma:Nominal:Coagulation Assay
C3870010|dRVVT.hexagonal phase phospholipid actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3870010|dRVVT.hexagonal phase phospholipid actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870010|dRVVT W excess hexagonal phospholipid/Normal (StaClot LA confirm)
C3870010|Normalized confirm dRVVT StaClot
C3870343|Coagulation surface induced.lupus sensitive with 1:1 Pooled Normal Plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870343|Mixing aPTT
C3870343|aPTT.lupus sensitive with 1:1 PNP (LA mix)
C3870343|Coagulation surface induced.lupus sensitive with 1:1 Pooled Normal Plasma:Time:Pt:PPP:Qn:Coag
C3870092|Coagulation surface induced.hexagonal phase phospholipid actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870092|Coagulation surface induced.hexagonal phase phospholipid actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3870092|aPTT W hexagonal phospholipid/Normal (StaClot LA confirm)
C3870092|Normalized confirm aPTT StaClot
C3870000|Delta dRVVT:Time Difference:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870000|Delta dRVVT [Time] in Platelet poor plasma by Coagulation assay
C3870000|Delta dRVVT PPP
C3870000|Delta dRVVT:TimeDif:Pt:PPP:Qn:Coag
C3870342|DRVVT percent correction:PctDiff:Pt:PPP:Qn:Coag
C3870342|dRVVT W excess phospholipid percent correction
C3870342|dRVVT % correction
C3870342|DRVVT percent correction:Percent difference:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870341|dRVVT with 1:1 PNP actual/normal (normalized LA mix)
C3870341|DRVVT with 1:1 Pooled Normal Plasma actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3870341|Mixing dRVVT/normal
C3870341|DRVVT with 1:1 Pooled Normal Plasma actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870340|Mixing dRVVT
C3870340|DRVVT with 1:1 Pooled Normal Plasma:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870340|DRVVT with 1:1 Pooled Normal Plasma:Time:Pt:PPP:Qn:Coag
C3870340|dRVVT with 1:1 PNP (LA mix)
C3870037|dRVVT W excess hexagonal phospholipid (STA-StaClot confirm)
C3870037|dRVVT.hexagonal phase phospholipid:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3870037|dRVVT.hexagonal phase phospholipid:Time:Pt:PPP:Qn:Coag
C3870037|Confirm dRVVT STA-StaClot
C3869999|Delta aPTT PPP
C3869999|Delta aPTT:Time Difference:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C3869999|Delta aPTT:TimeDif:Pt:PPP:Qn:Coag
C3869999|Delta aPTT [Time] in Platelet poor plasma by Coagulation assay
C3870345|Confirm aPTT/normal
C3870345|Coagulation surface induced.lupus sensitive.excess phospholipid actual/Normal:RelTime:Pt:PPP:Qn:Coag
C3870345|aPTT.lupus sensitive W excess phospholipid actual/Normal (normalized LA confirm)
C3870345|Coagulation surface induced.lupus sensitive.excess phospholipid actual/Normal:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C4036712|Thrombin activatable fibrinolysis inhibitor:ACnc:Pt:PPP:Qn:Chromo
C4036712|Thrombin activatable fibrinolysis inhibitor [Units/volume] in Platelet poor plasma by Chromogenic method
C4036712|Thrombin activatable fibrinolysis inhibitor:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Chromogenic/Enzymatic Assay
C4036712|TAFI PPP Chro-aCnc
C4037141|Prothrombin.activity^immediately after addition of factor II depleted plasma:Arbitrary Concentration:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C4037141|Prothrombin.activity^immediately after addition of factor II depleted plasma:ACnc:Pt:PPP:Qn:Coag
C4037141|Prothrom imm FII DP PPP-aCnc
C4037141|Prothrombin activity [Units/volume] in Platelet poor plasma by Coagulation assay --immediately after addition of factor II depleted plasma
C4053801|Factor X Activity
C4053801|Factor X Activity Measurement
C4053801|FACTXA
C1271799|von Willebrand factor activity
C1271799|von Willebrand factor activity (procedure)
C1271799|FACTVWA
C1271799|von Willebrand Factor Activity Measurement
C1271799|Von Willebrand factor activity level
C1271799|Von Willebrand factor activity measurement (procedure)
C1294019|blood alpha-2 antiplasmin activity (lab test)
C1294019|blood alpha-2 antiplasmin activity
C1294019|alpha-2 antiplasmin activity
C1294019|Alpha-2 antiplasmin functional assay
C1294019|Alpha 2 antiplasmin activity
C1294019|Alpha 2 antiplasmin activity (procedure)
C1294019|Alpha-2 Antiplasmin Activity Measurement
C1294019|APLSMA2A
C1294019|Alpha-2 antiplasmin functional assay (procedure)
C4070996|PA Coll 5 ug/mL PRP
C4070996|Platelet aggregation.collagen induced^5 ug/mL:RelACnc:Pt:PRP:Qn
C4070996|Platelet aggregation.collagen induced^5 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070996|Platelet aggregation collagen induced in Platelet rich plasma --5 ug/mL
C4070995|Platelet aggregation.ristocetin induced^1.25 mg/mL:RelACnc:Pt:PRP:Qn
C4070995|PA Rist 1.25 mg/ml PRP
C4070995|Platelet aggregation.ristocetin induced^1.25 mg/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070995|Platelet aggregation ristocetin induced in Platelet rich plasma --1.25 mg/ml
C4071002|Platelet aggregation ADP induced in Platelet rich plasma --4 umol/L
C4071002|Platelet aggregation.adenosine diphosphate induced^4 umol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4071002|Platelet aggregation.adenosine diphosphate induced^4 umol/L:RelACnc:Pt:PRP:Qn
C4071002|PA ADP 4 umol/L PRP
C4071001|Platelet aggregation ADP induced in Platelet rich plasma --5 umol/L
C4071001|Platelet aggregation.adenosine diphosphate induced^5 umol/L:RelACnc:Pt:PRP:Qn
C4071001|PA ADP 5 umol/L PRP
C4071001|Platelet aggregation.adenosine diphosphate induced^5 umol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070999|Platelet aggregation.epinephrine induced^6 umol/L:RelACnc:Pt:PRP:Qn
C4070999|Platelet aggregation epinephrine induced in Platelet rich plasma --6 umol/L
C4070999|Platelet aggregation.epinephrine induced^6 umol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070999|PA Epineph 6 umol/L PRP
C4070903|PA Rist hi dose Bld-aCnc
C4070903|Platelet aggregation ristocetin induced [Units/volume] in Blood --High dose
C4070903|Platelet aggregation.ristocetin induced^high dose:ACnc:Pt:Bld:Qn
C4070903|Platelet aggregation.ristocetin induced^high dose:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C4070853|Platelet aggregation ristocetin induced [Units/volume] in Blood --Low dose
C4070853|Platelet aggregation.ristocetin induced^low dose:ACnc:Pt:Bld:Qn
C4070853|Platelet aggregation.ristocetin induced^low dose:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C4070853|PA Rist lo dose Bld-aCnc
C4070997|PA Coll 1.25 ug/ml PRP
C4070997|Platelet aggregation.collagen induced^1.25 ug/mL:RelACnc:Pt:PRP:Qn
C4070997|Platelet aggregation.collagen induced^1.25 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070997|Platelet aggregation collagen induced in Platelet rich plasma --1.25 ug/ml
C4070901|Platelet aggregation adenosine diphosphate+prostaglandin E1 induced [Units/volume] in Blood
C4070901|Platelet aggregation.adenosine diphosphate+prostaglandin E1 induced:ACnc:Pt:Bld:Qn
C4070901|Platelet aggregation.adenosine diphosphate+prostaglandin E1 induced:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C4070901|PA ADP+PGE1 induced Bld-aCnc
C4070432|Platelet aggregation.ristocetin induced^500 ug/mL:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070432|Platelet aggregation.ristocetin induced^500 ug/mL:RelACnc:Pt:PRP:Qn
C4070432|Platelet aggregation ristocetin induced in Platelet rich plasma --500 ug/mL
C4070432|PA Rist 500 ug/mL PRP
C4070398|Platelet aggregation.adenosine diphosphate induced^10 umol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070398|PA ADP 10 umol/L PRP
C4070398|Platelet aggregation ADP induced in Platelet rich plasma --10 umol/L
C4070398|Platelet aggregation.adenosine diphosphate induced^10 umol/L:RelACnc:Pt:PRP:Qn
C4069315|Clotting time of depleted plasma with 1:1 phospholipid^after addition of factor X activated:Time:Pt:PPP:Qn:Coag
C4069315|PPL p Fxa PPP
C4069315|Clotting time of depleted plasma with 1:1 phospholipid by Coagulation assay --after addition of factor X activated
C4069315|Clotting time of depleted plasma with 1:1 phospholipid^after addition of factor X activated:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C4071003|Platelet aggregation.adenosine diphosphate induced^2.5 umol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4071003|Platelet aggregation ADP induced in Platelet rich plasma --2.5 umol/L
C4071003|Platelet aggregation.adenosine diphosphate induced^2.5 umol/L:RelACnc:Pt:PRP:Qn
C4071003|PA ADP 2.5 umol/L PRP
C4071000|PA Epineph 100 umol/L PRP
C4071000|Platelet aggregation.epinephrine induced^100 umol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4071000|Platelet aggregation.epinephrine induced^100 umol/L:RelACnc:Pt:PRP:Qn
C4071000|Platelet aggregation epinephrine induced in Platelet rich plasma --100 umol/L
C4070998|PA AA 1.6 mmol/L PRP
C4070998|Platelet aggregation.arachidonate induced^1.6 mmol/L:RelACnc:Pt:PRP:Qn
C4070998|Platelet aggregation.arachidonate induced^1.6 mmol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4070998|Platelet aggregation arachidonate induced in Platelet rich plasma --1.6 mmol/L
C4070904|PA Coll Bld-aCnc
C4070904|Platelet aggregation collagen induced [Units/volume] in Blood
C4070904|Platelet aggregation.collagen induced:ACnc:Pt:Bld:Qn
C4070904|Platelet aggregation.collagen induced:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C4071004|Platelet aggregation.adenosine diphosphate induced^2 umol/L:Relative Arbitrary Concentration:Point in time:Platelet rich plasma:Quantitative
C4071004|Platelet aggregation ADP induced in Platelet rich plasma --2 umol/L
C4071004|PA ADP 2 umol/L PRP
C4071004|Platelet aggregation.adenosine diphosphate induced^2 umol/L:RelACnc:Pt:PRP:Qn
C4070902|Platelet aggregation thrombin receptor activating peptide-6 induced [Units/volume] in Blood
C4070902|Platelet aggregation.thrombin receptor activating peptide-6 induced:Arbitrary Concentration:Point in time:Whole blood:Quantitative
C4070902|Platelet aggregation.thrombin receptor activating peptide-6 induced:ACnc:Pt:Bld:Qn
C4070902|PA TRAP-6 induced Bld-aCnc
C0200435|Clotting test with substitution
C0200435|Substituted clotting test
C0200435|Clotting test, mixtures
C0200435|Clotting test with substitution (procedure)
C0200435|Clotting test with substitution, NOS
C0200435|Substituted clotting test, NOS
C0200435|Clotting test, mixtures, NOS
C0200493|Blood coagulation panel, disseminated intravascular coagulation
C0200493|Blood coagulation panel, disseminated intravascular coagulation (procedure)
C0200493|Blood coagulation panel, DIC (procedure)
C0200493|Blood coagulation panel, DIC
C0200493|Consumptive coagulopathy screen
C0200493|Disseminated intravascular coagulation screening panel
C0200493|DIC screen
C0200493|DIC - Disseminated intravascular coagulation screen
C0200493|Disseminated intravascular coagulation screening
C0200494|Coagulation panel for thrombosis
C0200494|Thrombosis panel
C0200494|Hypercoagulable state screen
C0200494|Coagulation panel for thrombosis (procedure)
C0581145|Plasma activated protein C resistance (procedure)
C0581145|Plasma activated protein C resistance
C1273350|Advanced coagulation studies (procedure)
C1273350|Advanced coagulation studies
C1273381|Kaolin clotting time Rosner index (procedure)
C1273381|Kaolin clotting time Rosner index
C1273438|kaolin clotting time (lab test)
C1273438|kaolin clotting time
C1273438|Kaolin clotting time (procedure)
C1319568|Factor V(306) Cambridge mutation test (procedure)
C1319568|Factor V(306) Cambridge mutation test
C1272307|Target international normalized ratio (observable entity)
C1272307|Target international normalised ratio (observable entity)
C1272307|Target international normalised ratio
C1272307|Target international normalised ratio (procedure)
C1272307|INR - Target international normalised ratio
C1272307|INR - Target international normalized ratio
C1272307|Target international normalized ratio
C2584422|International normalized ratio result obtained using portable international normalized ratio monitoring device (observable entity)
C2584422|International normalized ratio result obtained using portable international normalized ratio monitoring device
C2584422|International normalised ratio result obtained using portable international normalised ratio monitoring device
C1254541|Calculation of international normalised ratio (INR)
C1254541|Calculation of international normalized ratio (INR)
C1254541|Calculation of international normalised ratio
C1254541|Calculation of international normalized ratio
C1254541|Calculation of international normalized ratio (procedure)
C1254541|International Normalized Ratio (INR) Calculations
C3533142|Days in therapeutic INR range/Days INR result determined
C3533142|days in therapeutic INR range / days INR result determined
C3533142|days in therapeutic INR range / days INR result determined (lab test)
C3533142|coag studies: days in therapeutic inr range / days inr result determined
C3838119|coagulation studies: inr in blood or platelet-poor plasma (lab test)
C3838119|coagulation studies: inr in blood or platelet-poor plasma
