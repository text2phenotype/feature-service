C0001899|Alanine Transaminase
C0201836|Alanine aminotransferase measurement
C2257651|L-alanine:2-oxoglutarate aminotransferase activity
C0051063|pyruvate (glyoxylate) aminotransferase
C0051063|Alanine-glyoxylate aminotransferase
C0051063|Alanine glyoxylate aminotransferase
C0051063|Alanine-glyoxylate aminotransferase (substance)
C0051063|Alanine-glyoxylate transaminase
C0283331|alanine-glyoxylate transaminase 1
C0283331|alanine-glyoxylate aminotransferase 1
C0377018|alanine-glyoxylate aminotransferase 2
C0114117|dimethylarginine pyruvate aminotransferase
C0124788|Kynurenine-glyoxylate aminotransferase
C0124788|Kynurenine-glyoxylate aminotransferase (substance)
C0001899|Alanine 2 Oxoglutarate Aminotransferase
C0001899|Alanine Aminotransferase
C0001899|Aminotransferase, Alanine
C0001899|Aminotransferase, Alanine-2-Oxoglutarate
C0001899|Glutamic Alanine Transaminase
C0001899|Glutamic Pyruvic Transaminase
C0001899|Glutamic-Pyruvic Transaminase
C0001899|Transaminase, Glutamic-Alanine
C0001899|Transaminase, Glutamic-Pyruvic
C0001899|L-Alanine:2-oxoglutarate aminotransferase
C0001899|Alanine Transaminase
C0001899|Transaminase, Alanine
C0001899|Glutamic-Alanine Transaminase
C0001899|Alanine Transaminase [Chemical/Ingredient]
C0001899|Alanine-2-Oxoglutarate Aminotransferase
C0001899|GPT
C0001899|ALAT - Alanine aminotransferase
C0001899|ALT - Alanine aminotransferase
C0001899|Glutamate pyruvate transaminase
C0001899|Alanine aminotransferase (substance)
C1980933|Alanine aminotransferase &#x7C; bld-ser-plas
C2703297|Alanine aminotransferase &#x7C; Pleural fluid
C1980932|Alanine aminotransferase &#x7C; amniotic fluid
C1980938|Alanine aminotransferase.macromolecular &#x7C; Bld-Ser-Plas
C2924675|Alanine glyoxylate aminotransferase &#x7C; Tissue and Smears
C1980935|Alanine Aminotransferase &#x7C; Dialysis fluid
C1980937|Alanine aminotransferase &#x7C; red blood cells
C2703296|Alanine aminotransferase &#x7C; Peritoneal fluid
C1980934|Alanine aminotransferase &#x7C; body fluid
C0376147|SGPT
C0376147|SGPT - Glutamate pyruvate transaminase
C0376147|ALT
C0376147|serum glutamate pyruvate transaminase
C0376147|alanine transferase
C0376147|SGPT (ALT)
C3887708|Glutamate Pyruvate Transaminase 1
C3887708|Glutamic--Alanine Transaminase 1
C3887708|Glutamic-Pyruvate Transaminase
C3887708|GPT 1
C3887708|Glutamic--Pyruvic Transaminase 1
C3887708|Alanine Aminotransferase 1
C3887708|EC 2.6.1.2
C3887708|Alanine Aminotransferase 1, human
C3887708|Alanine Aminotransferase
C3887708|Glutamic-Alanine Transaminase
C3887708|Glutamic-Pyruvic Transaminase
C3887708|GPT
C3887708|AAT1
C3887708|GPT1
C3887708|ALT1
C0201836|Alanine aminotransferase measurement
C0201836|Alanine aminotransferase
C0201836|ALT
C0201836|Transferase; alanine amino (ALT) (SGPT)
C0201836|Test;alanine aminotransferase
C0201836|TRANSFERASE ALANINE AMINO ALT SGPT
C0201836|Measurement of alanine amino transferase (ALT) (SGPT)
C0201836|Measurement of alanine amino transferase
C0201836|Liver enzyme (SGPT), level
C0201836|Alanine amino (alt) (sgpt)
C0201836|SGPT
C0201836|Glutamic-pyruvate transaminase
C0201836|GPT
C0201836|GPT measurement
C0201836|Glutamic pyruvate transaminase measurement
C0201836|SGPT measurement
C0201836|ALT measurement
C0201836|Alanine aminotransferase measurement (procedure)
C0201836|alanine aminotransferase test
C1883008|Serum Alanine Aminotransferase Measurement
C1883008|Serum SGPT Measurement
C1883008|Serum Alanine Transaminase Measurement
C1883008|serum alanine aminotransferase measurement (lab test)
C1883008|ALT (SGPT) level
C0428324|Alanine transaminase level
C0428324|Alanine transaminase level (procedure)
C0428325|ALT/SGPT serum level
C0428325|ALT/SGPT serum level (procedure)
C0523461|ALT measurement, method with pyridoxal-5'-phosphate (procedure)
C0523461|Alanine aminotransferase (ALT) measurement, method with pyridoxal-5'-phosphate
C0523461|Alanine aminotransferase measurement, method with pyridoxal-5'-phosphate (procedure)
C0523461|Alanine aminotransferase (ALT) measurement, method with pyridoxal-5'-phosphate (procedure)
C0523461|Alanine aminotransferase measurement, method with pyridoxal-5'-phosphate
C0523461|ALT measurement, method with pyridoxal-5'-phosphate
C0523462|ALT measurement, method without pyridoxal-5'-phosphate (procedure)
C0523462|Alanine aminotransferase (ALT) measurement, method without pyridoxal-5'-phosphate
C0523462|Alanine aminotransferase measurement, method without pyridoxal-5'-phosphate (procedure)
C0523462|Alanine aminotransferase measurement, method without pyridoxal-5'-phosphate
C0523462|Alanine aminotransferase (ALT) measurement, method without pyridoxal-5'-phosphate (procedure)
C0523462|ALT measurement, method without pyridoxal-5'-phosphate
C0428326|Serum glutamic oxaloacetic transaminase (SGPT) - blood measurement (procedure)
C0428326|Serum glutamic oxaloacetic transaminase (SGPT) - blood measurement
C0428326|SGPT - blood measurement (procedure)
C0428326|SGPT - blood level
C0428326|SGPT - blood measurement
C0428327|ALT - blood measurement (procedure)
C0428327|Alanine aminotransferase (ALT) - blood measurement
C0428327|Liver enzymes (& blood level [ALT] or [SGPT])
C0428327|Liver enzymes (& blood level [ALT] or [SGPT]) (procedure)
C0428327|SGPT - blood level
C0428327|ALT - blood level
C0428327|Alanine aminotransferase - blood measurement
C0428327|Alanine aminotransferase (ALT) - blood measurement (procedure)
C0428327|Alanine aminotransferase - blood measurement (procedure)
C0428327|ALT - blood measurement
C0428327|ALT blood measurement
