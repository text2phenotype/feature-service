C0086409|Hispanics
C3846650|Spanish,NOS; Hispanic,NOS
C0019576|Hispanic Americans
C1533017|Hispanic black finding
C1533018|Hispanic black racial group
C1533020|Hispanic white finding
C1533021|Hispanic white racial group
C1881927|Multiple Hispanic
C2741637|Hispanic or Latino:Finding:Point in time:^Patient:Ordina
C3844642|Other Hispanic
C4036190|Yes, another Hispanic, Latino-a, or Spanish origin
C0086409|Hispanic
C0086409|Central American
C0086409|Canal Zone
C0086409|Central American Indian
C0086409|Costa Rican
C0086409|Guatemalan
C0086409|Honduran
C0086409|Nicaraguan
C0086409|Panamanian
C0086409|Salvadoran
C0086409|Cuban
C0086409|Dominican
C0086409|Latin American
C0086409|Mexican
C0086409|Chicano
C0086409|La Raza
C0086409|Mexican American Indian
C0086409|Mexican American
C0086409|Mexicano
C0086409|Puerto Rican
C0086409|South American
C0086409|Argentinean
C0086409|Bolivian
C0086409|Chilean
C0086409|Colombian
C0086409|Criollo
C0086409|Ecuadorian
C0086409|Paraguayan
C0086409|Peruvian
C0086409|South American Indian
C0086409|Uruguayan
C0086409|Venezuelan
C0086409|Spaniard
C0086409|Andalusian
C0086409|Asturian
C0086409|Belearic Islander
C0086409|Canarian
C0086409|Castillian
C0086409|Catalonian
C0086409|Gallego
C0086409|Spanish Basque
C0086409|Valencian
C0019576|American, Hispanic
C0019576|Americans, Hispanic
C0019576|Americans, Spanish
C0019576|Hispanic American
C0019576|Hispanic Americans
C0019576|Spanish American
C0019576|Spanish Americans
C1553379|Cuban
C1553379|-- Cuban
C3829110|Mexican or Mexican American
C3828691|Other Hispanic or Latino(a)
C3161473|Spanish
C3161473|Spanish Person
C0086409|Hispanic
C0086409|Hispanics
C0086409|Hispanic or Latino
C0086409|EthnicityHispanic
C0086409|Hispanic origin
C0086409|Spanish
C0086409|Hispanic Populations
C0086409|Hispanics or Latinos
C0086409|Latino Population
C0086409|Spanish Origin
C0086409|Hispanic (racial group)
C0025884|American, Mexican
C0025884|Americans, Mexican
C0025884|Chicano
C0025884|Mexican American
C0025884|Mexican Americans
C0025884|Chicanos
C0025884|Chicanas
C0025884|Chicana
C0010436|Americans, Cuban
C0010436|Cuban American
C0010436|Cuban Americans
C0086528|Latino
C0086528|Latinos
C0034043|Puerto Rican
C0034043|Puertorican
C0034043|-- Puerto Rican
C0034043|Puerto Ricans
C0935556|Latinos/Latinas
C1533018|Hispanic, black (racial group)
C1533018|Hispanic, black
C1533018|Hispanic black racial group
C1533019|Hispanic, color unknown (racial group)
C1533019|Hispanic, color unknown
C1533019|Hispanic, colour unknown
C1533021|Hispanic, white (racial group)
C1533021|Hispanic, white
C1533021|Hispanic white racial group
C0425359|South American
C0425359|-- South American
C0240339|Mexican
C0240339|EthnicityHispanicMexican
C0240339|-- Mexican
C0238914|Central American
C0238914|EthnicityHispanicCentralAmerican
C0238914|-- Central American
C1328872|Dominican
C1328872|Dominican - Ethnicity
C1553378|Latin American
C0337817|Spaniards
C0337817|Spaniards (ethnic group)
C0337817|Spaniard
C1881927|Multiple Hispanic
C1880193|Cuban or Cuban American
C2135343|cultural background Hispanic (history)
C2135343|the cultural background is Hispanic
C2135343|cultural background Hispanic
C2741637|Hispanic or Latino:Finding:Point in time:^Patient:Ordinal
C2741637|Hispanic or Latino
C2741637|Hispanic or Latino:Find:Pt:^Patient:Ord
