C0035078|Kidney Failure
C1565489|Renal Insufficiency
C0022660|Kidney Failure, Acute
C0022660|Acute renal failure
C0022660|Acute renal failure, unspecified
C0022660|ARF
C0022660|acute renal failure (diagnosis)
C0022660|ARF (acute renal failure)
C0022660|Acute kidney failure
C0022660|Acute kidney failure NOS
C0022660|Acute kidney failure, unspecified
C0022660|Acute and unspecified renal failure
C0022660|Renal Failure, Acute
C0022660|Kidney Failure, Acute [Disease/Finding]
C0022660|Kidney Failures, Acute
C0022660|Acute Kidney Failures
C0022660|Acute Renal Failures
C0022660|Renal Failures, Acute
C0022660|Failure;renal;acute
C0022660|Acute renal failure NOS (disorder)
C0022660|Acute renal failure (disorder)
C0022660|Acute renal failure NOS
C0022660|AKI
C0022660|Acute kidney injury
C0022660|Failure kidney acute
C0022660|Kidney failure acute
C0022660|Renal shutdown acute
C0022660|Renal failure acute
C0022660|Acute renal failure syndrome
C0022660|ARF - Acute renal failure
C0022660|Acute renal failure syndrome (disorder)
C0022660|Acute renal failure syndrome, NOS
C0022661|Kidney Failure, Chronic
C0022661|Chronic renal failure
C0022661|Disease, End-Stage Kidney
C0022661|Disease, End-Stage Renal
C0022661|End-Stage Renal Failure
C0022661|Kidney Disease, End-Stage
C0022661|Renal Disease, End Stage
C0022661|Renal Failure, End Stage
C0022661|End Stage Kidney Disease
C0022661|End Stage Renal Disease
C0022661|CRF
C0022661|Chronic renal failure, unspecified
C0022661|End-stage renal disease
C0022661|End stage chronic renal failure
C0022661|End stage chronc renal failure
C0022661|END STAGE KIDNEY DIS
C0022661|RENAL DIS END STAGE
C0022661|END STAGE RENAL DIS
C0022661|end stage renal failure
C0022661|end stage renal disease (diagnosis)
C0022661|chronic renal failure (diagnosis)
C0022661|ESRD (end stage renal disease)
C0022661|CRF - Chronic Renal Failure
C0022661|Chronic renal disease
C0022661|Chronic renal failure NOS
C0022661|End-Stage Kidney Disease
C0022661|Renal Failure, Chronic
C0022661|ESRD
C0022661|Renal Failure, End-Stage
C0022661|Chronic Kidney Failure
C0022661|Kidney Failure, Chronic [Disease/Finding]
C0022661|Renal Disease, End-Stage
C0022661|Failure;renal;chronic
C0022661|Renal failure - chronic
C0022661|Renal failure (chronic)
C0022661|End stage renal failure (disorder)
C0022661|Failure, renal -chronic
C0022661|Chronic renal failure syndrome
C0022661|Kidney failure chronic
C0022661|End stage renal disease (ESRD)
C0022661|Renal failure chronic
C0022661|ESCRF - End stage chronic renal failure
C0022661|ESRD - End stage renal disease
C0022661|ESRF - End stage renal failure
C0022661|Chronic renal failure syndrome (disorder)
C0022661|End stage renal disease (disorder)
C0022661|disease (or disorder); kidney, end-stage
C0022661|disease (or disorder); renal, end-stage
C0022661|Chronic renal failure syndrome, NOS
C0026766|Failure, Multiple Organ
C0026766|Multiple Organ Failure
C0026766|Multiple Organ Failures
C0026766|multiple organ system failure
C0026766|MOF syndrome
C0026766|Multi-organ failure
C0026766|MOF
C0026766|Multiple System Failure
C0026766|Organ Failure, Multiple
C0026766|Multiple Organ Dysfunction Syndrome
C0026766|Organ Dysfunction Syndrome, Multiple
C0026766|Multiple Organ Failure [Disease/Finding]
C0026766|MODS
C0026766|Multiple organ failure (disorder)
C0026766|Multiorgan failure
C0026766|Multi organ failure
C0026766|multiple organ failure (diagnosis)
C0026766|MODS - Multiple organ dysfunction syndrome
C0026766|MOF - Multiple organ failure
C0026766|MOSF - Multiple organ systems failure
C0026766|MSOF - Multiple systems organ failure
C0026766|Multiple organ systems failure
C0026766|Multiple systems organ failure
C0026766|Multisystem organ failure
C0026766|Multiple organ dysfunction syndrome (disorder)
C0026766|Multiple organ failure, NOS
C0041948|Uremia
C0041948|Uremias
C0041948|UREMIA OF RENAL ORIGIN
C0041948|Uraemia
C0041948|uremia (diagnosis)
C0041948|Uremia [Disease/Finding]
C0041948|Uremia NOS
C0041948|Uraemia NOS
C0041948|Uraemia of renal origin
C0041948|Uremia (disorder)
C0041948|urea in blood; high
C0041948|Uremia, NOS
C0041948|Uraemia, NOS
C0242528|Azotemia
C0242528|Azotaemia
C0242528|Azotemia (disorder)
C0242528|Azotemia [Disease/Finding]
C0242528|Azotemia (finding)
C0035078|KIDNEY FAILURE
C0035078|Renal failure
C0035078|Unspecified renal failure
C0035078|renal failure (diagnosis)
C0035078|Renal failure NOS
C0035078|Unspecified kidney failure
C0035078|Kidney Failure [Disease/Finding]
C0035078|Kidney Failures
C0035078|Failure, Renal
C0035078|Failure, Kidney
C0035078|Failures, Kidney
C0035078|Failures, Renal
C0035078|Renal Failures
C0035078|Renal insufficiency
C0035078|ESRD
C0035078|Renal failure unspecified
C0035078|Renal failure unspecified (disorder)
C0035078|Renal failure (disorder)
C0035078|Renal Failure Syndrome
C0035078|Failure kidney
C0035078|Renal failure, unspecified
C0035078|Renal insufficiency syndrome
C0035078|RF - Renal failure
C0035078|Renal failure syndrome (disorder)
C0035078|failure; renal
C0035078|kidney; failure
C0035078|renal; failure
C0035078|Renal failure syndrome, NOS
C0035078|Renal insufficiency syndrome, NOS
C0035078|renal failure not otherwise specified
C0035078|Failure;renal;NOS
C0403462|Acute on chronic renal failure
C0403462|Renal failure acute on chronic
C0403462|Acute-on-chronic renal failure (disorder)
C0403462|Acute-on-chronic renal failure
C2919930|Uraemia due to inadequate renal perfusion
C2919930|Uremia due to inadequate renal perfusion (disorder)
C2919930|Uremia due to inadequate renal perfusion
C0574786|Acute renal failure with medullary necrosis
C0574786|Acute kidney failure with medullary necrosis
C0574786|Acute renal failure with lesion of renal medullary (papillary) necrosis
C0574786|Acute renal papillary necrosis with renal failure
C0574786|Acute renal papillary necrosis with renal failure (disorder)
C0574786|insufficiency; renal, acute, with necrosis, medullary, medullary
C0574786|kidney; insufficiency, acute, with necrosis, medullary, medullary
C0574786|Acute Renal Failure with Renal Papillary Necrosis
C0574786|Acute renal failure with lesion of renal medullary necrosis
C0495124|Postprocedural renal failure
C0495124|postprocedural renal insufficiency (diagnosis)
C0495124|postprocedural renal insufficiency
C0495124|postprocedural renal failure (diagnosis)
C0495124|insufficiency; renal, postprocedural
C0495124|kidney; insufficiency, postprocedural
C0495124|necrosis; tubular, postprocedural
C0495124|tubular; necrosis, postprocedural
C0410932|Congenital renal failure
C0410932|renal failure congenital
C0410932|Congenital renal failure (diagnosis)
C0410932|Congenital renal failure (disorder)
C0410932|insufficiency; renal, congenital
C0410932|kidney; insufficiency, congenital
C2316810|ESRD
C2316810|End Stage Kidney Disease
C2316810|End Stage Kidney Failure
C2316810|End Stage Renal Failure
C2316810|chronic kidney disease stage 5 (diagnosis)
C2316810|chronic kidney disease stage 5
C2316810|Chronic kidney disease stage 5 (disorder)
C2316810|chronic kidney disease, stage 5
C2316810|End Stage Renal Disease
C2316810|CKD stage 5
C2316810|End-stage renal disease
C2316810|Renal failure, endstage
C2316810|ESRD, End Stage Renal Disease
C2316810|Renal Disease (ESRD), End Stage
C2316810|Renal Disease, End Stage
C2316810|End Stage Renal Disease (ESRD)
C2316810|Disease (ESRD), End Stage Renal
C2316810|Chronic renal failure
C2316810|Stage 5 chronic kidney disease
C2316810|End-stage renal failure
C0404974|Renal shutdown following abortive pregnancy (disorder)
C0404974|Renal shutdown following abortive pregnancy
C1534552|(Renal failure NOS) or (uraemia NOS)
C1534552|(Renal failure NOS) or (uremia NOS)
C1534552|(Renal failure NOS) or (uraemia NOS) (disorder)
C1534552|(Renal failure unspecified) or (uraemia NOS) (disorder)
C1534552|(Renal failure unspecified) or (uraemia NOS)
C1534552|(Renal failure unspecified) or (uremia NOS)
C3662191|Induced termination of pregnancy complicated by renal failure
C3662191|Induced termination of pregnancy complicated by renal failure (disorder)
C3662191|Termination of pregnancy complicated by renal failure
C1565662|acute renal insufficiency (diagnosis)
C1565662|acute renal insufficiency
C1565662|Renal insufficiency (acute)
C1565662|Acute Renal Insufficiencies
C1565662|Renal Insufficiencies, Acute
C1565662|Kidney Insufficiencies, Acute
C1565662|Acute Kidney Insufficiencies
C1565662|Acute Kidney Insufficiency
C1565662|Renal Insufficiency, Acute
C1565662|Kidney Insufficiency, Acute
C1565662|Acute renal impairment
C1565662|Acute renal impairment (disorder)
C1565662|insufficiency; renal, acute
C0588179|Anaemia secondary to renal failure
C0588179|Anemia secondary to renal failure
C0588179|Anaemia secondary to renal failure (disorder)
C0588179|Anemia secondary to renal failure (disorder)
C1565489|Renal insufficiency
C1565489|Impaired renal function
C1565489|renal insufficiency (diagnosis)
C1565489|Renal Insufficiency [Disease/Finding]
C1565489|Kidney Insufficiency
C1565489|Insufficiency;renal
C1565489|Renal impairment (disorder)
C1565489|Renal impairment
C1565489|Renal dysfunction
C1565489|Kidney Impairment
C1565489|Insufficiency renal
C1565489|Renal impairment NOS
C1565489|insufficiency; renal
C1565489|kidney; insufficiency
C1565489|Kidney Insufficiencies
C1565489|Renal Insufficiencies
C1565489|Insufficiency, Kidney
C4075836|Renal failure syndrome co-occurrent with human immunodeficiency virus infection
C4075836|Renal failure syndrome co-occurrent with human immunodeficiency virus infection (disorder)
C0026141|Milk Alkali Syndrome
C0026141|Syndrome, Milk-Alkali
C0026141|Milk-alkali syndrome
C0026141|milk alkali syndrome (diagnosis)
C0026141|Burnett syndrome
C0026141|Burnett's syndrome
C0026141|Milk alkali syndrome (disorder)
C0026141|Burnett
C0026141|milk-alkali; syndrome
C0026141|syndrome; milk-alkali
C0348879|Hypertensive heart and renal disease, unspecified, with renal failure
C0348879|Hypertensive heart and renal disease with renal failure
C0348879|hypertensive heart and renal disease with renal failure (diagnosis)
C0348879|hypertensive heart and chronic kidney disease with renal failure
C0348879|Hy ht/kd NOS st V w/o hf
C0348879|Hypertensive heart and chronic kidney disease, unspecified, without heart failure and with chronic kidney disease stage V or end stage renal disease
C0348879|Hypertensive heart and renal disease with renal failure (disorder)
C0348879|failure; cardiorenal, hypertensive, with renal failure
C0348879|insufficiency; renal, with hypertensive heart disease
C0348879|kidney; insufficiency, with hypertensive heart disease
C0348860|Hypertensive renal disease, unspecified, with renal failure
C0348860|Hypertensive renal disease with renal failure
C0348860|Hyp kid NOS w cr kid V
C0348860|Hypertensive chronic kidney disease, unspecified, with chronic kidney disease stage V or end stage renal disease
C0348860|hypertensive kidney disease with renal failure (diagnosis)
C0348860|hypertensive kidney disease with renal failure
C0348860|Hypertensive renal disease with renal failure (disorder)
C0348860|hypertension; renal disease, hypertensive, with renal failure
C0348860|insufficiency; renal, chronic, hypertensive
C0348860|insufficiency; renal, with hypertension
C0348860|kidney; hypertension, with renal failure
C0494576|Hypertensive heart and renal disease, unspecified, with congestive heart failure and renal failure
C0494576|Hypertensive heart and renal disease with both (congestive) heart failure and renal failure
C0494576|Hyp ht/kd NOS st V w hf
C0494576|Hypertensive heart and chronic kidney disease, unspecified, with heart failure and chronic kidney disease stage V or end stage renal disease
C0494576|Hypertensive heart and renal disease, unspecified, with heart failure and renal failure
C0494576|Hypertensive heart and renal disease with both (congestive) heart failure and renal failure (disorder)
C0494576|insufficiency; renal, with hypertensive heart disease and heart failure
C0494576|kidney; insufficiency, with hypertensive heart disease and heart failure
C0403448|Kidney failure as a complication of care
C0403448|Renal failure as a complication of care
C0403448|Renal failure as a complication of care (disorder)
C0404973|renal failure following abortion
C0404973|renal failure following abortion (diagnosis)
C0404973|Renal failure NOS following abortive pregnancy
C0404973|Renal failure following abortive pregnancy
C0404973|Renal failure NOS following abortive pregnancy (finding)
C0404973|Renal failure NOS following abortive pregnancy (disorder)
C0404973|Renal failure following abortive pregnancy (disorder)
C0477745|Other acute renal failure
C0477745|Other acute kidney failure
C0477745|[X]Other acute renal failure
C0477745|Other acute renal failure (disorder)
C0477745|[X]Other acute renal failure (disorder)
C0477746|Other chronic renal failure
C0477746|[X]Other chronic renal failure
C0477746|[X]Other chronic renal failure (disorder)
C0542211|Postoperative renal failure
C0542211|Postoperative renal failure (disorder)
C0156556|Unspecified abortion complicated by renal failure
C0156556|Unspecified type of abortion, unspecified, complicated by renal failure
C0156556|abortion complicated by renal failure (diagnosis)
C0156556|abortion complicated by renal failure
C0156556|abortion with renal failure
C0156556|Ab NOS w renal fail-unsp
C0156556|Unspecified abortion, complicated by renal failure, unspecified
C0156556|Abortion complicated by renal failure (disorder)
C2931783|ERS
C2931783|AI1G
C2931783|AMELOGENESIS IMPERFECTA, TYPE IG
C2931783|Amelogenesis imperfecta nephrocalcinosis
C2931783|Enamel renal syndrome
C2931783|Generalized enamel hypoplasia and renal dysfunction
C2931783|Absent enamel, nephrocalcinosis and apparently normal calcium metabolism
C2931783|Amelogenesis Imperfecta, Hypoplastic, and Nephrocalcinosis
C2931783|Enamel-Renal Syndrome
C2931783|AMELOGENESIS IMPERFECTA AND GINGIVAL FIBROMATOSIS SYNDROME
C2931783|AIGFS
C2931783|AMELOGENESIS IMPERFECTA, HYPOPLASTIC, WITH NEPHROCALCINOSIS
C2931783|ENAMEL-RENAL-GINGIVAL SYNDROME
C2931783|Amelogenesis imperfecta and nephrocalcinosis
C2931783|McGibbon Lubinsky syndrome
C2931783|Enamel-renal syndrome (disorder)
C2931783|Lubinsky syndrome
C2931783|Amelogenesis imperfecta, nephrocalcinosis and impaired renal concentration
C0269314|Renal failure following molar AND/OR ectopic pregnancy (disorder)
C0269314|Renal failure following molar AND/OR ectopic pregnancy
C0269314|Renal failure following molar or ectopic pregnancy
C1386521|uremic; aphasia
C1386521|aphasia; uremic
C1390022|blindness; uremic
C1390022|uremic; blindness
C0151567|Coma uraemic
C0151567|Uraemic coma
C0151567|Coma uremic
C0151567|Uremic coma
C0151567|Uremic coma (disorder)
C0151567|coma; uremic
C0151567|uremic; coma
C0234540|Uremic convulsion
C0234540|Uraemic convulsion
C0234540|Uremic convulsion (finding)
C0234540|convulsions; uremic
C0234540|uremic; convulsions
C0748288|decompensation; renal
C0748288|kidney; decompensation
C1395122|delirium; uremic
C1395122|uremic; delirium
C1395967|dyspnea; uremic
C1395967|uremic; dyspnea
C0232807|Decreased renal function
C0232807|Decreased kidney function
C0232807|Function kidney decreased
C0232807|Decreased renal function (finding)
C0232807|function; low, kidney
C0232807|low; function, kidney
C0151746|Abnormal renal function
C0151746|Renal functional abnormality
C0151746|Abnormal renal physiology
C0151746|Abnormality of renal physiology
C0151746|Dysfunction kidney
C0151746|Renal function abnormal
C0151746|Function kidney abnormal
C0151746|Kidney dysfunction
C0151746|Kidney function abnormal
C0151746|Abnormal renal function (finding)
C0151746|dysfunction; kidney
C1401758|fever; uremic
C1401758|uremic; fever
C1408265|kidney; functional disturbance
C0232808|nonfunctioning kidney (diagnosis)
C0232808|nonfunctioning kidney
C0232808|Non-functioning kidney
C0232808|Non-functioning kidney (disorder)
C0232808|NFK - Non-functioning kidney
C0232808|Shutdown renal
C0232808|Absent renal function
C0232808|kidney; nonfunctioning
C0232808|nonfunctioning; kidney
C0232808|Absent renal function (disorder)
C0232808|Absent renal function (finding)
C1407023|kidney; toxemia
C1407023|toxemia; kidney
C1406177|renal; suppression
C1406177|suppression; renal
C1407025|toxemia; uremic
C1407025|uremic; toxemia
C1407026|toxemia; urinary
C1407026|urinary; toxemia
C0235446|Azotemia due to intrarenal disease
C0235446|Renal azotemia
C0235446|Renal azotemia (disorder)
C0235446|Intrarenal azotemia
C0235446|Azotaemia due to intrarenal disease
C0235446|Azotemia due to intrarenal disease (disorder)
C0235446|Intrarenal azotaemia
C0235446|Renal azotaemia
C0235446|Azotemia renal
C0235446|Azotaemia renal
C0235446|Azotemia of renal origin
C0235446|Azotaemia of renal origin
C1278220|Deteriorating renal function
C1278220|Deteriorating renal function (finding)
C1278220|Deteriorating renal function (situation)
C0456040|Newborn renal dysfunction
C0456040|Newborn renal dysfunction (disorder)
C0403447|chronic renal insufficiency
C0403447|chronic renal insufficiency (diagnosis)
C0403447|Chronic Kidney Insufficiency
C0403447|Renal Insufficiency, Chronic
C0403447|Renal Insufficiency, Chronic [Disease/Finding]
C0403447|Kidney Insufficiency, Chronic
C0403447|Chronic renal impairment
C0403447|Chronic renal impairment (disorder)
C0403447|insufficiency; renal, chronic, end stage renal disease
C0403447|insufficiency; renal, chronic
C0403447|insufficiency; renal, end stage
C0403447|kidney; insufficiency, chronic
C0403447|Chronic Kidney Insufficiencies
C0403447|Chronic Renal Insufficiencies
C0403447|Kidney Insufficiencies, Chronic
C0403447|Renal Insufficiencies, Chronic
C0585398|Acute-on-chronic renal impairment (disorder)
C0585398|Acute-on-chronic renal impairment
C2242703|Cardiorenal syndrome
C2242703|Cardiorenal syndrome (disorder)
C2242703|Cardio-Renal Syndromes
C2242703|Syndrome, Renocardiac
C2242703|Syndrome, Cardiorenal
C2242703|Cardio-Renal Syndrome
C2242703|Syndrome, Cardio-Renal
C2242703|Syndromes, Cardio-Renal
C2242703|Cardiorenal Syndromes
C2242703|Syndromes, Cardiorenal
C2242703|Reno-Cardiac Syndromes
C2242703|Syndromes, Renocardiac
C2242703|Cardio Renal Syndrome
C2242703|Renocardiac Syndromes
C2242703|Reno Cardiac Syndrome
C2242703|Syndrome, Reno-Cardiac
C2242703|Syndromes, Reno-Cardiac
C2242703|Reno-Cardiac Syndrome
C2242703|Cardio-Renal Syndrome [Disease/Finding]
C2242703|Renocardiac Syndrome
C1859722|ARC syndrome
C1859722|Arthrogryposis renal dysfunction cholestasis syndrome
C1859722|Arthrogryposis multiplex congenita, renal dysfunction, and cholestasis
C1859722|ARCS1
C1859722|ARCS
C1859722|ARTHROGRYPOSIS, RENAL DYSFUNCTION, AND CHOLESTASIS 1
C1859722|Arthrogryposis, Renal Dysfunction, And Cholestasis
C1852759|PAPILLORENAL SYNDROME
C1852759|Optic nerve coloboma with renal disease
C1852759|Coloboma of optic nerve with renal disease
C1852759|Renal-coloboma syndrome
C1852759|Optic coloboma, vesicoureteral reflux, and renal anomalies
C1852759|Renal coloboma syndrome (disorder)
C1852759|Renal coloboma syndrome
C1852759|Renal-Coloboma Syndrome With Macular Abnormalities
C1852759|Optic Nerve Coloboma Renal Syndrome
C1852759|Coloboma-Ureteral-Renal Syndrome
C1852759|PAPRS
C1852759|CONGENITAL ANOMALIES OF THE KIDNEY AND URINARY TRACT WITH OR WITHOUT OCULAR ABNORMALITIES
C1852759|CAKUT WITH OR WITHOUT OCULAR ABNORMALITIES
C0400972|BILIARY MALFORMATION WITH RENAL TUBULAR INSUFFICIENCY
C0400972|Cholestatic jaundice and renal tubular insufficiency
C0400972|Lutz Richner Landolt syndrome
C0400972|Renal tubular insufficiency, cholestatic jaundice, and multiple congenital anomalies
C0400972|Biliary malformation associated with renal tubular insufficiency
C0400972|Biliary malformation associated with renal tubular insufficiency (disorder)
C2609414|Acute Kidney Injury
C2609414|Acute Renal Injuries
C2609414|Renal Injury, Acute
C2609414|Acute Kidney Injuries
C2609414|Renal Injuries, Acute
C2609414|Kidney Injury, Acute
C2609414|Kidney Injuries, Acute
C2609414|Acute Kidney Injury [Disease/Finding]
C2609414|Acute Renal Injury
C2609414|Acute injury of kidney
C2609414|Acute injury of kidney (disorder)
C0403361|renal insufficiency with growth failure
C0403361|renal insufficiency with growth failure (diagnosis)
C0403361|Renal function impairment with growth failure
C0403361|Renal function impairment with growth failure (disorder)
C0403720|NEPHROLITHIASIS, X-LINKED RECESSIVE, WITH RENAL FAILURE
C0403720|XRN
C0403720|NPHL1
C0403720|X-linked recessive nephrolithiasis with renal failure
C0403720|Nephrolithiasis 1
C0403720|Nephrolithiasis, X-Linked Recessive, Type 1
C0403720|Urolithiasis, X-Linked Recessive, Type 1
C0403720|X-linked recessive nephrolithiasis with renal failure (disorder)
C2751310|HNFJ2
C2751310|HYPERURICEMIC NEPHROPATHY, FAMILIAL JUVENILE, 2
C2751310|Early-Onset Hyperuricemia, Anemia, And Progressive Kidney Failure
C2751310|Hyperuricemic Nephropathy, Familial Juvenile 2
C2751310|Familial Juvenile Hyperuricemic Nephropathy 2
C2751310|Ren-Related Kidney Disease
C3854173|Pre-renal acute kidney injury (disorder)
C3854173|Prerenal renal failure
C3854173|Acute renal failure
C3854173|Pre-renal acute kidney injury
C1839604|Renal failure in adulthood
C1561643|Chronic renal disease
C1561643|Chronic Kidney Disease
C1561643|Chronic kidney dis NOS
C1561643|CKD - Chronic Kidney Disease
C1561643|Chronic kidney disease (CKD)
C1561643|Chronic kidney disease, unspecified
C1561643|Disease, Chronic Kidney
C1561643|Diseases, Chronic Renal
C1561643|Kidney Diseases, Chronic
C1561643|Disease, Chronic Renal
C1561643|Diseases, Chronic Kidney
C1561643|Renal Disease, Chronic
C1561643|Kidney Disease, Chronic
C1561643|Renal Diseases, Chronic
C1561643|CKD
C1561643|Chronic Kidney Diseases
C1561643|Chronic Renal Insufficiency
C1561643|Loss of renal function
C1561643|Chronic kidney disease (disorder)
C1561643|Chronic Renal Failure
C1561643|Chronic Renal Diseases
C1561643|disease (or disorder); kidney, chronic
C1561643|kidney; disease, chronic
C1843276|Renal failure, reversible
C1843276|Reversible renal failure
C0184571|Impaired Kidney Function
C0184571|rndx renal alteration
C0184571|rndx renal alteration (diagnosis)
C0184571|Renal Alteration
C0184571|Renal alteration (finding)
C0184571|change; renal
C0184571|kidney; change
C4076161|Renal impairment caused by Polyomavirus (disorder)
C4076161|Renal impairment caused by Polyomavirus
C1285418|Renal failure associated with renal vascular disease (disorder)
C1285418|Renal failure associated with renal vascular disease
