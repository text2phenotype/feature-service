C0200665|Mean platelet volume
C0032181|Blood Platelet Counts
C0005821|Blood Platelets
C0920267|Platelet aggregation measurement
C0200642|Platelet estimate
C0200665|Mean platelet volume
C0200665|mean platelet volume (MPV) (lab test)
C0200665|mean platelet volume (MPV)
C0200665|MPV
C0200665|Mean Platelet Volume Measurement
C0200665|Volumes, Mean Platelet
C0200665|Platelet Volumes, Mean
C0200665|Platelet Volume, Mean
C0200665|Volume, Mean Platelet
C0200665|Mean Platelet Volumes
C0200665|MPV - Mean platelet volume
C0200665|Platelet mean volume (observable entity)
C0200665|Platelet mean volume
C0200665|Platelet mean volume determination
C0200665|Platelet mean volume determination (procedure)
C0344388|Platelet mean volume
C0344388|Mean platelet volume (procedure)
C0344388|Mean platelet volume (observable entity)
C0344388|Mean platelet volume
C0344388|Platelet mean volume finding
C1254925|Operating Room Misc Labs: Platelets
C0032181|Blood Platelet Counts
C0032181|Blood Platelet Numbers
C0032181|Count, Blood Platelet
C0032181|Count, Platelet
C0032181|Counts, Blood Platelet
C0032181|Counts, Platelet
C0032181|Number, Blood Platelet
C0032181|Number, Platelet
C0032181|Numbers, Blood Platelet
C0032181|Numbers, Platelet
C0032181|Platelet Count
C0032181|Platelet Count, Blood
C0032181|Platelet Counts
C0032181|Platelet Counts, Blood
C0032181|Platelet Number, Blood
C0032181|Platelet Numbers
C0032181|Platelet Numbers, Blood
C0032181|platelets
C0032181|platelet count (lab test)
C0032181|Platelet count NOS (procedure)
C0032181|Platelet count NOS
C0032181|Platelet count (procedure)
C0032181|PLAT
C0032181|Anucleated Thrombocytes
C0032181|Thrombocyte count
C0032181|Platelet Number
C0032181|Blood Platelet Count
C0032181|Blood Platelet Number
C0032181|Whole Blood Platelet Counts
C0032181|Plt - Platelet count
C0032181|Platelet count - observation
C0032181|Platelet Count measurement
C2697501|Giant Platelet Count
C2697501|Giant Platelet Count (procedure)
C2697501|Giant Platelets
C2697501|PLATGNT
C2697898|Large Platelet Count
C2697898|PLATLRG
C2697898|Large Platelets
C1314099|reticulated platelet assay (lab test)
C1314099|reticulated platelet assay
C1314099|Reticulated (young) platelet measurement
C1314099|Assay for reticulated platelets
C2082381|plasma platelet count
C2082381|plasma platelet count (lab test)
C2702985|immature platelet fraction (lab test)
C2702985|immature platelet fraction
C0523117|manual platelet count (lab test)
C0523117|manual platelet count
C0523117|Platelet count, blood, manual
C0523117|Platelet count, blood, manual (procedure)
C2082406|platelet count estimation from smear (lab test)
C2082406|platelet count estimation from smear
C2082406|platelet estimation from smear
C1144713|automated platelet count
C1144713|automated platelet count (lab test)
C1144713|BLOOD COUNT PLATELET AUTOMATED
C1144713|Platelet count, automated test
C1144713|Blood count; platelet, automated
C3272909|Platelet Clumps Count
C3272909|Platelet Clumps
C3272909|PLT Clumps
C3272909|PLATCLMP
C0523118|Platelet count, blood, automated
C0523118|Platelet count, blood, automated (procedure)
C1294068|Platelet count, Rees-Ecker method (procedure)
C1294068|Platelet count, Rees-Ecker method
C1443989|Serial platelet counts (procedure)
C1443989|Serial platelet counts
C0005821|Thrombocyte
C0005821|Blood Platelets
C0005821|Platelet
C0005821|Platelet, Blood
C0005821|Platelets, Blood
C0005821|Blood Platelet
C0005821|Platelets
C0005821|Platelet (cell structure)
C0005821|PLT - Platelet
C0005821|PLT - Platelets
C0005821|Platelet (body structure)
C0005821|Thrombocyte (platelet)
C0005821|Deetjen Body
C0005821|Bizzozero Corpuscle
C0005821|Thrombocytes
C0005821|Platelet [dup] (body structure)
C0005821|Platelets (Blood)
C0005821|Reticuloendothelial System, Platelets
C2751259|MACROTHROMBOCYTOPENIA, AUTOSOMAL DOMINANT, TUBB1-RELATED
C0427568|Platelet satellite
C0427568|Platelet satellite (cell structure)
C0427568|Platelet satellite (body structure)
C0427566|Macrothrombocytes
C0427566|Macrothrombocyte
C0427566|Macrothrombocyte (cell structure)
C0427566|Macrothrombocyte (body structure)
C0427567|Microthrombocyte
C0427567|Microthrombocyte (cell structure)
C0427567|Microthrombocyte (body structure)
C0484484|Platelets given:Type:Pt:^Patient:Nom
C0484484|Platelets given [Type]
C0484484|Platelet Gvn
C0484484|Platelets given:Type:Point in time:^Patient:Nominal
C2966248|Platelets &#x7C; Fetus &#x7C; Bld-Ser-Plas
C2964883|Bizarre platelets &#x7C; Bld-Ser-Plas
C1994889|Platelets agranular &#x7C; bld-ser-plas
C1994884|Platelets &#x7C; blood cord
C0363450|Platelets given [Volume]
C0363450|Platelets given:Vol:Pt:Dose:Qn
C0363450|Platelet Gvn Vol Dose
C0363450|Platelets given:Volume:Point in time:Dose med or substance:Quantitative
C2972547|Transfuse platelets &#x7C; patient
C1994885|Platelets &#x7C; body fluid
C1305955|Megakaryocytes
C1305955|Investigation of megakaryocytes
C2966378|Reticulocytes.high light scatter &#x7C; Bld-Ser-Plas
C1994886|Platelets &#x7C; Bone marrow
C1994891|Platelets large &#x7C; bld-ser-plas
C0370058|Platelet Ab
C0370058|Platelet Antibody
C0370058|Anti-platelet antibody
C0370058|Anti-platelet antibody (substance)
C2358582|Platelets reticulated &#x7C; Bld-Ser-Plas
C1979797|Platelet indices
C1994887|Platelets &#124; dialysis fluid
C1994887|Platelets &#x7C; dialysis fluid
C3700279|Platelets &#x7C; Blood capillary
C1994893|Platelets small &#x7C; bld-ser-plas
C1994883|Platelets &#x7C; bld-ser-plas
C3847483|Platelets &#x7C; Platelet rich plasma
C4072392|Giant platelets &#x7C; Bld-Ser-Plas
C4072048|Platelet dense bodies &#x7C; Bld-Ser-Plas
C1512639|Immature Platelet
C0200474|platelet aggregation to adenosine diphosphate (lab test)
C0200474|platelet aggregation to adenosine diphosphate
C0200474|platelet aggregation to ADP
C0200474|Platelet aggregation with adenosine diphosphate test (procedure)
C0200474|Platelet aggregation with adenosine diphosphate test
C0200474|Platelet aggregation with ADP test (procedure)
C0200474|Platelet Adp Aggregation Test
C0200474|Platelet aggregation with ADP test
C0200476|platelet aggregation induced by collagen
C0200476|platelet aggregation induced by collagen (lab test)
C0200476|Platelet Collagen Aggregation Test
C0200476|Platelet aggregation with collagen test
C0200476|Platelet aggregation with collagen test (procedure)
C1255223|Platelet Epinhephrine Aggregation Test
C0522868|Platelet Ristocetin Aggregation Test
C0522868|Platelet aggregation with ristocetin test
C0522868|Platelet aggregation with ristocetin test (procedure)
C0920267|platelet aggregation
C0920267|platelet aggregation (lab test)
C0920267|Platelet aggr
C0920267|Platelet aggregation measurement
C0920267|Platelet aggregation test (procedure)
C0920267|Platelet aggregation assay (qualifier value)
C0920267|Platelet aggregation assay
C0920267|Platelet aggregation test
C0920267|PLATAGGR
C0920267|Platelet Function
C0920267|Platelet aggregation NOS
C0920267|Aggregometer test
C0920267|Platelet aggregation test, NOS
C0920267|Aggregometer test, NOS
C2082403|platelet aggregation induced by bovine factor VIII (lab test)
C2082403|platelet aggregation induced by bovine factor VIII
C0200475|platelet aggregation induced by epinephrine
C0200475|platelet aggregation induced by epinephrine (lab test)
C0200475|Platelet aggregation with epinephrine test
C0200475|Platelet aggregation with adrenaline test
C0200475|Platelet aggregation with epinephrine test (procedure)
C2082404|platelet aggregation induced by ristocetin (lab test)
C2082404|platelet aggregation induced by ristocetin
C0200470|Heparin assay
C0200470|Assay for heparin
C0200470|Heparin assay (procedure)
C0200470|Heparin assay (qualifier value)
C0200470|Heparin assay, NOS
C0200477|Platelet aggregation with thrombin test
C0200477|Platelet aggregation with thrombin test (procedure)
C0200478|Platelet aggregation with drug test
C0200478|Platelet aggregation with drug test (procedure)
C0522869|Platelet aggregation with arachidonate test
C0522869|Platelet aggregation with arachidonate test (procedure)
C0522866|Platelet aggregation with calcium ionophore test
C0522866|Platelet aggregation with calcium ionophore test (procedure)
C0522867|Platelet aggregation with norepinephrine test
C0522867|Platelet aggregation with noradrenaline test
C0522867|Platelet aggregation with norepinephrine test (procedure)
C0522870|Platelet aggregation with serotonin test
C0522870|Platelet aggregation with serotonin test (procedure)
C0427578|Platelet aggregation ratio
C0427578|Platelet aggregation ratio measurement (procedure)
C0427578|Platelet aggregation ratio measurement
C0373809|Platelet, aggregation (in vitro), each agent
C0373809|PLATELET AGGREGATION IN VITRO EACH AGENT
C0373809|BLOOD PLATELET AGGREGATION
