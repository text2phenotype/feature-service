C0004364|Autoimmune Diseases
C0400936|Autoimmune liver disease
C0850560|Other autoimmune disease
C1328839|autoimmune inflammatory bowel disease
C1384868|disease (or disorder); autoimmune (systemic)
C0035012|Reiter's syndrome
C0035012|Reiter's disease
C0035012|Reiters Disease
C0035012|REITER DIS
C0035012|Disease, Reiter's
C0035012|Syndrome, Reiter
C0035012|Disease, Reiter
C0035012|REITERS DIS
C0035012|Fiessinger Leroy Reiter syndrome
C0035012|Reiter's syndrome with arthropathy
C0035012|Reiter's syndrome with arthropathy (diagnosis)
C0035012|Reiter's syndrome (diagnosis)
C0035012|Reiter Syndrome
C0035012|Reiter disease
C0035012|Reiter's disease, unspecified site
C0035012|Reiters syndrome
C0035012|Reiter's disease (disorder)
C0035012|Fiessinger-Leroy-Reiter syndrome
C0035012|Urethrooculoarticular syndrome
C0035012|arthritis; urethritica
C0035012|Reiter; triad
C0035012|Reiter
C0035012|syndrome; urethro-oculo-articular
C0035012|triad; Reiter
C0035012|urethritica; arthritis
C0035012|urethro-oculo-articular; syndrome
C0035012|uroarthritis; infectious
C0001403|Addisons Disease
C0001403|Disease, Addison
C0001403|Addison's disease
C0001403|Primary adrenocortical insufficiency
C0001403|Adrenal insufficiency (Addison disease)
C0001403|Addison disease
C0001403|Primary adrenocortical failure
C0001403|ADDISONS DIS
C0001403|ADDISON DIS
C0001403|Addison's disease NOS
C0001403|primary adrenal insufficiency
C0001403|primary adrenal insufficiency (diagnosis)
C0001403|Addison Disease [Disease/Finding]
C0001403|Primary Hypoadrenalism
C0001403|Disease;Addisons
C0001403|Hypocortisolism
C0001403|Addison's disease, NOS
C0001403|Addison's disease (disorder)
C0001403|Addison's disease, NOS (disorder)
C0001403|Primary adrenal deficiency
C0001403|Chronic Primary Adrenal Insufficiency
C0001403|Disease Addison's
C0001403|Primary adrenocortical insufficiency (disorder)
C0001403|corticoadrenal; deficiency, primary
C0001403|deficiency; adrenocortical, primary
C0001403|deficiency; corticoadrenal, primary
C0001403|disease (or disorder); bronzed skin (Addison) (bronze disease)
C0001403|hypoadrenocorticism; primary
C0001403|insufficiency; adrenal, primary
C0001403|insufficiency; suprarenal, primary
C0001403|adrenal cortex; deficiency, primary
C0001403|adrenal cortex; hypofunction, primary
C0001403|adrenal; insufficiency, primary
C0001403|primary; hypoadrenocorticism
C0001403|Addison; disease or syndrome
C0001403|suprarenal; insufficiency, primary
C0001403|syndrome; Addison
C0001403|Addison's disease [Ambiguous]
C0001403|Hypoadrenalism, Primary
C0001403|Hypoadrenalisms, Primary
C0001403|Insufficiencies, Primary Adrenocortical
C0001403|Insufficiency, Primary Adrenocortical
C0001403|Primary Adrenocortical Insufficiencies
C0001403|Adrenal Insufficiency, Primary
C0001403|Adrenocortical Insufficiencies, Primary
C0001403|Adrenocortical Insufficiency, Primary
C1527336|Sjogren's Syndrome
C1527336|Syndrome, Sjogren's
C1527336|Sjogrens Syndrome
C1527336|Sicca syndrome [Sjogren]
C1527336|Sjogren's disease
C1527336|SJOGREN SYNDROME
C1527336|Sjogren's Syndrome [Disease/Finding]
C1527336|Sicca (Sjogren's) syndrome
C1527336|Sjogren syndrome (diagnosis)
C1527336|Sjogren's
C1527336|Gougerot-Mulock-Houwer syndrome
C1527336|Syndrome Sjogren's
C1527336|Sjoegren's syndrome
C1527336|Sjögren's syndrome (disorder)
C1527336|Sjögren
C0002880|Autoimmune hemolytic anemia
C0002880|Anemia, Hemolytic, Autoimmune
C0002880|Hemolytic anemia, autoimmune
C0002880|ANEMIA, AUTOIMMUNE HEMOLYTIC
C0002880|Autoimmun hemolytic anem
C0002880|Anemia, Hemolytic, Autoimmune [Disease/Finding]
C0002880|Autoimmune haemolytic anaemias
C0002880|AIHA - Autoimmune hemolytic anemia
C0002880|AIHA - Autoimmune haemolytic anaemia
C0002880|Autoimmune haemolytic anaemia (disorder)
C0002880|Autoimmune hemolytic anemia NOS (disorder)
C0002880|Autoimmune haemolytic anaemia
C0002880|Hemolytic anemia due to antibody
C0002880|Autoimmune hemolytic anemia NOS
C0002880|Haemolytic anaemia due to antibody
C0002880|Autoimmune hemolytic anemia (disorder)
C0002880|Autoimmune hemolytic anemias
C0002880|Autoimmune haemolytic anaemia NOS
C0002880|Immune mediated hemolytic anemia
C0002880|Anemia hemolytic autoimmune (NOS)
C0002880|Anaemia haemolytic autoimmune
C0002880|Anemia hemolytic autoimmune
C0002880|hemolytic; anemia, autoimmune
C0002880|anemia; hemolytic, autoimmune
C0002880|Autoimmune hemolytic anemia, NOS
C0002880|Hemolytic anemia due to antibody, NOS
C0002880|Anemias, Autoimmune Hemolytic
C0002880|Hemolytic Anemias, Autoimmune
C0015300|Exophthalmos
C0015300|Proptoses
C0015300|Exophthalmus
C0015300|Exophthalmia
C0015300|Ocular proptosis
C0015300|Proptosis
C0015300|Bulging eyes
C0015300|exophthalmos (diagnosis)
C0015300|eyes bulging out as symptom
C0015300|proptosis (physical finding)
C0015300|eyes bulging out
C0015300|eyes bulging out (symptom)
C0015300|Exophthalmos NOS
C0015300|Unspecified exophthalmos
C0015300|Exophthalmos [Disease/Finding]
C0015300|Eye bulging
C0015300|Prolapsed globe
C0015300|Anterior bulging of the globe
C0015300|Exophthalmos, unspecified
C0015300|Eye displaced forwards
C0015300|Exophthalmos (disorder)
C0015300|Exophthalmos, NOS
C0015300|Proptosis, NOS
C0014072|Encephalomyelitis, Experimental Allergic
C0014072|Experimental Allergic Encephalomyelitides
C0014072|experimental allergic encephalomyelitis
C0014072|ALLERGIC ENCEPH
C0014072|ALLERGIC ENCEPH EXPER
C0014072|EXPER ALLERGIC ENCEPH
C0014072|ENCEPH EXPER AUTOIMMUNE
C0014072|ENCEPH AUTOIMMUNE EXPER
C0014072|AUTOIMMUNE ENCEPH EXPER
C0014072|AUTOIMMUNE EXPER ENCEPH
C0014072|ENCEPH ALLERGIC
C0014072|EXPER AUTOIMMUNE ENCEPH
C0014072|autoimmune encephalomyelitis
C0014072|EAE
C0014072|Encephalomyelitis, Autoimmune Experimental
C0014072|Experimental Encephalomyelitis, Autoimmune
C0014072|Experimental Autoimmune Encephalomyelitis
C0014072|Autoimmune Experimental Encephalomyelitis
C0014072|Encephalomyelitis, Autoimmune, Experimental [Disease/Finding]
C0014072|Autoimmune Encephalomyelitis, Experimental
C0014072|Encephalomyelitis, Experimental Autoimmune
C0014072|Encephalomyelitis, Autoimmune, Experimental
C0014072|Allergic Encephalomyelitis, Experimental
C0014072|Encephalomyelitis, Allergic
C0014072|Allergic Encephalomyelitis
C0014072|Experimental allergic encephalomyelitis (disorder)
C0014072|Allergic encephalomyelitis (disorder)
C0017658|Glomerulonephritides
C0017658|Glomerulonephritis
C0017658|glomerulonephritis (diagnosis)
C0017658|glomerulonephritis NOS
C0017658|Glomerulonephritis [Disease/Finding]
C0017658|Unspecified glomerulonephritis NOS (disorder)
C0017658|Unspecified glomerulonephritis NOS
C0017658|Glomrulonephritis
C0017658|Nephritis-glomerular
C0017658|Glomerular Nephritis
C0017658|GN - Glomerulonephritis
C0017658|Glomerulonephritis (disorder)
C0017658|Glomerulonephritis, NOS
C0020951|Immune Complex Diseases
C0020951|Disease, Immune Complex
C0020951|Diseases, Immune Complex
C0020951|Hypersensitivities, Type III
C0020951|Type III Hypersensitivities
C0020951|Immune Complex Disease
C0020951|IMMUNE COMPLEX DIS
C0020951|Immune Complex Diseases [Disease/Finding]
C0020951|Type III Hypersensitivity
C0020951|Hypersensitivity, Type III
C0011854|Brittle Diabetes Mellitus
C0011854|Diabetes Mellitus, Insulin-Dependent
C0011854|Diabetes Mellitus, Juvenile Onset
C0011854|Diabetes Mellitus, Ketosis Prone
C0011854|IDDM
C0011854|Insulin-Dependent Diabetes Mellitus
C0011854|Juvenile-Onset Diabetes Mellitus
C0011854|Ketosis-Prone Diabetes Mellitus
C0011854|Diabetes Mellitus, Insulin Dependent
C0011854|insulin dependent diabetes mellitus
C0011854|Diabetes Mellitus, Sudden Onset
C0011854|Mellitus, Sudden-Onset Diabetes
C0011854|Sudden-Onset Diabetes Mellitus
C0011854|JOD
C0011854|IDDM1
C0011854|INSULIN-DEPENDENT DIABETES MELLITUS 1
C0011854|Insulin-dependent diabetes mellitus (type I)
C0011854|DIABETES MELLITUS, INSULIN-DEPENDENT, 1
C0011854|DIABETES MELLITUS TYPE 01
C0011854|insulin dependent diabetes
C0011854|type I diabetes mellitus
C0011854|juvenile diabetes mellitus
C0011854|ketosis prone diabetes
C0011854|IDD
C0011854|Type 1 diabetes mellitus
C0011854|Type 1 Diabetes
C0011854|Type I Diabetes
C0011854|Juvenile Diabetes
C0011854|DIABETES MELLITUS, KETOSIS-PRONE
C0011854|KPD
C0011854|brittle diabetes (mellitus)
C0011854|juvenile onset diabetes (mellitus)
C0011854|ketosis-prone diabetes (mellitus)
C0011854|Diabetes Mellitus, Type 1 [Disease/Finding]
C0011854|Diabetes Mellitus, Brittle
C0011854|Diabetes Mellitus, Type 1
C0011854|Diabetes Mellitus, Juvenile-Onset
C0011854|Diabetes Mellitus, Sudden-Onset
C0011854|Diabetes Mellitus, Type I
C0011854|Diabetes;Type 1
C0011854|Diabetes;insulin dependent
C0011854|Diabetes;juvenile onset
C0011854|Insulin Dependent Diabetes Mellitus 1
C0011854|Juvenile Onset Diabetes
C0011854|Diabetes, Juvenile-Onset
C0011854|Juvenile-Onset Diabetes
C0011854|Diabetes Type 1
C0011854|Insulin-dependent diabetes
C0011854|Diabetes mellitus: [juvenile] or [insulin dependent]
C0011854|Diabetes mellitus - juvenile
C0011854|Diabetes mellitus: [juvenile] or [insulin dependent] (disorder)
C0011854|Diabetes mellitus type 1
C0011854|Juvenile onset diabetes mellitus
C0011854|Type I diabetes mellitus (disorder)
C0011854|IDDM - Insulin-dependent diabetes mellitus
C0011854|Insulin dependent diabetes mel
C0011854|-- Diabetes Type 1
C0011854|Diabetes mellitus Type I
C0011854|Type 1 diabetes mellitus (diagnosis)
C0011854|Diabetes mellitus juvenile onset
C0011854|Diabetes mellitus insulin-dependent
C0011854|Insulin dependent diabetic
C0011854|Diabetes mellitus type 1 (disorder)
C0011854|diabetes; insulin-dependent
C0011854|diabetes; juvenile-onset
C0011854|diabetes; ketosis-prone
C0011854|diabetes; type I
C0011854|insulin-dependent; diabetes
C0011854|juvenile-onset; diabetes
C0011854|ketosis, prone; diabetes
C0011854|type I; diabetes
C0011854|juvenile onset of diabetes
C0026769|Multiple Sclerosis
C0026769|Disseminated Sclerosis
C0026769|MS
C0026769|Sclerosis, Multiple
C0026769|insular sclerosis
C0026769|multiple sclerosis (diagnosis)
C0026769|generalized multiple sclerosis
C0026769|generalized multiple sclerosis (diagnosis)
C0026769|Sclerosis, Disseminated
C0026769|MS (Multiple Sclerosis)
C0026769|Multiple Sclerosis [Disease/Finding]
C0026769|Sclerosis;disseminated
C0026769|Multiple sclerosis NOS
C0026769|Multiple sclerosis NOS (disorder)
C0026769|Multiple sclerosis (disorder)
C0026769|Multiple sclerosis - MS
C0026769|Generalised multiple sclerosis
C0026769|Sclerosis multiple
C0026769|Neuro: Multiple Sclerosis
C0026769|DS - Disseminated sclerosis
C0026769|MS - Multiple sclerosis
C0026769|Generalized multiple sclerosis (disorder)
C0026769|cerebrospinal; sclerosis
C0026769|disseminated; sclerosis
C0026769|insular; sclerosis
C0026769|sclerosis; cerebrospinal
C0026769|sclerosis; disseminated
C0026769|sclerosis; insular
C0026769|sclerosis; multiple
C0026769|Multiple sclerosis, NOS
C0030807|Pemphigus
C0030807|Pemphigus, unspecified
C0030807|pemphigus (diagnosis)
C0030807|Pemphigus [Disease/Finding]
C0030807|Pemphigus NOS
C0030807|Pemphigus (disorder)
C0030807|Pemphigus NOS (disorder)
C0030807|Pemphigus, NOS
C0003873|Rheumatoid arthritis
C0003873|Arthritis, Rheumatoid
C0003873|Rheumatoid arthritis, unspecified
C0003873|RA
C0003873|RA (rheumatoid arthritis)
C0003873|rheumatoid arthritis (diagnosis)
C0003873|R arthritis
C0003873|Rh arthritis
C0003873|Arthritis, Rheumatoid [Disease/Finding]
C0003873|Rheumatoid arthritis NOS (disorder)
C0003873|Rheumatoid arthritis NOS
C0003873|Rheumatoid arthritis (disorder)
C0003873|Arthritis rheumatoid
C0003873|Atrophic arthritis
C0003873|Systemic rheumatoid arthritis
C0003873|Chronic rheumatic arthritis
C0003873|Rheumatic gout
C0003873|RA - Rheumatoid arthritis
C0003873|RhA - Rheumatoid arthritis
C0003873|Rheumatoid disease
C0003873|atrophic; arthritis
C0003873|rheumatoid; arthritis
C0003873|arthritis; atrophic
C0003873|arthritis; rheumatoid
C0003873|Arthritis or polyarthritis, atrophic
C0003873|Arthritis or polyarthritis, rheumatic
C0024141|SYSTEMIC LUPUS ERYTHEMATOSIS
C0024141|LUPUS, ERYTHEMATOSUS, SYSTEMIC
C0024141|Lupus Erythematosus, Systemic
C0024141|SLE
C0024141|Systemic lupus erythematosus
C0024141|Systemic lupus erythematosus, unspecified
C0024141|disseminated lupus erythematosus
C0024141|lupus
C0024141|systemic lupus erythematosus (diagnosis)
C0024141|systemic lupus
C0024141|Syst lupus erythematosus
C0024141|Systemic lupus erythematosus (SLE)
C0024141|SLE NOS
C0024141|Systemic lupus erythematosus NOS
C0024141|Lupus Erythematosus Disseminatus
C0024141|Lupus Erythematosus, Systemic [Disease/Finding]
C0024141|Systemic lupus erythematosus NOS (disorder)
C0024141|Systemic lupus erythematosus (disorder)
C0024141|Lupus erythematosis disseminated
C0024141|Syndrome lupus
C0024141|Lupus syndrome
C0024141|Syndrome disseminated lupus erythematosis
C0024141|Lupus erythematosus systemic
C0024141|LE systemic
C0024141|Systemic lupus erythematosus synd
C0024141|LE syndrome
C0024141|SLE - Systemic lupus erythematosus
C0024141|erythematosus; lupus, systemic
C0024141|lupus; erythematosus, systemic
C0024141|system; lupus erythematosus
C0024141|SLE - Lupus Erythematosus, Systemic
C0157987|allergic arthritis
C0157987|allergic arthritis (diagnosis)
C0157987|Allerg arthritis-unspec
C0157987|Arthritis;allergic
C0157987|Allergic arthritis (disorder)
C0157987|Allergic arthritis NOS (disorder)
C0157987|Allergic arthritis NOS
C0157987|Allergic arthritis of unspecified site (disorder)
C0157987|Allergic arthritis of unspecified site
C0157987|Allergic arthritis, site unspecified
C0157987|Arthritis allergic
C0157987|Arthritis allergic NOS
C0157987|allergic; arthritis
C0157987|arthritis; allergic
C0920350|Autoimmune Thyroiditides
C0920350|Lymphocytic Thyroiditides
C0920350|Lymphomatous Thyroiditides
C0920350|Lymphomatous Thyroiditis
C0920350|Thyroiditides, Autoimmune
C0920350|Thyroiditides, Lymphocytic
C0920350|Thyroiditides, Lymphomatous
C0920350|Thyroiditis, Autoimmune
C0920350|Lymphocytic Thyroiditis
C0920350|Autoimmune thyroiditis
C0920350|Thyroiditis, Autoimmune [Disease/Finding]
C0920350|Thyroiditis, Lymphomatous
C0920350|Thyroiditis, Lymphocytic
C0920350|thyroiditis autoimmune
C0920350|autoimmune thyroiditis (diagnosis)
C0920350|Lymphocytic thyroiditis (disorder)
C0920350|Autoimmune thyroiditis (disorder)
C0920350|autoimmune; thyroiditis
C0920350|thyroiditis; autoimmune
C0920350|Autoimmune thyroiditis, NOS
C0085278|Anti Phospholipid Syndrome
C0085278|Antiphospholipid Syndrome
C0085278|Syndrome, Anti-Phospholipid
C0085278|Syndrome, Antiphospholipid
C0085278|Anti Phospholipid Antibody Syndrome
C0085278|Antibody Syndrome, Anti-Phospholipid
C0085278|Antibody Syndrome, Antiphospholipid
C0085278|Antiphospholipid Antibody Syndromes
C0085278|Syndrome, Anti-Phospholipid Antibody
C0085278|Syndrome, Antiphospholipid Antibody
C0085278|antiphospholipid syndrome (diagnosis)
C0085278|Antiphospholipid Antibody Syndrome
C0085278|Anti-Phospholipid Syndrome
C0085278|Antiphospholipid Syndrome [Disease/Finding]
C0085278|Anti-Phospholipid Antibody Syndrome
C0085278|Anticardiolipin syndrome
C0085278|Antiphospholipid syndrome (disorder)
C0085278|Syndrome, Hughes
C0085278|Hughes Syndrome
C0085278|APL - Antiphospholipid syndrome
C0085278|APS - Antiphospholipid syndrome
C0085278|syndrome; anticardiolipin
C0085278|syndrome; antiphospholipid
C0085278|anticardiolipin; syndrome
C0085278|antiphospholipid; syndrome
C0031036|Polyarteritis Nodosa
C0031036|periarteritis nodosa
C0031036|panarteritis nodosa (diagnosis)
C0031036|periarteritis nodosa (diagnosis)
C0031036|panarteritis nodosa
C0031036|polyarteritis nodosa (diagnosis)
C0031036|PAN
C0031036|Polyarteritis Nodosa [Disease/Finding]
C0031036|Classical Polyarteritis Nodosa
C0031036|Polyarteritis nodosa NOS
C0031036|Systemic periarteritis nodosa
C0031036|PAN - Polyarteritis nodosa
C0031036|Polyarteritis nodosa (disorder)
C0031036|Polyarteritis nodosa NOS (disorder)
C0031036|Kussmaul's disease
C0031036|Classic polyarteritis nodosa
C0031036|Polyarteritis nodosum
C0031036|Kussmaul; disease
C0031036|disease; Kussmaul
C0342302|Brittle diabetes
C0342302|Brittle diabetes mellitus (disorder)
C0342302|Unstable diabetes mellitus
C0342302|Brittle diabetes mellitus (finding)
C0342302|Brittle diabetes mellitus
C0342302|Unstable diabetes
C0342302|Unstable diabetes mellitus (disorder)
C0342302|brittle diabetes mellitus (diagnosis)
C0342302|Diabetes brittle
C0342302|Labile diabetes
C0342302|brittle; diabetes
C0342302|diabetes; brittle
C0342302|diabetes; unstable
C0342302|unstable; diabetes
C0342302|Brittle diabetes (disorder)
C0342302|Unstable diabetes (disorder)
C0178468|autoimmune thyroid disease
C0687719|Autoimmune disease, not elsewhere classified
C0687719|Autoimmune disease NEC
C0687719|Autoimmune disease NEC in ICD9CM
C0409974|Lupus erythematosus
C0409974|Lupus erythematosis (NOS)
C0409974|Lupus erythematosus NOS
C0409974|Lupus
C0409974|Lupus erythematosus NOS (disorder)
C0409974|LE - Lupus erythematosus
C0409974|Lupus erythematosus (disorder)
C0409974|erythematosus; lupus
C0409974|lupus; erythematosus
C0024228|Diseases, Lymphatic
C0024228|Lymphatic Disease
C0024228|Lymphatic Diseases
C0024228|lymphatic disorder
C0024228|Disease, Lymphatic
C0024228|LYMPHATIC DIS
C0024228|Disease of lymphoid system
C0024228|Lymphatic Diseases [Disease/Finding]
C0024228|Lymphangiopathies
C0024228|Lymphatics--Diseases
C0024228|Disorder of lymphatic system
C0024228|disorder of lymphatic system (diagnosis)
C0024228|Lymphangiopathy
C0024228|Lymphangiopathy NOS
C0024228|Disorders of lymph node and lymphatics
C0024228|Disorder of lymphatic system (disorder)
C0024228|Disorders of lymph node and lymphatics (disorder)
C0024228|disease (or disorder); lymphatic
C0024228|Disorder of lymphatics, NOS
C0024228|Lymphangiopathy, NOS
C0024228|Disease of lymphoid system (disorder)
C0024228|Disorder of lymphatics
C0024228|Disorder of lymphoid system (disorder)
C0024228|Disorder of lymphoid system
C0024228|Lymphatic Disorders
C0011608|Dermatitis Herpetiformis
C0011608|Duhrings Disease
C0011608|Disease, Duhring's
C0011608|Disease, Duhring
C0011608|DUHRING DIS
C0011608|DUHRINGS DIS
C0011608|dermatitis herpetiformis (diagnosis)
C0011608|Duhring's disease
C0011608|Duhring Disease
C0011608|Dermatitis Herpetiformis [Disease/Finding]
C0011608|Dermatitis;herpetiformis
C0011608|Duhring-Brocq disease
C0011608|DH - Dermatitis herpetiformis
C0011608|Dermatitis herpetiformis (disorder)
C0011608|Dermatosis herpetiformis
C0011608|dermatitis; herpetiformis
C0011608|dermatosis; herpetiformis
C0011608|herpetiformis; dermatitis
C0011608|herpetiformis; dermatosis
C0011608|Duhring
C0011608|Dermatitis herpetiformis [dup] (disorder)
C0017661|Bergers Disease
C0017661|Glomerulonephritides, IGA
C0017661|Glomerulonephritis, IGA
C0017661|IgA nephropathy
C0017661|Nephropathy, Immunoglobulin A
C0017661|BERGERS DIS
C0017661|BERGER DIS
C0017661|focal glomerulonephritis
C0017661|segmental glomerulonephritis
C0017661|IGA Glomerulonephritis
C0017661|Glomerulonephritis, IGA [Disease/Finding]
C0017661|Berger Disease
C0017661|Berger's Disease
C0017661|Nephropathy, IGA
C0017661|Immunoglobulin A Nephropathy
C0017661|IGA Type Nephritis
C0017661|Nephritis, IGA Type
C0017661|Nephropathy 1, Iga
C0017661|Iga Nephropathy 1
C0017661|Immunoglobulin A nephropathy (disorder)
C0017661|IgA nephropathy (disorder)
C0017661|Glomerulonephritis focal
C0017661|nephropathy IgA
C0017661|IgA nephropathy (diagnosis)
C0017661|IgAN - IgA nephropathy
C0017661|IgA; nephropathy
C0017661|glomerulonephritis; IgA
C0017661|nephropathy; IgA
C0018213|GRAVES DISEASE
C0018213|Basedows Disease
C0018213|Disease, Basedow
C0018213|Exophthalmic Goiters
C0018213|Goiters, Exophthalmic
C0018213|Disease, Basedow's
C0018213|Disease, Graves'
C0018213|Basedow's disease
C0018213|EXOPHTHALMIC GOITER
C0018213|BASEDOW DIS
C0018213|BASEDOWS DIS
C0018213|GRAVES DIS
C0018213|Graves' disease (diagnosis)
C0018213|Graves' disease
C0018213|Graves' disease (diffuse toxic goiter)
C0018213|Disease Graves'
C0018213|Graves Disease [Disease/Finding]
C0018213|Basedow Disease
C0018213|Goiter, Exophthalmic
C0018213|Disease;Basedows
C0018213|Disease;Graves
C0018213|Exophthalmic goitre
C0018213|Hyperthyroidism, Autoimmune
C0018213|Graves' disease (disorder)
C0018213|Graves' Disease - hyperthyroidism
C0018213|Basedow's disease (disorder)
C0018213|Morbus Basedow
C0018213|Goiter exophthalmic
C0018213|Graves-Basedow disease
C0018213|Autoimmune hyperthyroidism
C0018213|Goitre exophthalmic
C0018213|Graves' disease with exophthalmos
C0018213|Toxic diffuse goiter with exophthalmos
C0018213|Toxic diffuse goitre with exophthalmos
C0018213|Toxic diffuse goiter with exophthalmos (disorder)
C0018213|Flajani
C0018213|Graves
C0018213|Basedow
C0018213|exophthalmic; goiter
C0018213|exophthalmos; goiter (etiology)
C0018213|exophthalmos; goiter (manifestation)
C0018213|goiter; exophthalmos (etiology)
C0018213|goiter; exophthalmos (manifestation)
C0018213|struma; exophthalmic
C0018213|Graves' disease [Ambiguous]
C0018213|Disease, Graves
C0029077|Sympathetic ophthalmia
C0029077|Ophthalmia, Sympathetic
C0029077|Ophthalmias, Sympathetic
C0029077|Sympathetic Ophthalmias
C0029077|Sympathetic Uveitides
C0029077|Uveitides, Sympathetic
C0029077|Sympathetic Uveitis
C0029077|sympathetic uveitis (diagnosis)
C0029077|Uveitis, Sympathetic
C0029077|Ophthalmia, Sympathetic [Disease/Finding]
C0029077|Sympathetic ophthalmitis
C0029077|Sympathetic uveitis (disorder)
C0029077|ophthalmia; sympathetic
C0029077|sympathetic; ophthalmia
C0029077|sympathetic; uveitis
C0029077|uveitis; sympathetic
C0030805|Bullous pemphigoid
C0030805|Pemphigoid
C0030805|Pemphigoid, Bullous
C0030805|Pemphigoid, unspecified
C0030805|Pemphigoids
C0030805|pemphigoid (diagnosis)
C0030805|bullous pemphigoid (diagnosis)
C0030805|Pemphigoid, Bullous [Disease/Finding]
C0030805|Pemphigoid NOS (disorder)
C0030805|Pemphigoid NOS
C0030805|Pemphigoid (disorder)
C0030805|Bullous pemphigoid NOS
C0030805|BP - Bullous pemphigoid
C0030805|Bullous pemphigoid (disorder)
C0030805|bullous; pemphigoid
C0030805|pemphigoid; bullous
C0030805|Pemphigoid, NOS
C0017665|Glomerulonephritides, Membranous
C0017665|Glomerulonephritis, Membranous
C0017665|Glomerulonephropathy, Membranous
C0017665|Glomerulopathy, Extramembranous
C0017665|Glomerulopathy, Membranous
C0017665|Membranous Glomerulonephritides
C0017665|Membranous Glomerulonephritis
C0017665|Chronic nephritic syndrome, diffuse membranous glomerulonephritis
C0017665|membranous nephropathy
C0017665|Membranous glomerulonephropathy
C0017665|nephropathy membranous
C0017665|membranous glomerulonephritis (diagnosis)
C0017665|membranous nephropathy (diagnosis)
C0017665|Glomerulonephritis membranous
C0017665|Chronic nephritic syndrome with diffuse membranous glomerulonephritis
C0017665|Membranous Glomerulopathy
C0017665|Glomerulonephritis, Membranous [Disease/Finding]
C0017665|Extramembranous Glomerulopathy
C0017665|Nephropathy, Membranous
C0017665|Chronic nephritic syndrome w diffuse membranous glomrlneph
C0017665|chronic nephritic syndrome with diffuse membranous glomerulonephritis (diagnosis)
C0017665|Membranous glomerulonephritis (disorder)
C0017665|MGN - Membranous glomerulonephritis
C0017665|Chronic nephritic syndrome, diffuse membranous glomerulonephritis (disorder)
C0017665|Membranous glomerulonephritis NOS
C0017665|Membranous nephropathy NOS
C0022972|Eaton Lambert Myasthenic Syndrome
C0022972|Eaton Lambert Syndrome
C0022972|Lambert Eaton Myasthenic Syndrome
C0022972|Lambert Eaton Syndrome
C0022972|Lambert-Eaton Myasthenic Syndrome
C0022972|Myasthenic Syndrome, Eaton-Lambert
C0022972|Syndrome, Eaton-Lambert Myasthenic
C0022972|Syndrome, Lambert-Eaton
C0022972|Syndrome, Lambert-Eaton Myasthenic
C0022972|Syndrome, Eaton-Lambert
C0022972|Eaton-Lambert syndrome
C0022972|MYOPATHIC MYASTHENIC SYNDROME OF LAMBERT EATON
C0022972|MYASTHENIC MYOPATHIC SYNDROME LAMBERT EATON
C0022972|Myasthenic Syndrome, Lambert Eaton
C0022972|Eaton-Lambert syndrome (diagnosis)
C0022972|Eaton-Lambert Myasthenic-Myopathic Syndrome
C0022972|Eaton-Lambert Myopathic-Myasthenic Syndrome
C0022972|Lambert-Eaton Myasthenic-Myopathic Syndrome
C0022972|Lambert-Eaton Myopathic-Myasthenic Syndrome
C0022972|Myopathic-Myasthenic Syndrome of Lambert-Eaton
C0022972|Lambert-Eaton Myasthenic Syndrome [Disease/Finding]
C0022972|Myasthenic-Myopathic Syndrome of Lambert-Eaton
C0022972|Eaton-Lambert Myasthenic Syndrome
C0022972|Myasthenic Syndrome, Lambert-Eaton
C0022972|Lambert-Eaton Syndrome
C0022972|Myopathic-Myasthenic Syndrome of Eaton-Lambert
C0022972|Myasthenic-Myopathic Syndrome of Eaton-Lambert
C0022972|myasthenic syndrome of Lambert Eaton
C0022972|Lambert-Eaton Myasthenic-Myopathic Syndromes
C0022972|Myasthenic Myopathic Syndrome of Eaton Lambert
C0022972|Myasthenic Myopathic Syndrome of Lambert Eaton
C0022972|Myopathic Myasthenic Syndrome of Eaton Lambert
C0022972|Lambert-Eaton syndrome NOS
C0022972|Lambert-Eaton Myopathic-Myasthenic Syndromes
C0022972|Eaton-Lambert Myopathic-Myasthenic Syndromes
C0022972|Eaton Lambert myasthenic syndrome (disorder)
C0022972|LEMS - Lambert-Eaton myasthenic syndrome
C0022972|Myasthenic syndrome
C0022972|Eaton-Lambert syndrome (disorder)
C0022972|Lambert-Eaton (etiology)
C0022972|Lambert-Eaton (manifestation)
C0022972|Eaton-Lambert (etiology)
C0022972|Eaton-Lambert (manifestation)
C0398650|Autoimmune Thrombocytopenic Purpuras
C0398650|Disease, Werlhof
C0398650|Idiopathic Thrombocytopenic Purpuras
C0398650|Purpura, Autoimmune Thrombocytopenic
C0398650|Purpura, Idiopathic Thrombocytopenic
C0398650|Purpura, Thrombocytopenic, Idiopathic
C0398650|Purpuras, Autoimmune Thrombocytopenic
C0398650|Purpuras, Idiopathic Thrombocytopenic
C0398650|Thrombocytopenic Purpura, Idiopathic
C0398650|Thrombocytopenic Purpuras, Idiopathic
C0398650|Werlhofs Disease
C0398650|Disease, Werlhof's
C0398650|Idiopathic thrombocytopenic purpura
C0398650|ITP
C0398650|Idiopathic thrombocytopenic purpura (ITP)
C0398650|THROMBOCYTOPENIC PURPURA, AUTOIMMUNE
C0398650|WERLHOF DIS
C0398650|WERLHOFS DIS
C0398650|immune thrombocytopenic purpura (diagnosis)
C0398650|immune thrombocytopenic purpura
C0398650|idiopathic thrombocytopenic purpura (diagnosis)
C0398650|ITP (idiopathic thrombocytopenic purpura)
C0398650|ITP (immune thrombocytopenic purpura)
C0398650|Idiopathic Thrombocytopenia Purpura
C0398650|Idiopathic Thrombocytopenia
C0398650|AITP
C0398650|Immune thrombocyt purpra
C0398650|Werlhof's Disease
C0398650|Purpura, Thrombocytopenic, Idiopathic [Disease/Finding]
C0398650|Werlhof Disease
C0398650|Autoimmune Thrombocytopenic Purpura
C0398650|Purpura, Thrombocytopenic, Autoimmune
C0398650|Autoimmune Thrombocytopenia
C0398650|Idiopathic purpura (& thrombocytopenic)
C0398650|Ideopath thrombocytopenic pur
C0398650|Idiopathic purpura
C0398650|ITP - idiopathic thrombocytopenic purpura
C0398650|Idiopathic purpura (& thrombocytopenic) (disorder)
C0398650|Immune Thrombocytopenias
C0398650|Purpuras, Immune Thrombocytopenic
C0398650|Thrombocytopenic Purpuras, Immune
C0398650|Thrombocytopenia, Immune
C0398650|Purpura, Immune Thrombocytopenic
C0398650|Thrombocytopenias, Immune
C0398650|Thrombocytopenias, Autoimmune
C0398650|Thrombocytopenic Purpura, Immune
C0398650|Thrombocytopenia, Autoimmune
C0398650|Immune Thrombocytopenic Purpuras
C0398650|Autoimmune Thrombocytopenias
C0398650|Immune Thrombocytopenia
C0398650|Werlhof's syndrome
C0398650|Idiopathic thrombocytopenic purpura (disorder)
C0398650|Immune thrombocytopenic purpura (disorder)
C0398650|Frank
C0398650|Werlhof
C0398650|idiopathic; purpura
C0398650|purpura; idiopathic
C0398650|purpura; thrombocytopenic, idiopathic
C0398650|thrombocytopenic; purpura, idiopathic
C0398650|ITP, NOS
C0398650|Idiopathic thrombocytopenic purpura, NOS
C0398650|Idiopathic purpura, NOS
C0398650|Idiopath Thrombocytopenic Purp
C0085409|Autoimmune Polyendocrinopathy
C0085409|Polyendocrinopathies, Autoimmune
C0085409|Polyendocrinopathy, Autoimmune
C0085409|Autoimmune polyglandular failure
C0085409|Lloyd's syndrome (diagnosis)
C0085409|Lloyd's syndrome
C0085409|polyendocrine failure syndrome (diagnosis)
C0085409|endocrine Lloyd's syndrome
C0085409|polyendocrine failure syndrome
C0085409|Autoimmune Polyendocrinopathy Syndrome
C0085409|Polyendocrinopathies, Autoimmune [Disease/Finding]
C0085409|autoimmune polyendocrine syndrome (diagnosis)
C0085409|autoimmune polyendocrine syndrome
C0085409|Lloyd's syndrome (disorder)
C0085409|Autoimmune polyglandular failure (disorder)
C0085409|PGA
C0085409|APS
C0085409|Polyendocrine autoimmunity syndrome
C0085409|Polyglandular autoimmune syndrome
C0085409|Autoimmune polyendocrinopathy (disorder)
C0085409|Autoimmune polyglandular syndrome
C0085409|autoimmune; polyglandular syndrome
C0085409|deficiency; polyglandular, autoimmune
C0085409|polyglandular; deficiency, autoimmune
C0085409|polyglandular; syndrome, autoimmune
C0085409|syndrome; autoimmune polyglandular
C0085409|syndrome; polyglandular, autoimmune
C0085409|Autoimmune polyendocrinopathy, NOS
C0085409|Autoimmune polyglandular syndrome, NOS
C0085409|Polyglandular autoimmune syndrome, NOS
C0241910|Autoimmune Hepatitides
C0241910|Autoimmune hepatitis
C0241910|Hepatitides, Autoimmune
C0241910|Hepatitis, Autoimmune
C0241910|autoimmune hepatitis (diagnosis)
C0241910|hepatitis chronic active autoimmune
C0241910|chronic active autoimmune hepatitis
C0241910|chronic active autoimmune hepatitis (diagnosis)
C0241910|Hepatitides, Autoimmune Chronic
C0241910|Hepatitis, Autoimmune Chronic
C0241910|Autoimmune Chronic Hepatitides
C0241910|Chronic Hepatitides, Autoimmune
C0241910|Chronic Hepatitis, Autoimmune
C0241910|Hepatitis, Autoimmune [Disease/Finding]
C0241910|Autoimmune Chronic Hepatitis
C0241910|Hepatitis autoimmune
C0241910|Autoimmune chronic active hepatitis
C0241910|Autoimmune hepatitis (disorder)
C0241910|autoimmune; hepatitis
C0241910|hepatitis; autoimmune
C0403529|Goodpasture's syndrome
C0403529|Anti GBM Disease
C0403529|Anti-Glomerular Basement Membrane Disease
C0403529|Syndrome, Goodpasture's
C0403529|Goodpastures Syndrome
C0403529|Syndrome, Goodpasture
C0403529|GOODPASTURE SYNDROME
C0403529|ANTI GLOMERULAR BASEMENT MEMBRANE DIS
C0403529|ANTIGBM DISEASE
C0403529|ANTIGLOMERULAR BASEMENT MEMBRANE DISEASE
C0403529|ANTI GBM DIS
C0403529|Goodpasture's syndrome (diagnosis)
C0403529|Syndrome Good pasture
C0403529|Syndrome Good postures
C0403529|Goodpasture disease
C0403529|Anti-GBM Disease
C0403529|Anti-Glomerular Basement Membrane Disease [Disease/Finding]
C0403529|Lung Purpura with Nephritis
C0403529|Anti Glomerular Basement Membrane Disease
C0403529|Goodpasture's syndrome (disorder)
C0403529|Syndrome Goodpasture's
C0403529|Pulmonary-renal syndrome
C0403529|Lung purpura with nephritis syndrome
C0403529|Anti-GBM nephritis with pulmonary hemorrhage
C0403529|Pulmonary hemorrhage with glomerulonephritis
C0403529|Pulmonary hemosiderosis with glomerulonephritis
C0403529|Anti GBM - Antiglomerular basement membrane disease
C0403529|Anti-GBM nephritis with pulmonary haemorrhage
C0403529|Goodpasture's disease
C0403529|Pulmonary haemorrhage with glomerulonephritis
C0403529|Pulmonary haemosiderosis with glomerulonephritis
C0403529|Goodpasture's disease (disorder)
C0403529|Haemorrhagic pneumonia AND glomerulonephritis
C0403529|Hemorrhagic pneumonia AND glomerulonephritis
C0403529|Goodpasture
C0403529|pulmonary; renal syndrome (Goodpasture)
C0403529|syndrome; pulmonary-renal (Goodpasture)
C0403529|Lung Purpura with Glomerulonephritis
C0751871|NEUROL AUTOIMMUNE DIS
C0751871|AUTOIMMUNE DIS NERVOUS SYSTEM
C0751871|AUTOIMMUNE NERVOUS SYSTEM DIS
C0751871|NERVOUS SYSTEM AUTOIMMUNE DIS
C0751871|AUTOIMMUNE DIS NEUROL
C0751871|Autoimmune Diseases of the Nervous System
C0751871|Autoimmune Disease, Neurologic
C0751871|Disease, Neurologic Autoimmune
C0751871|Diseases, Neurologic Autoimmune
C0751871|Neurologic Autoimmune Disease
C0751871|Autoimmune Diseases, Nervous System
C0751871|Nervous System Autoimmune Diseases
C0751871|Autoimmune Diseases of the Nervous System [Disease/Finding]
C0751871|Autoimmune Diseases, Neurologic
C0751871|Autoimmune Nervous System Diseases
C0751871|Autoimmune Disorders, Nervous System
C0751871|Neurologic Autoimmune Diseases
C0751871|Autoimmune Disorders of the Nervous System
C0751871|Autoimmune Nervous System Disorder
C0751871|Nervous system autoimmune disorders
C0004364|Autoimmune Diseases
C0004364|Disease, Autoimmune
C0004364|Diseases, Autoimmune
C0004364|autoimmune disorder
C0004364|autoimmunity
C0004364|AUTOIMMUNE DISEASE
C0004364|AUTOIMMUNE DIS
C0004364|self recognition (immune)
C0004364|autoimmune disease (diagnosis)
C0004364|Autoimmune disorders
C0004364|Autoimmune disease NOS
C0004364|Autoimmune Diseases [Disease/Finding]
C0004364|Autoimmune disease NOS (disorder)
C0004364|Autoimmune disorder NOS
C0004364|Autoimmune disease (disorder)
C0004364|Autoimmune disease, NOS
C0004364|Autoimmune disorder, NOS
C0847092|Blood autoimmune disorders
C0847092|autoimmune hematologic disorder
C0342552|Endocrine autoimmune disorders
C0342552|Autoimmune endocrine disease
C0342552|autoimmune endocrine disease (diagnosis)
C0342552|Autoimmune endocrine disease (disorder)
C0342552|autoimmune endocrine disorder
C0852003|Hepatic autoimmune disorders
C0852004|Muscular autoimmune disorders
C0852005|Lupus erythematosus and associated conditions
C0851816|Autoimmune disorders NEC
C0852006|Rheumatoid arthritis and associated conditions
C0852007|Scleroderma and associated disorders
C0949027|Skin autoimmune disorders NEC
C0036421|Progressive systemic sclerosis
C0036421|Scleroderma, Systemic
C0036421|Systemic sclerosis
C0036421|Systemic Scleroderma
C0036421|Systemic sclerosis, unspecified
C0036421|Diffuse Sclerosis
C0036421|Diffuse Scleroderma
C0036421|PSS - Progressive systemic sclerosis
C0036421|Scleroderma, Diffuse
C0036421|Sclerosis, Systemic
C0036421|Scleroderma, Systemic [Disease/Finding]
C0036421|Scleroderma;progressive
C0036421|Progressive system sclerosis
C0036421|Scleroderma syndrome (disorder)
C0036421|Scleroderma syndrome
C0036421|SSc, Diffuse Sclerosis
C0036421|SS - Systemic sclerosis
C0036421|Systemic sclerosis (disorder)
C0036421|PSS (progressive systemic sclerosis)
C0036421|sclerosis; systemic, progressive
C0036421|sclerosis; systemic
C0036421|sclerosis; system
C0036421|system; sclerosis
C0036421|systemic; sclerosis, progressive
C0036421|systemic; sclerosis
C0036421|progressive scleroderma
C2717865|Pauci Immune Vasculitis
C2717865|ANCA Associated Vasculitides
C2717865|Vasculitis, Pauci-Immune
C2717865|Vasculitides, ANCA-Associated
C2717865|Anti Neutrophil Cytoplasmic Antibody Associated Vasculitis
C2717865|Vasculitis, ANCA-Associated
C2717865|Pauci-Immune Vasculitides
C2717865|Vasculitide, ANCA-Associated
C2717865|Vasculitides, Pauci-Immune
C2717865|ANCA-Associated Vasculitide
C2717865|ANCA Associated Vasculitis
C2717865|Anti-Neutrophil Cytoplasmic Antibody-Associated Vasculitis
C2717865|Pauci-Immune Vasculitis
C2717865|ANCA-Associated Vasculitides
C2717865|ANCA-Associated Vasculitis
C2717865|Anti-Neutrophil Cytoplasmic Antibody-Associated Vasculitis [Disease/Finding]
C1328840|AUTOIMMUNE LYMPHOPROLIFERATIVE SYNDROME
C1328840|ALPS
C1328840|Autoimmun lymphprof synd
C1328840|Lymphoproliferative Syndromes, Autoimmune
C1328840|Syndromes, Autoimmune Lymphoproliferative
C1328840|Autoimmune Lymphoproliferative Syndromes
C1328840|Lymphoproliferative Syndrome, Autoimmune
C1328840|Syndrome, Autoimmune Lymphoproliferative
C1328840|Syndrome, Canale Smith
C1328840|Autoimmune lymphoproliferative syndrome [ALPS]
C1328840|Canale Smith Syndrome
C1328840|Autoimmune Lymphoproliferative Syndrome [Disease/Finding]
C1328840|Syndromes, Canale-Smith
C1328840|Canale-Smith Syndromes
C1328840|Syndrome, Canale-Smith
C1328840|Canale-Smith Syndrome
C1328840|Autoimmune Lymphoproliferative Syndrome, Type I, Autosomal Dominant
C1328840|Autoimmune lymphoproliferative syndrome (disorder)
C1328840|ALPS (autoimmune lymphoproliferative syndrome)
C0038013|Ankylosing spondylitis
C0038013|Bechterews Disease
C0038013|Marie Struempell Disease
C0038013|Spondylitis, Ankylosing
C0038013|Spondylitis, Rheumatoid
C0038013|BECHTEREW DIS
C0038013|MARIE STRUEMPELL DIS
C0038013|BECHTEREWS DIS
C0038013|ankylosing spondylitis (diagnosis)
C0038013|Ank spond
C0038013|Spondyloarthritides, Ankylosing
C0038013|Ankylosing Spondyloarthritides
C0038013|Spondylarthritides, Ankylosing
C0038013|Spondylarthritis, Ankylosing
C0038013|Spondyloarthritis, Ankylosing
C0038013|Ankylosing Spondylarthritides
C0038013|Rheumatoid arthritis of spine
C0038013|Rheumatoid Spondylitis
C0038013|Spondylarthritis Ankylopoietica
C0038013|Bechterew's Disease
C0038013|Bechterew Disease
C0038013|Marie-Struempell Disease
C0038013|Spondylitis, Ankylosing [Disease/Finding]
C0038013|Ankylosing Spondylarthritis
C0038013|Ankylosing Spondyloarthritis
C0038013|Disease;Bechterews
C0038013|Ankylosing spondylitis (disorder)
C0038013|Spondylitis Ankylopoietica
C0038013|Spondyloarthritis Ankylopoietica
C0038013|Spondylitis ankylosing
C0038013|Bekhterev's disease
C0038013|AS - Ankylosing spondylitis
C0038013|Idiopathic ankylosing spondylitis
C0038013|Marie-Strumpell spondylitis
C0038013|Marie Strümpell spondylitis
C0038013|arthritis; spine or vertebra, Marie-Strümpell
C0038013|arthritis; spine or vertebra, ankylosing
C0038013|Marie-Strümpell; spondylitis
C0038013|Marie-Strümpell
C0038013|Strümpell-Marie
C0038013|Von Bechterew
C0038013|Bechterew
C0038013|rheumatoid; arthritis, spine
C0038013|rheumatoid; spondylitis
C0038013|spine or vertebra; arthritis, Marie-Strümpell
C0038013|spine or vertebra; arthritis, ankylosing
C0038013|spondylitis; Marie-Strümpell
C0038013|spondylitis; ankylopoietica
C0038013|spondylitis; ankylosing
C0038013|spondylitis; rheumatoid
C0038013|ankylopoietica; spondylitis
C0038013|ankylosing; spondylitis
C0038013|arthritis; rheumatoid, spine
C0038013|Ankylosing spondylitis, NOS
C0038013|Rheumatoid arthritis of spine, NOS
C0038013|Spondylitis, Marie-Strumpell
C0038013|Rheumatioid arthritis of spine NOS
C0026272|Mixed Connective Tissue Disease
C0026272|Syndrome, Sharp
C0026272|CONNECTIVE TISSUE DIS MIXED
C0026272|MIXED CONNECTIVE TISSUE DIS
C0026272|mixed connective tissue disease (diagnosis)
C0026272|Mixed Connective Tissue Disease [Disease/Finding]
C0026272|Sharp Syndrome
C0026272|MCTD
C0026272|Connective Tissue Disease, Mixed
C0026272|Mixed collagen vascular disease (disorder)
C0026272|Connective tissue disease overlap syndrome
C0026272|Sharp's syndrome
C0026272|Mixed collagen vascular disease
C0026272|MCTD - Mixed connective tissue disease
C0026272|Connective tissue disease overlap syndrome (disorder)
C0026272|disease (or disorder); mixed connective tissue
C0026272|disease (or disorder); mixed, connective tissue
C0026272|disease; mixed connective tissue
C0026272|mixed, connective tissue; disorder
C0026272|Mixed collagen vascular disease, NOS
C0026272|Mixed connective tissue disease, NOS
C2609059|Antisynthetase syndrome
C2609059|Antisynthetase syndrome (disorder)
C0554876|poorly controlled diabetes mellitus (diagnosis)
C0554876|diabetes mellitus poorly controlled
C0554876|poorly controlled diabetes mellitus
C2930824|Autoimmune limbic encephalitis
C1260879|Autoimmune progesterone dermatitis
C1260879|Progesterone dermatitis
C1260879|Autoimmune progesterone urticaria
C1260879|Autoimmune progesterone dermatitis/urticaria (disorder)
C1260879|Autoimmune progesterone dermatitis/urticaria
C0301928|Psychogenic purpura
C0301928|Autoerythrocyte sensitization
C0301928|Gardner-Diamond syndrome
C0301928|Painful bruising syndrome
C0301928|Autoerythrocyte sensitivity disorder
C0301928|Auto-erythrocyte sensitization
C0301928|Auto-erythrocyte sensitisation
C0301928|Autoerythrocyte sensitivity disorder (finding)
C0301928|Autoerythrocyte sensitivity
C0301928|Gardner-Diamond syndrome (disorder)
C0301928|Auto-erythrocyte sensitisation syndrome
C0301928|Auto-erythrocyte sensitization syndrome
C0301928|Autoerythrocyte sensitivity (finding)
C0301928|autoerythrocyte sensitization; syndrome
C0301928|Gardner-Diamond
C0301928|syndrome; autoerythrocyte sensitization
C0301928|Gardener-Diamond syndrome
C0301928|Autoerythrocyte sensitivity disorder, NOS
C0432222|SPONDYLOENCHONDRODYSPLASIA
C0432222|SEM
C0432222|Spondyloenchondromatosis
C0432222|Spondylometaphyseal dysplasia with enchondromatous changes
C0432222|SPENCD
C0432222|Spondyloenchondrodysplasia (disorder)
C0432222|Spondyloenchondromatosis (disorder)
C2931429|Pediatric Autoimmune Neuropsychiatric Disorders Associated with Streptococcal infections
C2931429|PANDAS - Paediatric autoimmune neuropsychiatric disorder associated with streptococcal infection
C2931429|Paediatric autoimmune neuropsychiatric disorder associated with streptococcal infection
C2931429|Pediatric autoimmune neuropsychiatric disorder associated with streptococcal infection
C2931429|Pediatric autoimmune neuropsychiatric disorder associated with streptococcal infection (disorder)
C2931429|PANDAS - Pediatric autoimmune neuropsychiatric disorder associated with streptococcal infection
C2931429|Paediatric autoimmune neuropsychiatric disorders associated with streptococcal infection
C2931429|Pediatric autoimmune neuropsychiatric disorders associated with streptococcal infection
C2931429|PANDAS
C0341305|Autoimmune enteropathy
C0341305|Autoimmune enteropathy (disorder)
C0406650|Linear IgA disease
C0406650|linear IgA dermatoses (diagnosis)
C0406650|linear IgA dermatoses
C0406650|linear IgA dermatosis
C0406650|IgA Dermatoses, Linear
C0406650|Linear IgA Bullous Dermatosis
C0406650|Dermatosis, Linear IgA
C0406650|IgA Dermatosis, Linear
C0406650|Dermatoses, Linear IgA
C0406650|Linear IgA Bullous Dermatosis [Disease/Finding]
C0406650|Linear immunoglobulin A dermatosis (disorder)
C0406650|Linear IgA dermatosis (disorder)
C0406650|Linear immunoglobulin A dermatosis
C0406650|Linear IgA
C0406650|Linear Ig A disease
C0406650|IgA - Linear immunoglobulin A bullous dermatosis
C0406650|LAD - Linear IgA disease
C0406650|Linear immunoglobulin A bullous dermatosis
C0342340|Autoimmune parathyroiditis
C0342340|Autoimmune parathyroiditis (disorder)
C0034152|Purpura, Schoenlein Henoch
C0034152|Purpura, Schoenlein-Henoch
C0034152|Schoenlein Henoch Purpura
C0034152|Allergic purpura
C0034152|Henoch-Schonlein purpura
C0034152|Purpura, Allergic
C0034152|Purpura, Anaphylactoid
C0034152|Henoch-Schoenlein purpura
C0034152|Henoch-Schonlein purpura (disorder)
C0034152|Anaphylactoid purpura
C0034152|Purpura, Henoch
C0034152|Henoch-Scholein purpura
C0034152|Henoch-Sch@nlein purpura
C0034152|allergic purpura (diagnosis)
C0034152|allergic vascular purpura (diagnosis)
C0034152|Henoch Schoenlein Purpura
C0034152|Purpura, Henoch-Schoenlein
C0034152|allergic vascular purpura
C0034152|Henoch Schonlein purpura
C0034152|Henoch Schonlein purpura (diagnosis)
C0034152|vascular allergic purpura
C0034152|Purpuras, Schonlein-Henoch
C0034152|Schonlein-Henoch Purpuras
C0034152|Purpuras, Henoch-Schonlein
C0034152|Henoch Schonlein Purpuras
C0034152|Purpura, Schonlein Henoch
C0034152|Henoch-Schonlein Purpuras
C0034152|Purpura, Henoch Schonlein
C0034152|Schonlein Purpura, Henoch
C0034152|Schonlein Purpuras, Henoch
C0034152|Schonlein-Henoch Purpura
C0034152|Purpuras, Henoch Schonlein
C0034152|Purpura, Henoch-Schonlein
C0034152|Schoenlein-Henoch Purpura
C0034152|Purpura Henoch(-Schönlein)
C0034152|Purpura anaphylactoid
C0034152|Purpura, Schoenlein-Henoch [Disease/Finding]
C0034152|Henoch Purpura
C0034152|Purpura, Schonlein-Henoch
C0034152|Henoch-Sch?nlein purpura
C0034152|Autoimmune purpura
C0034152|Allergic purpura (disorder)
C0034152|Autoimmune purpura (disorder)
C0034152|Henoch-Schonlein all. purpura
C0034152|Allergic purpura NOS (disorder)
C0034152|Purpura: [allergic] or [Henoch-Schonlein allergy]
C0034152|Purpura: [allergic] or [Henoch-Schonlein allergy] (disorder)
C0034152|Henoch-Sch?nlein purpura (disorder)
C0034152|Allergic purpura NOS
C0034152|Anaphylactic vascular purpura
C0034152|Purpura allergic
C0034152|Purpura vascular allergic
C0034152|Anaphylactoid vascular purpura
C0034152|Henoch-Schonlein
C0034152|Henoch Shonlein purpura
C0034152|HSP
C0034152|Henoch's purpura
C0034152|Acute vascular purpura
C0034152|Henoch-Schoenlein vasculitis
C0034152|Spring fever
C0034152|HSP - Henoch-Schonlein purpura
C0034152|Schönlein; purpura
C0034152|Schönlein
C0034152|allergic; purpura
C0034152|purpura; Schönlein
C0034152|purpura; allergic
C0034152|purpura; anaphylactoid
C0034152|anaphylactoid; purpura
C0034152|Autoimmune purpura (disorder) [Ambiguous]
C0034152|Purpura, autoimmune
C0034152|Purpura;Henoch-Schonlein
C0272177|Neutropenia associated with autoimmune disease
C0272177|neutropenia associated with autoimmune disease (diagnosis)
C0272177|Neutropenia associated with autoimmune disease (disorder)
C3495559|Chronic Arthritis, Juvenile
C3495559|Rheumatoid Arthritis, Juvenile
C3495559|Juvenile arthritis
C3495559|Juvenile arthritis, unspecified
C3495559|Arthritis, Juvenile Chronic
C3495559|Juvenile Idiopathic Arthritis
C3495559|Juvenile Chronic Arthritis
C3495559|Juvenile Rheumatoid Arthritis
C3495559|Arthritis, Juvenile Idiopathic
C3495559|juvenile arthritis (diagnosis)
C3495559|Arthritis, Juvenile
C3495559|Enthesitis Related Arthritis, Juvenile
C3495559|Juvenile Oligoarthritis
C3495559|Arthritis, Juvenile Systemic
C3495559|Juvenile Enthesitis-Related Arthritis
C3495559|Juvenile Systemic Arthritis
C3495559|Arthritis, Juvenile Psoriatic
C3495559|Juvenile Psoriatic Arthritis
C3495559|Arthritis, Juvenile Enthesitis-Related
C3495559|Oligoarthritis, Juvenile
C3495559|Arthritis, Juvenile Rheumatoid
C3495559|Enthesitis-Related Arthritis, Juvenile
C3495559|Psoriatic Arthritis, Juvenile
C3495559|Systemic Arthritis, Juvenile
C3495559|Arthritis, Juvenile [Disease/Finding]
C3495559|JIA
C3495559|Polyarthritis, Juvenile, Rheumatoid Factor Positive
C3495559|Polyarthritis, Juvenile, Rheumatoid Factor Negative
C3495559|JCA - Juvenile chronic arthritis
C3495559|Juvenile chronic arthritis (disorder)
C3495559|juvenile; arthritis
C3495559|arthritis; juvenile
C3495559|Juvenile chronic arthritis, polyarticular seropositive
C3495559|Juvenile idiopathic arthritis (disorder)
C3495559|Juvenile idiopathic arthritis, polyarthritis, rheumatoid factor positive
C3495559|Idiopathic Arthritis, Juvenile
C3495559|Arthritis;juvenile
C2732697|Autoimmune inflammation of skeletal muscle (disorder)
C2732697|Autoimmune inflammation of skeletal muscle
C2732697|Autoimmune myositis
C1328843|Autoimmune vasculitis
C1328843|Autoimmune vasculitis (disorder)
C1328843|Immune mediated vasculitis
C2609129|Autoimmune pancreatitis
C2609129|Autoimmune pancreatitis (disorder)
C0456037|ANT - Autoimmune neonatal thrombocytopenia
C0456037|Autoimmune neonatal thrombocytopenia
C0456037|Autoimmune neonatal thrombocytopenia (disorder)
C0342337|Insulin resistance - type B
C0342337|Insulin resistance - type B (disorder)
C0400936|Autoimmune liver disease
C0400936|Autoimmune liver disease (disorder)
C1970472|PULMONARY ALVEOLAR PROTEINOSIS, ACQUIRED
C1970472|Pulmonary Alveolar Lipoproteinosis, Acquired
C1970472|Pulmonary Alveolar Proteinosis, Autoimmune
C1970472|Autoimmune pulmonary alveolar proteinosis (disorder)
C1970472|Autoimmune pulmonary alveolar proteinosis
C1970472|PAP, ACQUIRED
C1842763|SPONDYLOENCHONDRODYSPLASIA WITH IMMUNE DYSREGULATION
C1842763|SPENCDI
C1842763|Combined Immunodeficiency with Autoimmunity and Spondylometaphyseal Dysplasia
C1842763|Spondyloenchondrodysplasia with immune dysregulation (disorder)
C1842763|Roifman-Melamed syndrome
C1842763|Roifman-Costa syndrome
C0272137|Galactosyltransferase Deficiency
C0272137|Tn Syndrome
C0272137|TN POLYAGGLUTINATION SYNDROME
C0272137|TNPS
C0272137|Polyagglutinable erythrocyte syndrome
C0272137|Polyagglutinable erythrocyte syndrome (disorder)
C1835931|ALPHA/BETA T-CELL LYMPHOPENIA WITH GAMMA/DELTA T-CELL EXPANSION, SEVERE CYTOMEGALOVIRUS INFECTION, AND AUTOIMMUNITY
C1835931|Alpha-Beta T-Cell Lymphopenia with Gamma-Delta T-Cell Expansion, Severe Cytomegalovirus Infection, and Autoimmunity
C1857958|DIABETES MELLITUS, CONGENITAL AUTOIMMUNE
C0026103|Mikulicz's disease
C0026103|Mikulicz's syndrome
C0026103|Disease, Mikulicz
C0026103|Disease, Mikulicz'
C0026103|Mikulicz' Disease
C0026103|MIKULICZ DIS
C0026103|Mikulicz's disease (diagnosis)
C0026103|Mikulicz disease
C0026103|Mikulicz' Disease [Disease/Finding]
C0026103|Mikulicz syndrome
C0026103|Mikulicz's disease (disorder)
C0026103|Mikulicz
C2717757|Syndrome, Susac
C2717757|Susacs Syndrome
C2717757|Vasculopathies, Retinocochleocerebral
C2717757|Retinocochleocerebral Vasculopathies
C2717757|Syndrome, Susac's
C2717757|Susac Syndrome
C2717757|Vasculopathy, Retinocochleocerebral
C2717757|Susac Syndrome [Disease/Finding]
C2717757|Retinocochleocerebral Vasculopathy
C2717757|Susac's Syndrome
C2717757|Retinocochleocerebral vasculopathy (disorder)
C0409999|Undifferentiated connective tissue disease
C0409999|UCTD
C0409999|Undifferentiated connective tissue disease (disorder)
C1861303|ACUG
C1861303|SYNOVITIS, GRANULOMATOUS, WITH UVEITIS AND CRANIAL NEUROPATHIES (disorder)
C1861303|SYNOVITIS, GRANULOMATOUS, WITH UVEITIS AND CRANIAL NEUROPATHIES
C1861303|BLAU SYNDROME
C1861303|Granulomatous inflammatory arthritis, dermatitis, and uveitis, familial
C1861303|Granulomatosis, familial, Blau type
C1861303|Arthrocutaneouveal granulomatosis
C1861303|Granulomatosis, familial juvenile systemic
C1861303|Jabs syndrome
C1861303|Familial granulomatosis, Blau type
C1861303|Arthrocutaneouveal granulamotosis
C1861303|Granulomatous inflammatory arthritis, dermatitis and uveitis, familial
C1861303|Familial juvenile systemic granulomatosis
C1861303|Early onset sarcoidosis
C1861303|Pediatric granulomatous arthritis
C1861303|Familial granulomatous inflammatory arthritis, dermatitis and uveitis (disorder)
C1861303|Familial granulomatous inflammatory arthritis, dermatitis and uveitis
C1861303|Early-Onset Sarcoidosis
C1861303|BLAUS
C1861303|Synovitis granulomatous with uveitis and cranial neuropathies
C0410000|Overlap syndrome
C0410000|Overlap syndrome (disorder)
C0393799|Miller Fisher Syndrome
C0393799|Syndrome, Fisher
C0393799|Syndrome, Miller Fisher
C0393799|Syndrome, Miller-Fisher
C0393799|Miller-Fisher syndrome (diagnosis)
C0393799|Miller-Fisher syndrome
C0393799|Fisher syndrome
C0393799|Guillain-Barre Syndrome, Miller Fisher Variant
C0393799|Miller Fisher Syndrome [Disease/Finding]
C0393799|Miller Fisher Variant of Guillain Barre Syndrome
C0393799|Guillain Barre Syndrome, Miller Fisher Variant
C0393799|Ophthalmoplegia, Ataxia and Areflexia Syndrome
C0393799|Miller-Fisher variant of Guillain-Barre syndrome (disorder)
C0393799|Miller-Fisher variant of Guillain-Barre syndrome
C0393799|Fisher's syndrome
C0393799|Ophthalmoplegia, ataxia, areflexia syndrome
C0393799|Fisher's syndrome (disorder)
C0265235|Marshall syndrome
C0265235|Deafness, myopia, cataract, saddle nose-Marshall type
C0265235|PFAPA syndrome
C0265235|pfapa syndrome (diagnosis)
C0265235|MRSHS
C0265235|Periodic Fever, Aphthous Stomatitis, Pharyngitis, Adenitis Syndrome
C0265235|Syndrome of periodic fever, aphthous stomatitis, pharyngitis, cervical adenitis
C0265235|Marshall's syndrome
C0265235|Marshall syndrome (disorder)
C0340971|Autoimmune neutropenia
C0340971|neutropenia autoimmune
C0340971|Autoimmune neutropenia (diagnosis)
C0340971|Autoimmune neutropenia (disorder)
C0677607|Hashimoto's disease
C0677607|HASHIMOTO THYROIDITIS
C0677607|lymphomatous thyroiditis
C0677607|HASHIMOTOS DIS
C0677607|HASHIMOTO DIS
C0677607|Hashimoto's thyroiditis
C0677607|Hashimoto's thyroiditis (diagnosis)
C0677607|Chr lymphocyt thyroidit
C0677607|Hashimoto's Syndromes
C0677607|Hashimotos Syndrome
C0677607|Syndromes, Hashimoto's
C0677607|Hashimoto Syndrome
C0677607|Syndrome, Hashimoto's
C0677607|Struma lymphomatosa
C0677607|Hashimoto Disease [Disease/Finding]
C0677607|Hashimoto Disease
C0677607|Chronic Lymphocytic Thyroiditis
C0677607|Hashimoto's Syndrome
C0677607|Disease;Hashimotos
C0677607|Hashimoto Struma
C0677607|Struma lymphomatosis (disorder)
C0677607|Hashimoto's thyroiditis (disorder)
C0677607|Struma lymphomatosis
C0677607|Hashimoto's Struma
C0677607|autoimmune thyroiditis
C0677607|HT
C0677607|Lymphocytic thyroiditis
C0677607|Autoimmune lymphocytic chronic thyroiditis
C0677607|Hashimoto thyroiditis (disorder)
C0677607|Hashimoto; thyroiditis
C0677607|Hashimoto
C0677607|chronic; thyroiditis, lymphadenoid
C0677607|lymphocytic; thyroiditis
C0677607|lymphoid; thyroiditis
C0677607|lymphomatosa; goiter
C0677607|lymphomatous; thyroiditis
C0677607|struma; lymphomatosa
C0677607|thyroiditis; Hashimoto
C0677607|thyroiditis; chronic, lymphadenoid
C0677607|thyroiditis; lymphocytic
C0677607|thyroiditis; lymphoid
C0677607|thyroiditis; lymphomatous
C0677607|Disease, Hashimoto
C0677607|Hashimotos Disease
C0677607|Disease, Hashimoto's
C0677607|Chronic Lymphocytic Thyroiditides
C0677607|Hashimoto Thyroiditides
C0677607|Lymphocytic Thyroiditides, Chronic
C0677607|Lymphocytic Thyroiditis, Chronic
C0677607|Thyroiditides, Chronic Lymphocytic
C0677607|Thyroiditides, Hashimoto
C0677607|Thyroiditis, Chronic Lymphocytic
C0677607|Thyroiditis, Hashimoto
C4022660|Autoimmune antibody positivity
C0242584|Autoimmune thrombocytopenia
C0242584|Auto-immune thrombocytopenia
C0242584|Thrombocytopenia, autoimmune
C0242584|Thrombocytopenia (& [auto-immune])
C0242584|Autoimmune thrombocytopenia (disorder)
C0242584|Thrombocytopenia (& [auto-immune]) (procedure)
C0242584|Thrombocytopenia (& [auto-immune]) (finding)
C0242584|Immune thrombocytopenia
C0342410|Autoimmune Hypophysitis
C0342410|Hypophysitides, Autoimmune
C0342410|Lymphoid Hypophysitides
C0342410|Hypophysitis, Lymphoid
C0342410|Lymphocytic Hypophysitides
C0342410|Hypophysitides, Lymphoid
C0342410|Hypophysitides, Lymphocytic
C0342410|Autoimmune Hypophysitides
C0342410|Autoimmune Hypophysitis [Disease/Finding]
C0342410|Hypophysitis, Lymphocytic
C0342410|Hypophysitis, Autoimmune
C0342410|Lymphocytic Hypophysitis
C0342410|Lymphoid Hypophysitis
C0342410|Autoimmune hypophysitis (disorder)
C0393639|Hashimoto's encephalopathy
C0393639|Hashimoto's encephalitis
C0393639|Steroid-responsive encephalopathy associated with autoimmune thyroiditis
C0393639|Autoimmune encephalitis
C0393639|Encephalitis autoimmune
C0393639|Autoimmune encephalopathy
C0393639|Encephalitis allergic (autoimmune)
C0393639|Autoimmune encephalitis (disorder)
C0393639|Autoimmune encephalitis, NOS
C4075851|Autoimmune cholangitis (disorder)
C4075851|Autoimmune cholangitis
C0271893|Autoimmune pancytopenia
C0271893|pancytopenia autoimmune
C0271893|pancytopenia autoimmune (diagnosis)
C0271893|Autoimmune pancytopenia (disorder)
C0543694|Autoimmune leukopenia
C0543694|Autoimmune leucopenia
C0543694|Autoimmune leukopenia (disorder)
C0395947|Autoimmune disorder of inner ear
C0395947|Autoimmune labyrinthitis
C0395947|Autoimmune disorder of inner ear (disorder)
C0406632|Autoimmune diseases affecting skin
C0406632|Autoimmune skin disease (disorder)
C0406632|Autoimmune skin disease
C0406632|Autoimmune skin disease, NOS
C0086981|Sicca Syndrome
C0086981|Syndrome, Sicca
C0086981|xerodermosteosis
C0086981|sicca syndrome (diagnosis)
C0086981|SICCA
C0086981|Sicca syndrome, unspecified
C0086981|Sicca syndrome (disorder)
C0086981|Syndrome sicca
C0086981|sicca; syndrome
C0086981|syndrome; sicca
C1328835|autoimmune dermatologic disorder
C1328836|autoimmune gastrointestinal and liver disorder
C1328837|autoimmune genitourinary disorder
C1328837|autoimmune urogenital disorder
C1328837|urogenital autoimmune disorder
C1328841|autoimmune respiratory disorder
C1328842|autoimmune rheumatologic disease
C0175816|Cold type haemolytic anaemia
C0175816|COLD AGGLUTININ DIS
C0175816|Cold Hemagglutinin Disease
C0175816|cold antibody hemolytic anemia
C0175816|hemolytic anemia due to cold agglutinin disease (diagnosis)
C0175816|hemolytic anemia due to cold agglutinin disease
C0175816|cold agglutinin disease
C0175816|Diseases, Cold Antibody
C0175816|Disease, Cold Antibody
C0175816|Cold Antibody Diseases
C0175816|Haemolytic anaemia due to cold antibody
C0175816|Cryopathic hemolytic anemia
C0175816|Cold haemagglutinin disease
C0175816|AIHA - Cold autoimmune hemolytic anemia
C0175816|Hemolytic anemia due to cold antibody
C0175816|Cold autoimmune hemolytic anemia (disorder)
C0175816|Cold autoimmune haemolytic anaemia
C0175816|CHAD - Cold hemagglutinin disease
C0175816|Cold autoimmune hemolytic anemia
C0175816|AIHA - Cold autoimmune haemolytic anaemia
C0175816|Cold type hemolytic anemia
C0175816|Cold hemolytic disease
C0175816|Cold antibody haemolytic anaemia
C0175816|Cryopathic haemolytic anaemia
C0175816|Cold haemolytic disease
C0175816|Cold haemagglutinin disease (disorder)
C0175816|CHAD - Cold haemagglutinin disease
C0175816|Anemia, Hemolytic, Cold Antibody
C0175816|Cold Antibody Disease
C0175816|Hemolytic anemia due to cold antibody, NOS
C0175816|Agglutinin Disease, Cold
C0175816|Agglutinin Diseases, Cold
C0175816|Cold Agglutinin Diseases
C0175816|Disease, Cold Agglutinin
C0175816|Diseases, Cold Agglutinin
C0037997|Disease, Splenic
C0037997|Diseases, Splenic
C0037997|Splenic Disease
C0037997|Splenic Diseases
C0037997|spleen disorder
C0037997|Disease of spleen, unspecified
C0037997|Diseases of spleen
C0037997|SPLENIC DIS
C0037997|Disease of spleen
C0037997|splenic disorders (diagnosis)
C0037997|splenic disorders
C0037997|Spleen disorders
C0037997|Spleen disease NOS
C0037997|Splenic Diseases [Disease/Finding]
C0037997|Disease;spleen
C0037997|Spleen Diseases
C0037997|Splenic Diseaess
C0037997|Spleen disease
C0037997|Disease of spleen NOS
C0037997|Disease of spleen unspecified (disorder)
C0037997|Disease of spleen NOS (disorder)
C0037997|Disease of spleen unspecified
C0037997|Splenopathy
C0037997|Spleen--Diseases
C0037997|Disorder spleen
C0037997|Spleen disorder NOS
C0037997|Dyssplenism
C0037997|Splenic disorder
C0037997|disease (or disorder); spleen
C0037997|spleen; disease
C0037997|spleen; hyperfunction
C0037997|Disease of spleen, NOS
C0037997|Splenic disorder, NOS
C0037997|Splenic syndrome, NOS
C0037997|Disorder of spleen
C0037997|Disease of spleen (disorder)
C0037997|Disorder of spleen (disorder)
C0011644|Scleroderma
C0011644|dermatosclerosis
C0011644|scleroderma (diagnosis)
C0011644|Scleroderma (disorder)
C0011644|Scleroderma NOS
C0011644|Scleroderma NOS (disorder)
C0011644|Scleroderma (Disease)
C0011644|Progressive systemic scleroderma
C0011633|Dermatomyositides
C0011633|Dermatomyositis
C0011633|Dermatopolymyositis
C0011633|Dermatopolymyositis, unspecified
C0011633|Polymyositis Dermatomyositis
C0011633|Polymyositis-Dermatomyositides
C0011633|Dermatopolymyositides
C0011633|Dermatopolymyositis, unspecified, organ involvement unspecified
C0011633|Polymyositis-Dermatomyositis
C0011633|Dermatomyositis [Disease/Finding]
C0011633|Dermatopolymyositis, unsp, organ involvement unspecified
C0011633|[X]Dermatopolymyositis, unspecified
C0011633|Polymyositis with skin involvement
C0011633|DM - Dermatomyositis
C0011633|Dermatomyositis (disorder)
C0011633|[X]Dermatopolymyositis, unspecified (disorder)
C0011633|Wagner-Unverricht syndrome
C0011633|Dermatopolymyositis (diagnosis)
C0011633|polymyositis/dermatomyositis
C0011633|dermatomyositis (diagnosis)
C0011633|polymyositis; with involvement of skin
C0011633|dermatomucosomyositis
C0036202|Disease, Schaumann
C0036202|Sarcoid, Boeck's
C0036202|Sarcoidoses
C0036202|Sarcoidosis
C0036202|Besnier Boeck Disease
C0036202|Boeck Sarcoid
C0036202|Boecks Sarcoid
C0036202|Sarcoidosis, unspecified
C0036202|Boeck's sarcoidosis
C0036202|Boecks sarcoidosis
C0036202|SCHAUMANN DIS
C0036202|BESNIER BOECK DIS
C0036202|lymphogranulomatosis (benign)
C0036202|sarcoidosis (diagnosis)
C0036202|benign lymphogranulomatosis
C0036202|Boeck's sarcoid
C0036202|benign lymphogranulomatosis (diagnosis)
C0036202|benign lymphogranulomatosis of Schaumann
C0036202|Syndrome, Besnier-Boeck-Schaumann
C0036202|Syndrome, Schaumann
C0036202|Schaumann's Syndromes
C0036202|Besnier Boeck Schaumann Syndrome
C0036202|Boecks Disease
C0036202|Syndrome, Schaumann's
C0036202|Schaumann Disease
C0036202|Sarcoidosis [Disease/Finding]
C0036202|Besnier-Boeck Disease
C0036202|Boeck Disease
C0036202|Schaumann Syndrome
C0036202|Besnier-Boeck-Schaumann Syndrome
C0036202|Schaumann's Syndrome
C0036202|Boeck's Disease
C0036202|lymphogranulomatosis
C0036202|Sarcoidosis (disorder)
C0036202|sarcoid
C0036202|Schaumann's disease
C0036202|Besnier-Boeck-Schaumann's disease
C0036202|Sarcoidosis NOS
C0036202|Darier-Roussy sarcoid
C0036202|Lupus pernio of Besnier
C0036202|Miliary lupoid of Boeck
C0036202|benign; lymphogranulomatosis
C0036202|Hutchinson-Boeck
C0036202|Schaumann; benign lymphogranulomatosis
C0036202|Schaumann; disease or syndrome
C0036202|Besnier-Boeck
C0036202|Besnier; lupus pernio
C0036202|Boeck; disease
C0036202|Boeck; sarcoid
C0036202|lymphogranulomatosis; benign
C0036202|sarcoid; Boeck
C0036202|sarcoid; Darier-Roussy
C0036202|syndrome; Schaumann
C0036202|Darier-Roussy; sarcoid
C0036202|Sarcoidosis, NOS
C0036202|Besnier-Boeck-Schaumann disease
C0036202|Boeck Sarcoid, any site
C0036202|Benign Lymphogranulomatosis, Schaumann's
C0036202|Lupus pernio, Besnier
C0036202|Sarcoid NOS
C0272126|Evans syndrome
C0272126|Evans' syndrome (diagnosis)
C0272126|Evans' syndrome
C0272126|Autoimmune hemolytic anemia and autoimmune thrombocytopenia
C0272126|Evan's syndrome
C0272126|Evans syndrome (disorder)
C0272126|Evans
C0266995|benign lymphoepithelial lesion of salivary gland (diagnosis)
C0266995|benign lymphoepithelial lesion of salivary gland
C0266995|Benign lymphoepithelial salivary gland lesion
C0266995|Benign lymphoepithelial lesion of salivary gland (disorder)
C0266995|lesion; salivary gland, benign lymphoepithelial
C0266995|salivary gland; lesion, benign lymphoepithelial
C0266995|Godwin Tumor
C0266995|Benign Lymphoepithelial Lesion of the Salivary Gland
C0266995|Benign Salivary Gland Lymphoepithelial Lesion
C1841911|GLUTAMIC ACID DECARBOXYLASE, BRAIN, MEMBRANE FORM
C0031069|Disease, Periodic
C0031069|Familial Mediterranean Fever
C0031069|Benign paroxysmal peritonitis
C0031069|Recurrent polyserositis
C0031069|FMF
C0031069|WOLFFS PERIODIC DIS
C0031069|WOLFF PERIODIC DIS
C0031069|PERIODIC DIS WOLFFS
C0031069|PERIODIC DIS
C0031069|familial Mediterranean fever (diagnosis)
C0031069|familial Mediterranean fever with recurrent polyserositis
C0031069|familial Mediterranean fever with recurrent polyserositis (diagnosis)
C0031069|Disease, Wolff Periodic
C0031069|Disease, Wolff's Periodic
C0031069|Periodic Disease, Wolff
C0031069|Wolffs Periodic Disease
C0031069|Fam Mediterranean fever
C0031069|Diseases, Periodic
C0031069|Periodic Disease, Wolffs
C0031069|Periodic Diseases
C0031069|Wolff Periodic Disease
C0031069|Periodic Disease, Wolff's
C0031069|Familial Mediterranean Fever [Disease/Finding]
C0031069|Wolff's Periodic Disease
C0031069|Mediterranean Fever, Familial
C0031069|Periodic Disease
C0031069|Peritonitis, Periodic
C0031069|Peritonitides, Benign Paroxysmal
C0031069|Peritonitis, Benign Paroxysmal
C0031069|Familial Paroxysmal Polyserositides
C0031069|Periodic Peritonitides
C0031069|Peritonitides, Periodic
C0031069|Paroxysmal Polyserositis, Familial
C0031069|Paroxysmal Peritonitides, Benign
C0031069|Paroxysmal Polyserositides, Familial
C0031069|Benign Paroxysmal Peritonitides
C0031069|Paroxysmal Peritonitis, Benign
C0031069|Polyserositides, Familial Paroxysmal
C0031069|Polyserositides, Recurrent
C0031069|Recurrent Polyserositides
C0031069|Periodic Peritonitis
C0031069|Familial Paroxysmal Polyserositis
C0031069|Polyserositis, Recurrent
C0031069|Polyserositis, Familial Paroxysmal
C0031069|Familial Mediterranean Fever, Autosomal Recessive
C0031069|familial mediterranean fever autosomal recessive
C0031069|FMF autosomal recessive
C0031069|familial mediterranean fever autosomal recessive (diagnosis)
C0031069|Familial recurrent polyserositis
C0031069|Paroxysmal polyserositis
C0031069|FMF - Familial Mediterranean fever
C0031069|Periodic familial peritonitis
C0031069|Periodic polyserositis
C0031069|MEF - Familial Mediterranean fever
C0031069|Familial Mediterranean fever (disorder)
C0031069|fever; mediterranean, familial
C0031069|mediterranean; fever, familial
C0031069|periodic; peritonitis
C0031069|periodic; polyserositis
C0031069|peritonitis; periodic
C0031069|polyserositis; periodic
C0031069|Periodic fever
C0267807|Lupus hepatitis
C0267807|Lupoid hepatitis
C0267807|Lupus hepatitis (disorder)
C0267807|hepatitis; lupoid
C0267807|lupoid; hepatitis
C0008312|primary biliary cirrhosis
C0008312|primary biliary cirrhosis (diagnosis)
C0008312|Biliary cirrhosis primary
C0008312|PBC
C0008312|PBC1
C0008312|BILIARY CIRRHOSIS, PRIMARY, 1
C0008312|Primary Bilary Cirrhosis (PBC)
C0008312|Chronic nonsuppurative destructive cholangitis
C0008312|Biliary cirrhosis (& [primary]) (disorder)
C0008312|Biliary cirrhosis
C0008312|Biliary cirrhosis (& [primary])
C0008312|Chronic non-suppurative destructive cholangitis
C0008312|Cholangitis, Chronic Nonsuppurative Destructive
C0008312|PBC- Primary biliary cirrhosis
C0008312|Primary biliary cirrhosis (disorder)
C0008312|biliary; cirrhosis, primary
C0008312|Hanot
C0008312|cholangitis; chronic nonsuppurative destructive
C0008312|chronic; cholangitis, chronic nonsuppurative destructive, destructive
C0008312|cirrhosis; biliary, primary
C0008312|Biliary Cirrhosis, Primary
C0008312|Cirrhosis;biliary;primary
C0850560|Other autoimmune disease
C0010346|Crohn Disease
C0010346|Crohns Disease
C0010346|Crohn's disease
C0010346|Crohn's disease [regional enteritis]
C0010346|Crohn's disease, unspecified
C0010346|INFLAMMATORY BOWEL DISEASE 1
C0010346|IBD1
C0010346|CROHN DIS
C0010346|CROHNS DIS
C0010346|eleocolitis
C0010346|enteritis (regional)
C0010346|Crohn's disease, NOS
C0010346|Crohn's disease (diagnosis)
C0010346|Crohn's ileitis
C0010346|REGIONAL ENTERITIS
C0010346|granulomatous enteritis
C0010346|Crohn's disease NOS
C0010346|Crohn Disease [Disease/Finding]
C0010346|Disease;Crohns
C0010346|Regional enteritis - Crohn's disease
C0010346|Regional enteritis - Crohn
C0010346|Crohn's regional enteritis
C0010346|Crohn's Enteritis
C0010346|-- Crohn's Disease
C0010346|Morbus Crohn
C0010346|Granulomatous enteritis and colitis
C0010346|Disease Crohns
C0010346|Crohn's
C0010346|CD - Crohn's disease
C0010346|RE - Regional enteritis
C0010346|Crohn's disease (disorder)
C0010346|Crohn
C0010346|Granulomatous enteritis, NOS
C0010346|Regional enteritis, NOS
C0678202|Regional enteritis
C0678202|regional enteritis (diagnosis)
C0678202|Regional enteritis NOS
C0678202|Enteritis;regional
C0678202|Granulomatous Enteritis
C0678202|Regional enteritis (disorder)
C0678202|Enteritis - regional
C0678202|Regional enteritis NOS (disorder)
C0678202|Granulomatous enteritis (disorder)
C0678202|Regional enteritis of unspecified site
C0678202|Enteritis, Regional
C0678202|bowel; regional enteritis
C0678202|Enteritis, Granulomatous
C1384868|disease (or disorder); autoimmune (systemic)
