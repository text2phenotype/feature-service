C0023890|Liver Cirrhosis
C0023891|Liver Cirrhosis, Alcoholic
C0023891|Alcoholic Liver Cirrhosis
C0023891|Liver Cirrhosis, Alcoholic
C0023891|Alcoholic cirrhosis of liver
C0023891|alcoholic cirrhosis
C0023891|alcoholic cirrhosis (diagnosis)
C0023891|Cirrhosis alcoholic
C0023891|Alcohol cirrhosis liver
C0023891|Alcoholic cirrhosis NOS
C0023891|Hepatic Cirrhosis, Alcoholic
C0023891|Liver Cirrhosis, Alcoholic [Disease/Finding]
C0023891|Alcoholic cirrhosis of liver (disorder)
C0023891|Laennec; alcoholic
C0023891|Laennec; cirrhosis, alcoholic
C0023891|cirrhosis; Laennec, alcoholic
C0023891|cirrhosis; alcoholic
C0023891|cirrhosis; liver, alcoholic
C0023891|liver; cirrhosis, alcoholic
C0023891|alcohol; Laennec
C0023891|alcohol; cirrhosis
C0023891|Alcoholic cirrhosis of liver (disorder) [Ambiguous]
C0023891|Alcoholic Hepatic Cirrhosis
C0023891|Laennec's cirrhosis, alcoholic
C0023891|Alcoholic cirrhosis (disorder)
C0023892|Liver Cirrhoses, Biliary
C0023892|Liver Cirrhosis, Biliary
C0023892|Cirrhosis, Biliary
C0023892|Biliary cirrhosis, unspecified
C0023892|Biliary Cirrhosis
C0023892|Cirrhosis bilary
C0023892|Biliary Liver Cirrhosis
C0023892|Liver Cirrhosis, Biliary [Disease/Finding]
C0023892|cirrhosis biliary
C0023892|biliary cirrhosis (diagnosis)
C0023892|Biliary cirrhosis NOS (disorder)
C0023892|Biliary cirrhosis NOS
C0023892|Cholangitic cirrhosis
C0023892|Cholestatic cirrhosis
C0023892|Biliary cirrhosis (disorder)
C0023892|biliary; cirrhosis
C0023892|cirrhosis; biliary
C0023892|Cirrhosis, cholangitic
C0023892|Cirrhosis, cholestatic
C0023893|Liver Cirrhosis, Experimental
C0023893|CIRRHOSES EXPER LIVER
C0023893|EXPER LIVER CIRRHOSIS
C0023893|HEPATIC CIRRHOSES EXPER
C0023893|LIVER CIRRHOSIS EXPER
C0023893|CIRRHOSIS EXPER LIVER
C0023893|EXPER LIVER CIRRHOSES
C0023893|LIVER CIRRHOSES EXPER
C0023893|Liver Cirrhosis, Experimental [Disease/Finding]
C0023893|Hepatic Cirrhosis, Experimental
C0023893|Liver Cirrhoses, Experimental
C0023893|Cirrhosis, Experimental Liver
C0023893|Experimental Liver Cirrhosis
C0023893|Cirrhoses, Experimental Liver
C0023893|Experimental Liver Cirrhoses
C0023893|Experimental Hepatic Cirrhosis
C0023890|Cirrhoses, Hepatic
C0023890|Cirrhoses, Liver
C0023890|Cirrhosis, Hepatic
C0023890|Hepatic Cirrhoses
C0023890|Liver Cirrhoses
C0023890|Liver Cirrhosis
C0023890|Cirrhosis
C0023890|Hepatic cirrhosis
C0023890|cirrhosis of liver
C0023890|hepatic cirrhosis (diagnosis)
C0023890|Cirrhosis (of liver) NOS
C0023890|Liver Cirrhosis [Disease/Finding]
C0023890|Cirrhosis, Liver
C0023890|Cirrhosis (of);liver
C0023890|Cirrhosis of liver NOS
C0023890|Cirrhosis of liver NOS (disorder)
C0023890|Liver--Cirrhosis
C0023890|Hepatic cirrhosis NOS
C0023890|Cirrhosis liver
C0023890|CL - Cirrhosis of liver
C0023890|Cirrhosis of liver (disorder)
C0023890|cirrhosis; liver
C0023890|liver; cirrhosis
C0023890|Cirrhosis of liver, NOS
C0023890|Hepatic cirrhosis, NOS
C0023890|Cirrhosis (Liver)
C0023890|cirrhosis of the liver
C0267809|CIRRHOSIS, CRYPTOGENIC
C0267809|cryptogenic cirrhosis
C0267809|cryptogenic cirrhosis (diagnosis)
C0267809|Cryptogenic cirrhosis (of liver)
C0267809|Cryptogenic cirrhosis of liver
C0267809|Cryptogenic cirrhosis (disorder)
C1442995|pigmentary cirrhosis (diagnosis)
C1442995|pigmentary cirrhosis
C1442995|Pigmentary cirrhosis (of liver)
C1442995|Bronze cirrhosis
C1442995|Pigmentary cirrhosis of liver
C1442995|Bronzed cirrhosis
C1442995|Bronze cirrhosis (disorder)
C2004456|postnecrotic cirrhosis (diagnosis)
C2004456|postnecrotic cirrhosis
C2004456|macronodular cirrhosis
C2004456|macronodular cirrhosis (diagnosis)
C2004456|Macronodular cirrhosis (of liver)
C2004456|Postnecrotic cirrhosis (of liver)
C2004456|Postnecrotic cirrhosis of liver
C2004456|Hypertrophic portal cirrhosis
C2004456|Macronodular cirrhosis of liver
C2004456|PNC - Postnecrotic cirrhosis
C2004456|Macronodular cirrhosis (disorder)
C2004456|Cirrhosis liver postnecrotic
C2004456|Hepatic cirrhosis post necrotic
C2004456|Cirrhosis liver post necrotic
C2004456|Healed yellow atrophy of liver
C2004456|Postnecrotic cirrhosis (disorder)
C2004456|cirrhosis; macronodular
C2004456|cirrhosis; periportal
C2004456|cirrhosis; postnecrotic
C2004456|macronodular; cirrhosis
C2004456|periportal; cirrhosis
C2004456|postnecrotic; cirrhosis
C0267812|Micronodular cirrhosis
C0267812|micronodular cirrhosis (diagnosis)
C0267812|Micronodular cirrhosis (disorder)
C0267812|cirrhosis; micronodular
C0267812|micronodular; cirrhosis
C0085699|Cardiac cirrhosis
C0085699|cardiac cirrhosis (diagnosis)
C0085699|Congestive cirrhosis
C0085699|Cardiac cirrhosis (disorder)
C0085699|cardiac; cirrhosis
C0085699|cirrhose cardiaque
C0085699|cirrhosis; cardiac
C0085699|cirrhosis; congestive
C0085699|congestive; cirrhosis
C0085699|Cardiac cirrhosis, NOS
C2062319|cirrhosis, rare types
C2062319|rare types of cirrhosis
C2062319|rare types of cirrhosis (diagnosis)
C2075269|cirrhosis due to hepatitis A
C2075269|cirrhosis due to hepatitis A (diagnosis)
C2075270|cirrhosis due to hepatitis B
C2075270|cirrhosis due to hepatitis B (diagnosis)
C2075271|cirrhosis due to hepatitis C (diagnosis)
C2075271|cirrhosis due to hepatitis C
C0154307|idiopathic portal hypertension
C0154307|idiopathic portal hypertension (diagnosis)
C0154307|Banti's disease
C0154307|Idiopathic congestive splenomegaly
C0154307|Banti's syndrome
C0154307|Fibrocongestive splenomegaly
C0154307|Banti syndrome
C0154307|Banti's spleen
C0154307|Congestive splenomegaly
C0154307|Congestive splenomegaly (disorder)
C0154307|Banti
C1622502|Portal cirrhosis (of liver)
C1622502|Portal cirrhosis unspecified
C1622502|Laennec's cirrhosis
C1622502|Portal cirrhosis
C1622502|Portal cirrhosis (disorder)
C1622502|Portal cirrhosis unspecified (disorder)
C1622502|PC - Portal cirrhosis
C1622502|cirrhosis portal
C1622502|Portal cirrhosis (diagnosis)
C1622502|Laennec; cirrhosis
C1622502|Laennec
C1622502|cirrhosis; Laennec
C1622502|cirrhosis; portal
C1622502|portal; cirrhosis
C1622502|Portal cirrhosis, NOS
C0400947|cirrhosis diffuse nodular
C0400947|cirrhosis diffuse nodular (diagnosis)
C0400947|Diffuse nodular cirrhosis
C0400947|Diffuse nodular cirrhosis (disorder)
C0400951|cirrhosis cardituberculous (diagnosis)
C0400951|cirrhosis cardituberculous
C0400951|Cardituberculous cirrhosis
C0400951|Cardituberculous cirrhosis (disorder)
C0268074|INDIAN CHILDHOOD CIRRHOSIS
C0268074|CIRRHOSIS, FAMILIAL, WITH PULMONARY HYPERTENSION
C0268074|ICC
C0268074|SEN SYNDROME
C0268074|Cirrhosis-familial with pulmonary hypertension
C0268074|ICC - Indian childhood cirrhosis
C0268074|Indian childhood cirrhosis (disorder)
C0268074|Indian childhood; cirrhosis
C0268074|cirrhosis; Indian childhood
C1392670|Congenital cirrhosis (of liver)
C1392670|congenital cirrhosis liver
C1392670|congenital cirrhosis of liver
C1392670|congenital cirrhosis of liver (diagnosis)
C1392670|cirrhosis; liver, congenital
C0239946|Fibroses, Liver
C0239946|Liver Fibroses
C0239946|Hepatic fibrosis
C0239946|hepatic fibrosis (diagnosis)
C0239946|Liver fibrosis
C0239946|Fibrosis of liver
C0239946|Fibrosis of liver (disorder)
C0239946|Fibrosis liver
C0239946|Hepatic fibrosis (disorder)
C0239946|fibrosis; liver
C0239946|liver; fibrosis
C0239946|Hepatic fibrosis, NOS
C0239946|Fibrosis, Liver
C3662136|Chronic hepatitis C with stage 4 fibrosis
C3662136|Cirrhosis of liver due to chronic hepatits C (disorder)
C3662136|Cirrhosis of liver due to chronic hepatits C
C3662136|Cirrhosis of liver due to chronic hepatitis C
C3662136|Cirrhosis of liver due to chronic hepatitis C (disorder)
C0275872|Syphilitic cirrhosis
C0275872|cirrhosis syphilitic
C0275872|Syphilitic cirrhosis (diagnosis)
C0275872|Hepar lobatum
C0275872|Syphilitic cirrhosis (disorder)
C1861556|CIRRHOSIS, FAMILIAL
C0009714|Congenital hepatic fibrosis
C0009714|HEPATIC FIBROSIS, CONGENITAL
C0009714|congenital hepatic fibrosis (diagnosis)
C0009714|Congenital Fibrose Liver
C0009714|Congenital hepatic fibrosis (disorder)
C1859088|COPPER TOXICOSIS, IDIOPATHIC
C1859088|ICT
C3874483|Cirrhosis of liver due to hepatitis B (disorder)
C3874483|Cirrhosis of liver due to hepatitis B
C1392669|Mixed cirrhosis
C1392669|cirrhosis; mixed type
C1392669|mixed; cirrhosis
C0010398|Cruveilhier Baumgarten Syndrome
C0010398|Syndrome, Cruveilhier-Baumgarten
C0010398|Cruveilhier-Baumgarten syndrome
C0010398|Cruveilhier-Baumgarten syndrome (disorder)
C0010398|cirrhosis; Baumgarten-Cruveilhier
C0010398|cirrhosis; Cruveilhier-Baumgarten
C0010398|Baumgarten-Cruveilhier; cirrhosis
C0010398|Baumgarten-Cruveilhier
C0010398|Cruveilhier-Baumgarten; cirrhosis
C0010398|Cruveilhier-Baumgarten
C0267806|Florid cirrhosis
C0267806|Florid cirrhosis (disorder)
C0267817|Glissonian cirrhosis
C0267817|Glissonian cirrhosis (disorder)
C0267815|Pigment cirrhosis
C0267815|Pigment cirrhosis (disorder)
C0267813|Posthepatitic cirrhosis
C0267813|Posthepatitic cirrhosis (disorder)
C0267813|cirrhosis; posthepatitic
C0267813|posthepatitic; cirrhosis
C0156189|Chronic liver disease and cirrhosis
C0156189|Cirrhosis/chronic liver dis.
C0156189|Cirrhosis and chronic liver disease
C0156189|Cirrhosis and chronic liver disease (disorder)
C0341446|Hepatic sclerosis
C0341446|hepatic sclerosis (diagnosis)
C0341446|Hepatic sclerosis (disorder)
C0341446|liver; sclerosis
C0341446|sclerosis; liver
C0348749|Other and unspecified cirrhosis of liver
C0348749|[X]Other and unspecified cirrhosis of liver (disorder)
C0348749|[X]Other and unspecified cirrhosis of liver
C0400941|portal cirrhosis capsular (diagnosis)
C0400941|portal cirrhosis capsular
C0400941|Capsular portal cirrhosis
C0400941|Capsular portal cirrhosis (disorder)
C0400957|Cirrhosis secondary to cholestasis (disorder)
C0400957|Cirrhosis secondary to cholestasis
C0400942|portal cirrhosis fatty
C0400942|portal cirrhosis fatty (diagnosis)
C0400942|Fatty portal cirrhosis
C0400942|Fatty portal cirrhosis (disorder)
C0400961|Hepatic fibrosis with hepatic sclerosis
C0400961|hepatic fibrosis with hepatic sclerosis (diagnosis)
C0400961|Hepatic fibrosis with hepatic sclerosis (disorder)
C0400961|fibrosis; liver, with sclerosis
C0400961|sclerosis; liver, with fibrosis
C0400949|Infectious cirrhosis NOS (disorder)
C0400949|Infectious cirrhosis NOS
C0400949|Infectious cirrhosis
C0400949|Infectious cirrhosis (disorder)
C0400940|Pigmentary portal cirrhosis
C0400940|Pigmentary portal cirrhosis (disorder)
C0400956|Toxic cirrhosis
C0400956|Toxic cirrhosis (disorder)
C0400939|portal cirrhosis toxic (diagnosis)
C0400939|portal cirrhosis toxic
C0400939|Toxic portal cirrhosis
C0400939|Toxic portal cirrhosis (disorder)
C0400938|portal cirrhosis unilobular (diagnosis)
C0400938|portal cirrhosis unilobular
C0400938|Unilobular portal cirrhosis
C0400938|Unilobular portal cirrhosis (disorder)
C0400943|Cirrhosis, nonalcoholic
C0400943|Non-alcoholic cirrhosis NOS
C0400943|Cirrhosis - non alcoholic
C0400943|Cirrhosis - non-alcoholic
C0400943|Cirrhosis - non-alcoholic (disorder)
C0400943|Non-alcoholic cirrhosis NOS (disorder)
C0400943|Cirrhosis of liver not due to alcohol
C0400943|Cirrhosis of liver not due to alcohol (disorder)
C0400955|Hypoxia-associated cirrhosis
C0400955|Hypoxia-associated cirrhosis (disorder)
C1263668|Cholangiolitic cirrhosis (disorder)
C1263668|Cholangiolitic cirrhosis
C1263668|cholangiolitic; cirrhosis
C1263668|cirrhosis; cholangiolitic
C1299579|Early cirrhosis (disorder)
C1299579|Early cirrhosis
C1263666|Advanced cirrhosis (disorder)
C1263666|Advanced cirrhosis
C1263665|Latent cirrhosis (disorder)
C1263665|Latent cirrhosis
C1263663|Nutritional cirrhosis (disorder)
C1263663|Nutritional cirrhosis
C1263663|cirrhosis; nutritional
C1263663|nutritional; cirrhosis
C0008312|primary biliary cirrhosis
C0008312|primary biliary cirrhosis (diagnosis)
C0008312|Biliary cirrhosis primary
C0008312|PBC
C0008312|PBC1
C0008312|BILIARY CIRRHOSIS, PRIMARY, 1
C0008312|Primary Bilary Cirrhosis (PBC)
C0008312|Chronic nonsuppurative destructive cholangitis
C0008312|Biliary cirrhosis (& [primary]) (disorder)
C0008312|Biliary cirrhosis
C0008312|Biliary cirrhosis (& [primary])
C0008312|Chronic non-suppurative destructive cholangitis
C0008312|Cholangitis, Chronic Nonsuppurative Destructive
C0008312|PBC- Primary biliary cirrhosis
C0008312|Primary biliary cirrhosis (disorder)
C0008312|biliary; cirrhosis, primary
C0008312|Hanot
C0008312|cholangitis; chronic nonsuppurative destructive
C0008312|chronic; cholangitis, chronic nonsuppurative destructive, destructive
C0008312|cirrhosis; biliary, primary
C0008312|Biliary Cirrhosis, Primary
C0008312|Cirrhosis;biliary;primary
C0238065|Obstructive Liver Cirrhosis
C0238065|Secondary biliary cirrhosis
C0238065|secondary biliary cirrhosis (diagnosis)
C0238065|Biliary cirrhosis secondary
C0238065|Liver Cirrhosis, Obstructive
C0238065|Cirrhosis, Secondary Biliary
C0238065|Secondary biliary cirrhosis (disorder)
C0238065|cirrhosis; biliary, secondary
C0238065|Biliary Cirrhosis, Secondary
C0400935|Juvenile portal cirrhosis
C0400935|Childhood function cirrhosis
C0400935|Juvenile portal cirrhosis (disorder)
C1960179|Drug-induced cirrhosis of liver (disorder)
C1960179|Drug-induced hepatic cirrhosis
C1960179|Drug-induced cirrhosis of liver
C0400925|Alcoholic fibrosis and sclerosis of liver
C0400925|alcoholic sclerosis and fibrosis of liver (diagnosis)
C0400925|alcoholic sclerosis and fibrosis of liver
C0400925|Alcoholic fibrosis and sclerosis of liver (disorder)
C2887912|Alcoholic cirrhosis of liver without ascites
C2887913|Alcoholic cirrhosis of liver with ascites
C3509286|cirrhosis alcoholic (laennec's) with ascites
C3509286|alcoholic cirrhosis with ascites
C3509286|alcoholic cirrhosis with ascites (diagnosis)
C3838604|alcoholic cirrhosis without ascites
C3838604|alcoholic cirrhosis without ascites (diagnosis)
C3838604|cirrhosis alcoholic (laennec's) without ascites
C3838604|alcoholic (Laennec's) cirrhosis without ascites
C1392672|cirrhosis; macronodular, alcoholic
C1392672|macronodular; cirrhosis, alcoholic
C1392673|cirrhosis; micronodular, alcoholic
C1392673|micronodular; cirrhosis, alcoholic
C1392676|cirrhosis; portal, alcoholic
C1392676|portal; cirrhosis, alcoholic
C1392677|cirrhosis; postnecrotic, alcoholic
C1392677|postnecrotic; cirrhosis, alcoholic
C1392681|cirrhosis; nutritional, alcohol
C1392681|nutritional; cirrhosis, alcohol
