C0421451|Patient date of birth
C2967445|Birth date patient
C2348576|Subject Birth Date
C2919018|Birth Date and Time
C2348576|Subject Birth Date
C2986369|Biologic Entity Birth Date
C2986369|BiologicEntity.birthDate
C0421451|Patient date of birth
C0421451|BD
C0421451|DOB
C0421451|Date of Birth
C0421451|Birth Date
C0421451|Date of birth (finding)
C0421451|BRTHDAT
C0421451|birthDate
C0421451|DOB - Date of birth
C0421451|Date of birth (observable entity)
C0421451|Date of birth of person cared for
C0421451|Date of birth of recipient of care (observable entity)
C0421451|Date of birth of recipient of care
C2967445|Birth date &#x7C; patient
C0803906|Birth date:Time Stamp -- Date and Time:Point in time:^Patient:Quantitative
C0803906|Birth date
C0803906|Birth date:TmStp:Pt:^Patient:Qn
