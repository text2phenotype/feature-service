C1849687|Liver biopsy shows normal numbers of enlarged peroxisomes
C1856310|Liver biopsy shows diffuse interstitial fibrosis
C1857356|Liver biopsy shows increased lipid droplets (microvesicular steatosis)
C1857367|Liver biopsy shows increased lipid droplets and abnormal mitochondria
C2021366|liver biopsy iron (ug/100 mg of dry weight)
C2121176|liver biopsy when done for indicated purpose at time of other major procedure
C2368138|hepatic cyst aspiration for echinococcus identification
C2674614|Liver biopsy shows red autofluorescence and needle-like cytoplasmic inclusion bodies
C2748696|Liver biopsy shows ductal proliferation
C2751577|Liver biopsy during acute episode shows variable portal and sinusoidal fibrosis
C3277942|Liver biopsy shows portal and/or bridging fibrosis
C4273160|bile duct biopsy showed paucity of ducts    
C3899974|BCLC Stage
C3897124|BCLC Stage A Hepatocellular Carcinoma
C3897124|BCLC Stage A
C3898888|HCC by BCLC Stage
C3898888|BCLC Hepatocellular Carcinoma
C3898888|BCLC Stage Hepatocellular Carcinoma
C3898888|Hepatocellular Carcinoma by BCLC Stage
C3899975|BCLC Stage D Hepatocellular Carcinoma
C3899975|BCLC Stage D HCC
C3899977|BCLC Stage C Hepatocellular Carcinoma
C3899975|BCLC Stage C HCC
C3899979|BCLC Stage B Hepatocellular Carcinoma
C3899975|BCLC Stage B HCC
C3899981|BCLC Stage A Adult Hepatocellular Carcinoma
C3899975|BCLC Stage A HCC
C3899982|BCLC Stage 0 Hepatocellular Carcinoma
C3899975|BCLC Stage 0 HCC
C3899976|BCLC Stage D Adult Hepatocellular Carcinoma
C3899976|BCLC Stage D Adult HCC
C3899978|BCLC Stage C Adult Hepatocellular Carcinoma
C3899978|BCLC Stage C Adult HCC
C3899980|BCLC Stage B Adult Hepatocellular Carcinoma
C3899980|BCLC Stage B Adult HCC
C3899983|BCLC Stage 0 Adult Hepatocellular Carcinoma
C3899983|BCLC Stage 0 Adult HCC
C3550399|Increased iron deposition seen on liver biopsy
C4020697|Giant cell hepatitis on liver biopsy
C4314030|Ductal reaction seen on liver biopsy
C1847706|Absence of beta-ureidopropionase activity and protein in liver biopsy
C3899981|Barcelona Clinic Liver Cancer Stage A Adult Hepatocellular Carcinoma
C3899981|BCLC Stage A Adult Hepatocellular Carcinoma
C3899982|BCLC Stage 0 Hepatocellular Carcinoma
C3899982|Barcelona Clinic Liver Cancer Stage 0 Hepatocellular Carcinoma
C3897124|Barcelona Clinic Liver Cancer Stage A Hepatocellular Carcinoma
C3897124|BCLC Stage A Hepatocellular Carcinoma
C3899975|BCLC Stage D Hepatocellular Carcinoma
C3899975|Barcelona Clinic Liver Cancer Stage D Hepatocellular Carcinoma
C3899977|Barcelona Clinic Liver Cancer Stage C Hepatocellular Carcinoma
C3899977|BCLC Stage C Hepatocellular Carcinoma
C3899979|BCLC Stage B Hepatocellular Carcinoma
C3899979|Barcelona Clinic Liver Cancer Stage B Hepatocellular Carcinoma
C3899976|Barcelona Clinic Liver Cancer Stage D Adult Hepatocellular Carcinoma
C3899976|BCLC Stage D Adult Hepatocellular Carcinoma
C3899978|Barcelona Clinic Liver Cancer Stage C Adult Hepatocellular Carcinoma
C3899978|BCLC Stage C Adult Hepatocellular Carcinoma
C3899980|BCLC Stage B Adult Hepatocellular Carcinoma
C3899980|Barcelona Clinic Liver Cancer Stage B Adult Hepatocellular Carcinoma
C3899983|Barcelona Clinic Liver Cancer Stage 0 Adult Hepatocellular Carcinoma
C3899983|BCLC Stage 0 Adult Hepatocellular Carcinoma
