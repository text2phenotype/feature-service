C0474232|patient immune to hepatitis B
C0474232|patient immune to Hep B
C0474232|patient vaccinated for Hep B
C0474232|Hepatitis B vaccination (SNOMED:16584000)
C2716397|Diphtheria and Tetanus Toxoids and Acellular Pertussis Adsorbed, Inactivated Poliovirus, Haemophilus b Conjugate (Meningococcal Protein Conjugate), and Hepatitis B (Recombinant) Vaccine. 
C2716397|DTaP,IPV,Hib,HepB                                                                                     
C3644155|DTaP-Hep B-IPV                                                                                       
C3644155|DTaP-hepatitis B and poliovirus vaccine                                                                          
C3644182|DTaP-IPV-HIB-HEP B, historical                                                                               
C1548467|DTaP/DTP-Hib-Hep B                                                                                     
C1548467|DTP- Haemophilus influenzae type b conjugate and hepatitis b vaccine                                                            
C0694743|Haemophilus influenzae type b conjugate and Hepatitis B vaccine
C0694733|Hep B, adolescent or pediatric                                                                               
C1552908|Hep B, adolescent/high risk infant                                                                             
C1552909|Hep B, adult                                                                                        
C0694736|Hep B, dialysis                                                                                      
C3644158|Hep B, unspecified formulation
C0062525|hepatitis B immune globulin                                                                                
C1552908|hepatitis B vaccine, adolescent/high risk infant dosage                                                                  
C1552909|hepatitis B vaccine, adult dosage                                                                             
C0694736|hepatitis B vaccine, dialysis patient dosage                                                                       
C0694733|hepatitis B vaccine, pediatric or pediatric/adolescent dosage                                                              
C3644158|hepatitis B vaccine, unspecified formulation
C0694743|Hib-Hep B                                                                                         
C3644182|Historical record of vaccine containing * diphtheria, tetanus toxoids and acellular pertussis, * poliovirus, inactivated, * Haemophilus influenzae type b conjugate, * Hepatitis B     
C1170008|Hep A-Hep B                                                                                        
C0730242|combined hepatitis a & hepatitis b vaccination
C0730242|combined hepatitis A and hepatitis B vaccination (medication)
C0730242|combined hepatitis A and hepatitis B vaccination
C0730242|Combined hepatitis A and B vaccination
C0730242|Combined hepatitis A and B vaccination (procedure)
C1300747|vacc comb bact & viral administered diphth - acell pertus - hepb - ipv
C1300747|diphtheria-acellular pertussis-hepB-IPV vaccination
C1300747|diphtheria-acellular pertussis-hepB-IPV vaccination (medication)
C1300747|Diphtheria, acellular pertussis, hepatitis B and inactivated polio vaccination (procedure)
C1300747|Diphtheria, acellular pertussis, hepatitis B and inactivated polio vaccination
C0474232|Hepatitis B immunisation
C0474232|Immunisation;hepatitis B
C0474232|Hepatitis B immunization
C0474232|Hepatitis b vaccine (active) administration
C0474232|Hepatitis b vaccine administration (medication)
C0474232|Hepatitis b vaccine administration
C0474232|Administration of hepatitis b vaccine
C0474232|Hep B vaccination
C0474232|Hepatitis B series immunization
C0474232|Hepatitis B vaccination
C0474232|Hepatitis B injection
C0474232|Hepatitis B series immunisation
C0474232|Hepatitis B vaccination (procedure)
C0474232|Admin hepatitis b vaccine
C0474232|Immunization;hepatitis B
C0419731|Booster hepatitis B vaccination (procedure)
C0419731|Booster hepatitis B vaccination
C0419731|hepatitis b vaccine (active) booster vaccination (medication)
C0419731|hepatitis b vaccine (active) booster vaccination
C0419729|Fourth hepatitis B vaccination (procedure)
C0419729|Fourth hepatitis B vaccination
C0419729|hepatitis b vaccine (active) fourth vaccination
C0419729|hepatitis b vaccine (active) fourth vaccination (medication)
C0419729|4th hepatitis B vaccination
C0419727|Second hepatitis B vaccination (procedure)
C0419727|Second hepatitis B vaccination
C0419727|hepatitis b vaccine (active) second vaccination
C0419727|hepatitis b vaccine (active) second vaccination (medication)
C0419727|2nd hepatitis B vaccination
C0419728|Third hepatitis B vaccination (procedure)
C0419728|Third hepatitis B vaccination
C0419728|hepatitis b vaccine (active) third vaccination
C0419728|hepatitis b vaccine (active) third vaccination (medication)
C0419728|3rd hepatitis B vaccination
C0419726|First hepatitis B vaccination
C0419726|First hepatitis B vaccination (procedure)
C0419726|hepatitis b vaccine (active) first vaccination
C0419726|hepatitis b vaccine (active) first vaccination (medication)
C0419726|1st hepatitis B vaccination
C0419730|Fifth hepatitis B vaccination
C0419730|Fifth hepatitis B vaccination (procedure)
C0419730|5th hepatitis B vaccination
C1293866|intramuscular injection of hepatitis B immune globulin (human)
C1293866|globulin, hepatitis b immune (human) intramuscular injection
C1293866|intramuscular injection of hepatitis B immune globulin (human) (medication)
C1293866|Hepatitis B Virus immune globulin administration by intramuscular injection
C1293866|Intramuscular injection of Hepatitis B Virus immune globulin, human (procedure)
C1293866|Intramuscular injection of Hepatitis B Virus immune globulin, human
C1562257|Sixth hepatitis B vaccination (procedure)
C1562257|Sixth hepatitis B vaccination
C3661302|Infanrix hexa
C2716397|diphtheria-tetanus-acellular pertussis-inactivated poliovirus-Haemophilus influenzae b conjugate-hepatitis B vaccine
C2716397|DTaP-IPV-Hib-HBV vaccine
C2716397|DTaP-IPV-Hib-HBV conjugate vaccine
C2716397|dtap-ipv-hib-hepb
C2716397|dtap-ipv-hib-hepb (medication)
C2716397|DTaP,IPV,Hib,HepB
C2716397|Diphtheria and Tetanus Toxoids and Acellular Pertussis Adsorbed, Inactivated Poliovirus, Haemophilus b Conjugate (Meningococcal Protein Conjugate), and Hepatitis B (Recombinant) Vaccine.
C3644155|DTaP-Hep B-IPV
C3644155|DTaP-hepatitis B and poliovirus vaccine
C3644182|Historical record of vaccine containing * diphtheria, tetanus toxoids and acellular pertussis, * poliovirus, inactivated, * Haemophilus influenzae type b conjugate, * Hepatitis B
C3644182|DTaP-IPV-HIB-HEP B, historical
C1548467|DTaP/DTP-Hib-Hep B
C1548467|DTP- Haemophilus influenzae type b conjugate and hepatitis b vaccine
C1548467|DTP-Hib-Hep B
C0694743|Hib-Hep B
C0694743|Haemophilus influenzae type b conjugate and Hepatitis B vaccine
C0694733|hepatitis B vaccine, pediatric or pediatric/adolescent dosage
C0694733|Hep B, adolescent or pediatric
C1552908|hepatitis B vaccine, adolescent/high risk infant dosage
C1552908|Hep B, adolescent/high risk infant
C1552909|hepatitis B vaccine, adult dosage
C1552909|Hep B, adult
C0694736|Hep B, dialysis
C0694736|hepatitis B vaccine, dialysis patient dosage
C3644158|Hep B, unspecified formulation
C3644158|hepatitis B vaccine, unspecified formulation
C0720993|Hyperhep
C0703267|hepatitis B immune globulin intramuscular solution
C0720796|H-BIG
C0718838|Bayhep B
C1725338|HepaGam B
C0062525|HBIG
C0062525|hepatitis B hyperimmune globulin
C0062525|Hepatitis B immunoglobulin
C0062525|globulin, hepatitis B immune (human)
C0062525|globulin, hepatitis B immune (human) for intramuscular use
C0062525|hepatitis B immune globulin
C0062525|human hepatitis B immune globulin for intramuscular use (medication)
C0062525|human hepatitis B immune globulin
C0062525|human hepatitis B immune globulin for intramuscular use
C0062525|human hepatitis B immune globulin (medication)
C0062525|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN
C0062525|hepatitis B hyperimmune globulin [Chemical/Ingredient]
C0062525|HEPATITIS B IMMUNE GLOBULIN,HUMAN
C0062525|Anti-Hepatitis B immunoglob.
C0062525|Hepatitis B immunoglobulin (substance)
C0062525|Antihepatitis B immunoglobulin
C0062525|Hepatitis B immune globulin (human)
C0062525|Hepatitis B immune globulin (human) (product)
C0062525|Hepatitis B immune globulin (human) (substance)
C1700143|Hyperhep B
C3888170|HEPATITIS B NABI-HB GLOBULIN INJ VIL 1ML
C3888170|HUMAN HEPATITIS B VIRUS IMMUNE GLOBULIN 312 [iU] in 1 mL INTRAMUSCULAR INJECTION [NABI-HB]
C3888170|Nabi-HB 312unit/ml Solution for Injection
C3888170|HEPATITIS B IMMUNE GLOBULIN (NABI-HB) INJ,VIL,1ML
C3888170|HEPATITIS B IMMUNE GLOBULIN (NABI-HB) INJ,VIL,1ML [VA Product]
C3888170|Hepatitis B Immune Globulin Intramuscular Solution [NABI-HB NOVAPLUS]
C3888170|1 ML hepatitis B immune globulin 312 UNT/ML Injection [Nabi-HB]
C3888170|1 ML Nabi-HB 312 UNT/ML Injection
C3888170|Nabi-HB > 312 UNT/ML in 1 ML Injection
C3888170|Hepatitis B Immune Globulin Intramuscular Solution [NABI-HB]_#1
C3888170|Nabi-HB, intramuscular solution_#1
C1815761|HEPATITIS B IMMUNE GLOBULIN (BAYHEP) INJ,SYR,1ML
C1815761|HEPATITIS B GLOBULIN (BAYHEP) INJ 1ML
C1815761|1 ML Bayhep B 217 UNT/ML Prefilled Syringe
C1815761|1 ML hepatitis B immune globulin 217 UNT/ML Prefilled Syringe [Bayhep B]
C1815761|Bayhep B 217 UNT per 1 ML Prefilled Syringe
C1815761|HEPATITIS B IMMUNE GLOBULIN (BAYHEP) INJ,SYR,1ML [VA Product]
C0709015|Bayhep B 217 UNT/ML Injectable Solution
C0709015|HEPATITIS B IMMUNE GLOBULIN (BAYHEP) INJ
C0709015|hepatitis B immune globulin 217 UNT/ML Injectable Solution [Bayhep B]
C0709015|BayHep B 217unit/ml Solution for Injection
C0709015|HEPATITIS B IMMUNE GLOBULIN (BAYHEP) INJ [VA Product]
C2937711|Hepatitis B Immune Globulin Injection Solution
C0353106|Anti-hbs immunoglobulin injection
C0353106|Anti-hbs immunoglobulin injection (product)
C0353106|Anti-hbs immunoglobulin injection (substance)
C0590210|Hepatitis B immunoglobulin 1000iu injection
C0590210|Hepatitis B immunoglobulin 1000iu powder for injection solution vial (product)
C0590210|Hepatitis B immunoglobulin 1000iu powder for injection solution vial
C0590210|Hepatitis B immunoglobulin 1000iu injection (product)
C0590210|Hepatitis B immunoglobulin 1000iu injection (substance)
C0590211|Hepatitis B immunoglobulin 200iu injection
C0590211|Hepatitis B immunoglobulin 200iu powder for injection solution vial (product)
C0590211|Hepatitis B immunoglobulin 200iu powder for injection solution vial
C0590211|Hepatitis B immunoglobulin 200iu injection (product)
C0590211|Hepatitis B immunoglobulin 200iu injection (substance)
C0590212|Hepatitis B immunoglobulin 500iu injection
C0590212|Hepatitis B immunoglobulin 500iu powder for injection solution vial (product)
C0590212|Hepatitis B immunoglobulin 500iu powder for injection solution vial
C0590212|Hepatitis B immunoglobulin 500iu injection (product)
C0590212|Hepatitis B immunoglobulin 500iu injection (substance)
C1298253|Hepatitis b immune globulin 1unt/vial (product)
C1298253|Hepatitis b immune globulin 1unt/vial
C1163957|Hepatitis b immune globulin 217u injection solution vial (product)
C1163957|Hepatitis b immune globulin 217u injection solution vial
C1163957|Hepatitis b immune globulin 217unt injection
C1163957|Hepatitis b immune globulin 217unt injection (product)
C0876102|Nabi-HB
C0876102|Nabi-HB Novaplus
C3888113|Hepatitis b immune globulin 312units/mL injection solution 5mL vial (product)
C3888113|Hepatitis b immune globulin 312units/mL injection solution 5mL vial
C3888113|Hepatitis B Immune Globulin (Human) 1560U Solution for injection
C3888113|hepatitis B immune globulin (human) > 312 UNT/ML in 5 ML Injection
C3888113|5 ML hepatitis B immune globulin 312 UNT/ML Injection
C1948568|Hepatitis b immune globulin 312units/mL injection solution 1mL vial (product)
C1948568|Hepatitis b immune globulin 312units/mL injection solution 1mL vial
C1948568|hepatitis B immune globulin injectable solution
C1948568|Hepatitis B Immune Globulin (Human) 312U/1mL Solution for injection
C1948568|hepatitis B immune globulin (human) > 312 UNT/ML in 1 ML Injection
C1948568|1 ML hepatitis B immune globulin 312 UNT/ML Injection
C1170689|Twinrix Junior
C1170008|Hepatitis A and hepatitis B vaccine
C1170008|Hep A-Hep B
C1170008|hepatitis A-hepatitis B vaccine
