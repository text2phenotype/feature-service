C0005437|Bilirubin
C0201913|Bilirubin, total measurement
C0863174|Blood bilirubin measurement
C0053592|21H-biline-8,12-dipropanoic acid, 2,17-diethenyl-1,10-19,22,23,24-hexahydro-3,7,13,18-tetramethyl-1,19-dioxo-, mono-beta-D-glucopyranuronosyl ester
C0053592|bilirubin glucuronate
C0053592|bilirubin glucuronide
C0053592|bilirubin, glucuronic acid conjugates
C0053592|Bilirubin glucuronide (substance)
C0236556|Direct reacting bilirubin
C0236556|Direct (Conjugated) Bilirubin
C0236556|Conjugated bilirubin
C0236556|Split bilirubin
C0236556|Direct bilirubin
C0236556|CB - Conjugated bilirubin
C0236556|DB - Direct bilirubin
C0236556|Direct reacting bilirubin (substance)
C0236556|Direct reacting bilirubin, NOS
C0301719|Indirect reacting bilirubin
C0301719|Indirect (Unconjugated) Bilirubin
C0301719|Unconjugated bilirubin
C0301719|Indirect bilirubin
C0301719|BU - Bilirubin
C0301719|UCB - Unconjugated bilirubin
C0301719|UCBR - Unconjugated bilirubin
C0301719|Indirect reacting bilirubin (substance)
C0005446|Biliverdine
C0005446|21H-Biline-8,12-dipropanoic acid, 3,18-diethenyl-1,19,22,24-tetrahydro-2,7,13,17-tetramethyl-1,19-dioxo-
C0005446|Biliverdin
C0005446|Ooecyan
C0005446|Biliverdine [Chemical/Ingredient]
C0005446|Dehydrobilirubin
C0005446|Uteroverdine
C0005446|Biliverdin (substance)
C0005437|Bilirubin, total
C0005437|Bilirubin
C0005437|21H-Biline-8,12-dipropanoic acid, 2,17-diethenyl-1,10,19,22,23,24-hexahydro-3,7,13,18-tetramethyl-1,19-dioxo-
C0005437|Bilirubin [Chemical/Ingredient]
C0005437|Bilirubin IX alpha
C0005437|Conjugated and unconjugated bilirubin
C0005437|Bilirubin (substance)
C0005437|Bilirubin, NOS
C0005437|Total bilirubin
C0887593|Bilirubin, (15E)-Isomer
C0887594|Bilirubin, (4E)-Isomer
C0887595|Bilirubin, (4E,15E)-Isomer
C0368752|Bilirubin.non-glucuronidated
C1982584|Bilirubin &#x7C; gastric fluid
C3262266|Bilirubin.total [Moles/volume] in Urine by Automated test strip
C3262266|Bilirubin:SCnc:Pt:Urine:Qn:Test strip.automated
C3262266|Bilirub Ur Strip.auto-sCnc
C3262266|Bilirubin:Substance Concentration:Point in time:Urine:Quantitative:Test strip.automated
C1982580|Bilirubin &#x7C; body fluid
C2924724|Bilirubin &#x7C; Blood arterial
C1982593|Bilirubin &#x7C; XXX
C0017776|Glucuronidase
C0017776|beta glucuronidase
C0017776|beta-D-Glucuronoside glucuronosohydrolase
C0017776|Beta-glucuronidase
C0017776|Glucuronidase [Chemical/Ingredient]
C0017776|Beta-glucuronidase (substance)
C0803316|Bilirubin:MCnc:Pt:Urine:Qn:Test strip
C0803316|Bilirub Ur Strip-mCnc
C0803316|Bilirubin:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C0803316|Bilirubin.total [Mass/volume] in Urine by Test strip
C0367985|Bilirubin:ACnc:Pt:Urine:Ord:Test strip
C0367985|Bilirub Ur Ql Strip
C0367985|Bilirubin:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0367985|Bilirubin.total [Presence] in Urine by Test strip
C1982578|Bilirubin &#x7C; bld-ser-plas
C2925975|Bilirubin [Presence] in Urine by Confirmatory method
C2925975|Bilirub Ur Ql Cfm
C2925975|Bilirubin:Threshold:Point in time:Urine:Ordinal:Confirm
C2925975|Bilirubin:Threshold:Pt:Urine:Ord:Confirm
C3534268|Bilirubin excess &#x7C; Bld-Ser-Plas
C3700088|Bilirubin &#x7C; Calculus (stone)
C1982590|Bilirubin &#x7C; synovial fluid
C1982585|Bilirubin &#x7C; Pericardial fluid
C0805304|Bilirubin.glucuronidated
C2924726|Bilirubin &#x7C; Blood venous
C1982600|Bilirubin.albumin bound &#x7C; bld-ser-plas
C1982577|Bilirubin &#x7C; amniotic fluid
C1715313|Bilirubin:ACnc:24H:Urine:Ord:Test strip
C1715313|Bilirubin:Arbitrary Concentration:24 hours:Urine:Ordinal:Test strip
C1715313|Bilirubin.total [Presence] in 24 hour Urine by Test strip
C1715313|Bilirub 24h Ur Ql Strip
C1982589|Bilirubin &#x7C; stool
C2361847|Bilirubin:MCnc:Pt:Urine:Qn:Test strip.automated
C2361847|Bilirub Ur Strip.auto-mCnc
C2361847|Bilirubin:Mass Concentration:Point in time:Urine:Quantitative:Test strip.automated
C2361847|Bilirubin.total [Mass/volume] in Urine by Automated test strip
C1982592|Bilirubin &#x7C; Urine and Serum or Plasma
C1982586|Bilirubin &#124; peritoneal fluid
C1982586|Bilirubin &#x7C; peritoneal fluid
C1991615|Liley Zone &#x7C; Amniotic Fluid
C1544963|Bilirub Ur Strip-sCnc
C1544963|Bilirubin:SCnc:Pt:Urine:Qn:Test strip
C1544963|Bilirubin:Substance Concentration:Point in time:Urine:Quantitative:Test strip
C1544963|Bilirubin.total [Moles/volume] in Urine by Test strip
C1982582|Bilirubin &#124; dialysis fluid
C1982582|Bilirubin &#x7C; dialysis fluid
C0017905|Glycocholic Acid
C0017905|Glycine, N-((3alpha,5beta,7alpha,12alpha)-3,7,12-trihydroxy-24-oxocholan-24-yl)-
C0017905|Cholylglycine
C0017905|Glycocholic Acid [Chemical/Ingredient]
C0017905|N-cholylglycine
C0017905|Glycocholic acid (substance)
C0882701|Bilirubin.glucuronidated+Bilirubin.albumin bound
C2356967|Bilirubin.glucuronidated+Bilirubin.non-glucuronidated &#x7C; Bld-Ser-Plas
C1982581|Bilirubin &#x7C; cerebral spinal fluid
C1973795|Stercobilin &#x7C; stool
C1978478|Bilirubin:ACnc:Pt:Urine:Ord:Test strip.automated
C1978478|Bilirub Ur Ql Strip.auto
C1978478|Bilirubin:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip.automated
C1978478|Bilirubin.total [Presence] in Urine by Automated test strip
C1982591|Bilirubin &#x7C; urine
C1982579|Bilirubin &#x7C; Blood cord
C1982587|Bilirubin &#x7C; pleural fluid
C2924727|Bilirubin &#x7C; Skin
C0053591|21H,23H-biline-8,12-dipropanoic acid, 2,17-diethenyl-1,10,19,22,23,24-hexahydro-3,7,13,18-tetramethyl-1,19-dioxo-, mono-beta-D-glucopyranosyl ester
C0053591|bilirubin glucoside
C0056733|cyclobilirubin
C0053597|21H-biline-8,12-dipropanoic acid, 2,17-diethenyl-1,10,19,22,23,24-hexahydro-3,7,13,18-tetramethyl-1,19-dioxo-, mono-beta-D-xylopyranosyl ester
C0053597|bilirubin xyloside
C0065247|lumirubin
C0604322|Azobilirubin, mono-beta-D-glucopyranoside
C0604322|azobilirubin beta-D-monoglucoside
C0075841|taurobilirubin
C0967046|8,12-bis(2-carboxyethyl)-2,3,17,18-tetraethyl-7,13-dimethyl-10-thia-(21H,23H,24H)-bilin-1,19-dione
C0967046|thia-bilirubin
C0053588|bilirubin diglucuronide
C0053588|Bilirubin diglucuronide (substance)
C0078600|5-((3-ethyl-1,5-dihydro-4-methyl-5-oxo-2H-pyrrol-2-ylidene)methyl-2,4-dimethyl-1H-pyrrole- 3-propanoic acid
C0078600|xanthobilirubic acid
C0609875|4-iodophenylazobilirubin
C0609875|para-iodophenylazobilirubin
C0058487|ditaurobilirubin
C0053590|bilirubin ditaurine
C0053590|bilirubin ditaurate
C0053589|bilirubin dimethyl diester
C0053589|bilirubin dimethyl ester
C0053589|dimethyl bilirubin
C0607801|21H-Biline-8,12-dipropanoic acid, 2,17-diethenyl-1,10,19,22,23,24-hexahydro-3,7,13,18-tetramethyl-1,19-dioxo-, phosphate
C0607801|bilirubin phosphate
C0612575|polybilirubinate
C0969254|SEB-C10-S
C0969254|Sodium etiobilirubin-IVgamma-C10-sulfonate
C1291178|Bilirubin compound (substance)
C1291178|Bilirubin compound
C0006678|Bilirubinate, Calcium
C0006678|Calcium bilirubinate
C0006678|Salt Bilirubin, Calcium
C0006678|Calcium Salt Bilirubin
C0006678|Bilirubin, Calcium Salt
C0006678|Calcium bilirubinate (substance)
C0949235|Monosodium Salt Bilirubin
C0949235|Bilirubin, Monosodium Salt
C0949234|Disodium Salt Bilirubin
C0949234|Bilirubin, Disodium Salt
C0070952|photobilirubin
C0070952|Photobilirubin IXalpha
C0051106|albumin-bilirubin complex
C0051106|Bilirubin-albumin complex
C0051106|Bilirubin-albumin complex (substance)
C0042040|Urine bilirubin tests
C0042040|Bilirubin urine
C0042040|Urine Bilirubin Test
C0042040|Bilirubin measurement, urine
C0042040|Urine bilirubin
C0042040|Urine bilirubin level
C0042040|Bilirubin measurement, urine (procedure)
C0702270|Amniotic Fluid Bilirubin Test
C0702270|Bilirubin measurement, amniotic fluid
C0702270|Bilirubin measurement, amniotic fluid (procedure)
C1278039|serum total bilirubin
C1278039|Serum Total Bilirubin Measurement
C1278039|total serum bilirubin level
C1278039|serum total bilirubin measurement (lab test)
C1278039|Serum total bilirubin level
C1278039|Serum total bilirubin level (procedure)
C1278039|Serum bilirubin total
C1278039|Serum total bilirubin measurement (procedure)
C2711150|Measurement of total bilirubin in cord blood specimen (procedure)
C2711150|Measurement of total bilirubin in cord blood specimen
C0201913|Bilirubin; total
C0201913|Total Bilirubin Measurement
C0201913|BILIRUBIN TOTAL
C0201913|Measurement of total bilirubin
C0201913|Total bilirubin
C0201913|Total bilirubin (& level) (procedure)
C0201913|Bilirubin, total measurement
C0201913|Bilirubin, total measurement (procedure)
C0201913|Total bilirubin (& level)
C0201913|Bilirubin
C0201913|BILI
C0201913|Total bilirubin level
C0201913|Bilirubin, total measurement (procedure) [Ambiguous]
C0373554|Bilirubin; feces, qualitative
C0373554|BILIRUBIN FECES QUALITATIVE
C0373554|FECAL BILIRUBIN TEST
C0697273|Bilirubin; direct
C0697273|Bilirubin conjugated
C0697273|BILIRUBIN DIRECT
C0697273|Conjugated Bilirubin test
C1278036|Plasma total bilirubin level (procedure)
C1278036|Plasma total bilirubin level
C1278036|Plasma bilirubin total
C1278036|Plasma Total Bilirubin Test
C1278036|Plasma total bilirubin measurement (procedure)
C1278036|Plasma total bilirubin measurement
C0201917|Baby bilirubin measurement
C0201917|Bilirubin, neonatal measurement
C0201917|Bilirubin, neonatal measurement (procedure)
C0201917|Total bilirubin, neonatal measurement
C0201917|Microbilirubin measurement
C0201917|Total bilirubin, neonatal measurement (procedure)
C0428441|bilirubin
C0428441|serum bilirubin measurement (lab test)
C0428441|Serum bilirubin (& level) (procedure)
C0428441|Bilirubin - serum
C0428441|Serum bilirubin NOS (procedure)
C0428441|Serum bilirubin NOS
C0428441|Serum bilirubin level
C0428441|Serum bilirubin (& level)
C0428441|Serum bilirubin
C0428441|SB - Serum bilirubin
C0428441|Serum bilirubin measurement (procedure)
C0428441|Serum bilirubin measurement
C0863174|Blood bilirubin
C0863174|Blood bilirubin measurement
C0863174|Bilirubin
