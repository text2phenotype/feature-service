C0003467|Anxiety
C0003469|Anxiety Disorders
C0860603|Anxiety symptoms
C1963064|Anxiety Adverse Event
C4050613|Anxiety Scale (BASC-2)
C0085380|Anxieties, Dental
C0085380|Dental Anxieties
C0085380|Dental Anxiety
C0085380|Dental Fears
C0085380|Dental Phobias
C0085380|Fears, Dental
C0085380|Odontophobias
C0085380|Phobias, Dental
C0085380|DENT ANXIETY
C0085380|ANXIETY DENT
C0085380|DENT PHOBIA
C0085380|PHOBIA DENT
C0085380|FEAR DENT
C0085380|DENT FEAR
C0085380|Dental phobia (disorder)
C0085380|Dental phobia
C0085380|Dental Fear
C0085380|Odontophobia
C0085380|Fear, Dental
C0085380|Anxiety, Dental
C0085380|Phobia, Dental
C0085380|Fear of dentist
C0085380|Dental phobia (finding)
C0085380|Fear of dentist (finding)
C0003476|Anxiety, Castration
C0003476|Castration Anxiety
C0003476|Castration Complices
C0003476|Complices, Castration
C0003476|Complex, Castration
C0003476|Castration Complex
C0003476|Castration anxiety complex
C0003476|Castration anxiety complex (finding)
C0003467|Anxieties
C0003467|Anxiety
C0003467|Anxiety reaction
C0003467|rndx anxiety (diagnosis)
C0003467|rndx anxiety
C0003467|Feeling;anxious
C0003467|Anxiousness
C0003467|Anxiousness (& symptom) (finding)
C0003467|Anxiousness (& symptom)
C0003467|Anxiousness - symptom
C0003467|Anxious behavior
C0003467|-- Anxiety
C0003467|Feel anxious
C0003467|Feeling anxious
C0003467|Reaction anxiety
C0003467|Anxiety (finding)
C0003467|anxious; sensation
C0003467|Angst
C2712005|Reduced Anxiety
C0563150|Catastrophization
C0563150|Catastrophizing
C0563150|Catastrophisation
C0563150|Catastrophization (finding)
C0458631|Performance fear
C0458631|Anxiety, Performance
C0458631|Performance Anxiety
C0458631|Anxieties, Performance
C0458631|Performance Anxieties
C0458631|Performance anxiety (finding)
C2077827|anxiety which comes and goes
C2077827|anxiety episodic
C2077827|intermittent anxiety (symptom)
C2077827|anxiety which comes and goes (episodic)
C2077827|intermittent anxiety
C0549259|Anxiety aggravated
C0262376|generalized; anxiety
C0262376|anxiety; generalized
C0262377|Situational anxiety
C0235111|Anxiety complex
C0457041|Anxiety about appearing ridiculous
C0457041|Anxiety about appearing ridiculous (finding)
C0231397|Anticipatory anxiety
C0231397|Anticipatory anxiety (finding)
C0231397|Anticipatory anxiety, NOS
C0231398|Anticipatory anxiety, mild
C0231398|Anticipatory anxiety, mild (finding)
C0231400|Anticipatory anxiety, severe
C0231400|Anticipatory anxiety, severe (finding)
C0154455|Other anxiety states
C0154455|Anxiety state NEC
C0030319|Disorders, Panic
C0030319|Panic Disorder
C0030319|Panic Disorders
C0030319|Disorder, Panic
C0030319|Panic disorder [episodic paroxysmal anxiety]
C0030319|PANIC DIS
C0030319|panic anxiety syndrome
C0030319|Panic Disorder [Disease/Finding]
C0030319|Disorder;panic
C0030319|[X]Panic disorder [episodic paroxysmal anxiety] (disorder)
C0030319|[X]Panic disorder [episodic paroxysmal anxiety]
C0030319|Panic disorder (finding)
C0030319|panic disorder (diagnosis)
C0030319|-- Panic Disorder
C0030319|Panic disorder NOS
C0030319|Episodic paroxysmal anxiety disorder
C0030319|Panic disorder (disorder)
C0030319|disorder; panic
C0030319|panic; disorder
C0030319|[X]Panic disorder [episodic paroxysmal anxiety] (finding)
C2239195|Anxious mood
C2239195|mood anxious
C2239195|anxious mood (physical finding)
C2239195|Feeling anxious (finding)
C2239195|Feeling anxious
C2128827|anxious on a daily basis
C2128827|anxiety daily
C2128827|anxious every day
C2128827|daily anxiety (symptom)
C2128827|daily anxiety
C2219855|anxiety with fear of dying (symptom)
C2219855|anxiety with fear of dying
C2219855|anxiety with a fear of dying
C2219861|anxiety with feelings of unreality
C2219861|anxiety with feelings of unreality (symptom)
C0522179|Fear of death
C0522179|Thanatophobia
C0522179|Fear (of);death
C0522179|Fear (of);dying
C0522179|Death Anxiety
C0522179|Fear About Death
C0522179|Fear of dying
C0522179|Fear of dying (finding)
C0522179|Fear of death (disorder)
C0522179|Death anxiety (finding)
C0522179|Fear of death (finding)
C2219860|anxiety with dizziness or unsteady feelings (symptom)
C2219860|anxiety with dizziness or unsteady feelings
C1854339|Anxiety (with pheochromocytoma)
C0700613|Anxiety states
C0700613|Anxiety state
C0700613|Anxiety state NOS
C0700613|Anxiety state unspecified (finding)
C0700613|Anxiety state NOS (finding)
C0700613|Anxiety state unspecified
C0700613|Anxiety state, unspecified
C0700613|Anxiety state (finding)
C0700613|state; anxiety
C0700613|anxiety; state
C0474385|Anxiety about behavior or performance
C0474385|Anxiety about behaviour or performance
C0474385|Anxiety about social functioning
C0474385|Anxiety about behavior or performance (finding)
C0424145|Anxiety about body function or health
C0424145|Anxiety about health
C0424145|Anxiety about body function or health (finding)
C0558210|Anxiety about loss of control
C0558210|Anxiety about loss of control (finding)
C0558209|Anxiety about forced dependence
C0558209|Anxiety about forced dependence (finding)
C0558208|Anxiety about treatment
C0558208|Anxiety about treatment (finding)
C0870858|Mathematics Anxiety
C0424166|Social fear
C0424166|Social fear (finding)
C0424166|Social Anxiety
C0424169|Fear of public speaking
C0424169|Fear of public speaking (finding)
C0424169|Speech Anxiety
C0424169|Communication Apprehension
C0871504|Test Anxiety
C0935548|Computer Anxiety
C0577602|Anxious parent
C0577602|Anxiety;parental
C0577602|Parental anxiety
C0577602|Anxious parents
C0577602|Parental anxiety (finding)
C0700031|Anxiety attacks
C0700031|Anxiety attack
C0700031|Anxiety attack (finding)
C0700031|Attack(s);anxiety
C0231402|Moderate anxiety
C0231402|Moderate anxiety (finding)
C0231401|Mild anxiety
C0231401|Mild anxiety (finding)
C0030318|Panic
C0030318|Panics
C0030318|Panic reaction
C0030318|Panic state
C0030318|Reaction panic
C0030318|Panic (finding)
C0030318|panic; state
C0030318|state; panic
C0030318|Panic [Ambiguous]
C0233483|Free-floating anxiety
C0233483|Free-floating anxiety (finding)
C0436600|On examination - anxious
C0436600|O/E - anxious
C0436600|O/E - anxious (finding)
C0436600|On examination - anxious (context-dependent category)
C0436600|On examination - anxious (finding)
C0860603|anxiety (symptom)
C0860603|anxiety
C0860603|Anxiety symptoms
C0860603|Anxiety symptoms NOS
C0860603|anxiety; complaint
C0028768|Disorders, Obsessive-Compulsive
C0028768|Obsessive-Compulsive Disorder
C0028768|Obsessive-compulsive disorders
C0028768|Disorder, Obsessive-Compulsive
C0028768|Obsessive Compulsive Disorder
C0028768|Obsessive-compulsive disorder, unspecified
C0028768|OCD
C0028768|OBSESSIVE COMPULSIVE DIS
C0028768|obsessive compulsive disorder (diagnosis)
C0028768|OCD (obsessive compulsive disorder)
C0028768|Neuroses, Obsessive-Compulsive
C0028768|Neurosis, Obsessive Compulsive
C0028768|Obsessive-Compulsive Neurosis
C0028768|Anankastic Personalities
C0028768|Personalities, Anankastic
C0028768|Personality, Anankastic
C0028768|Obsessive-Compulsive Neuroses
C0028768|Obsessive-compulsive dis
C0028768|Obsessive-Compulsive Disorder [Disease/Finding]
C0028768|Neurosis, Obsessive-Compulsive
C0028768|Anankastic Personality
C0028768|Disorder;obsessive-compulsive
C0028768|Anancastic neurosis
C0028768|[X]Obsessive-compulsive disorder, unspecified
C0028768|[X]Obsessive-compulsive disorder, unspecified (disorder)
C0028768|Obsessive-compulsive disorder (disorder)
C0028768|OCD - Obsessive-compulsive disorder
C0028768|Anankastic neurosis
C0028768|Obsessive compulsive disorder (disorder)
C0028768|Obsessive compulsive neurosis
C0028768|Obsessive-compulsive disorder NOS
C0028768|Obsessive-compulsive disorder NOS (disorder)
C0028768|-- Obsessive Compulsive Disorder
C0028768|Reaction obsessive-compulsive
C0028768|Obsessive-compulsive reaction
C0028768|disorder; obsessive-compulsive
C0028768|neurosis; anankastic
C0028768|neurosis; obsessive-compulsive
C0028768|obsessive-compulsive neurosis or reaction
C0028768|obsessive-compulsive; disorder
C0028768|obsessive-compulsive; neurosis
C0028768|obsessive-compulsive; reaction
C0028768|reaction; obsessive-compulsive
C0028768|anankastic; neurosis
C0028768|Obsessive compulsive disorder, NOS
C0349231|Phobia
C0349231|Disorder, Phobic
C0349231|Disorders, Phobic
C0349231|Phobic Disorder
C0349231|Phobic Disorders
C0349231|Phobic anxiety disorder, unspecified
C0349231|Phobic anxiety disorders
C0349231|Phobic state
C0349231|PHOBIC DIS
C0349231|Phobic anxiety disorder
C0349231|phobia (diagnosis)
C0349231|Phobia NOS
C0349231|Phobic state NOS
C0349231|Neuroses, Phobic
C0349231|Phobic Disorders [Disease/Finding]
C0349231|Phobias
C0349231|Phobic Neuroses
C0349231|Phobias NOS
C0349231|[X]Phobic anxiety disorder, unspecified (disorder)
C0349231|Phobia (finding)
C0349231|[X]Phobic anxiety disorders
C0349231|Phobic disorder NOS
C0349231|Phobic disorder NOS (finding)
C0349231|Phobic anxiety
C0349231|[X]Phobic anxiety disorder, unspecified
C0349231|Phobia unspecified
C0349231|Phobic anxiety disorder (disorder)
C0349231|[X]Phobic anxiety disorders (disorder)
C0349231|Phobic neurosis
C0349231|Abnormal fear
C0349231|Phobia unspecified (finding)
C0349231|Phobia, unspecified
C0349231|Phobic disorder (disorder)
C0349231|neurosis; phobic
C0349231|phobia; state
C0349231|phobic; anxiety disorder
C0349231|phobic; neurosis
C0349231|phobic; state
C0349231|state; phobia
C0349231|state; phobic
C0349231|anxiety disorder; phobic
C0349231|Phobia, NOS
C0038436|Post-traumatic stress disorder
C0038436|Neuroses, Post Traumatic
C0038436|Post Traumatic Stress Disorders
C0038436|Post-Traumatic Neuroses
C0038436|Posttraumatic Neuroses
C0038436|Posttraumatic Stress Disorder
C0038436|PTSD
C0038436|Stress Disorder, Post-Traumatic
C0038436|Stress Disorder, Posttraumatic
C0038436|Stress Disorders, Post Traumatic
C0038436|Stress Disorders, Post-Traumatic
C0038436|Post-Traumatic Stress Disorder (PTSD)
C0038436|POSTTRAUMATIC STRESS DISORDERS
C0038436|POST TRAUMATIC STRESS DIS
C0038436|POSTTRAUMATIC STRESS DIS
C0038436|STRESS DIS POSTTRAUMATIC
C0038436|STRESS DIS POST TRAUMATIC
C0038436|combat fatigue
C0038436|traumatic neurosis
C0038436|post-traumatic stress disorder (diagnosis)
C0038436|Post-traumatic stress disorder, unspecified
C0038436|Stress Disorder, Post Traumatic
C0038436|Post-Traumatic Stress Disorders
C0038436|Neuroses, Posttraumatic
C0038436|Stress Disorders, Post-Traumatic [Disease/Finding]
C0038436|Stress Disorders, Posttraumatic
C0038436|Neuroses, Post-Traumatic
C0038436|Disorder;post traumatic stress
C0038436|Post-traumatic stress disorder (disorder)
C0038436|-- Post Traumatic Stress Disorder
C0038436|PTSD - Post-traumatic stress disorder
C0038436|Post-traumatic stress syndrome
C0038436|Posttraumatic stress disorder (disorder)
C0038436|disorder, post-traumatic stress
C0038436|disorder; post-traumatic stress
C0038436|disorder; stress, post-traumatic
C0038436|neurosis; traumatic
C0038436|post-traumatic stress; disorder
C0038436|stress; disorder, post-traumatic
C0038436|traumatic; neurosis
C0038436|Posttraumatic stress disorder, NOS
C0038436|Posttraumatic stress disorder NOS
C0038436|post traumatic stress disorder
C0027821|Asthenias, Neurocirculatory
C0027821|Cardiac Neuroses
C0027821|Neurocirculatory Asthenia
C0027821|Neurocirculatory Asthenias
C0027821|Neuroses, Cardiac
C0027821|Asthenia, Neurocirculatory
C0027821|Neurosis, Cardiac
C0027821|Syndrome, Effort
C0027821|cardiac neurosis (diagnosis)
C0027821|cardiac neurosis
C0027821|Psychogen cardiovasc dis
C0027821|Neurocirculatory Asthenia [Disease/Finding]
C0027821|Effort Syndrome
C0027821|Neurosis;cardiac
C0027821|[X]Neurocirculatory asthenia
C0027821|[X]Cardiac neurosis
C0027821|[X]Da Costa's syndrome
C0027821|Cardiovascular disorder, psychogenic
C0027821|Cardiac neurosis (disorder)
C0027821|Da Costa's syndrome
C0027821|Cardiovascular neurosis
C0027821|Cerebrocardiac neurosis
C0027821|Neurocirculatory asthenia (finding)
C0027821|Cerebrocardiac neurosis (disorder)
C0027821|Cerebrocardiac syndrome
C0027821|Irritable heart syndrome
C0027821|Cardioneurosis
C0027821|Krishaber's disease
C0027821|Syndrome effort
C0027821|Neurosis cardiovascular
C0027821|Cardiovascular malfunction arising from mental factors
C0027821|Neurocirculatory asthenia (disorder)
C0235245|Psychogenic syncope
C0235245|[X] Psychogenic syncope
C0235245|[X]Psychogenic syncope
C0235245|psychogenic syncope (diagnosis)
C0235245|Psychogenic syncope (disorder)
C0856254|Neurotic personality
C0860602|Anxious personality
C0236121|Neurosis GI
C0236121|Gastrointestinal neurosis
C0270549|Generalized anxiety disorder
C0270549|Generalised anxiety disorder
C0270549|generalized anxiety disorder (diagnosis)
C0270549|GAD
C0270549|Generalized anxiety dis
C0270549|Generalised anxiety disorder (disorder)
C0270549|GAD - Generalised anxiety disorder
C0270549|GAD - Generalized anxiety disorder
C0270549|Generalized anxiety disorder (disorder)
C0270549|generalized; anxiety disorder
C0270549|anxiety disorder; generalized
C0270549|Generalised anxiety disorder [Ambiguous]
C0001818|Agoraphobia
C0001818|Agoraphobias
C0001818|Fear of open spaces
C0001818|Agoraphobia, unspecified
C0001818|Agoraphobia [Disease/Finding]
C0001818|agoraphobia (diagnosis)
C0001818|[X]Agoraphobia
C0001818|Agoraphobia (disorder)
C0001818|Fear of open places
C0001818|Phobia of going out
C0001818|Fear of open spaces (finding)
C0001818|Agoraphobia, NOS
C0038441|TRAUMATIC STRESS DIS
C0038441|Stress disorders
C0038441|Stress Disorders, Traumatic [Disease/Finding]
C0038441|Stress Disorders, Traumatic
C0038441|stress disorder (diagnosis)
C0038441|stress disorder
C0038441|Stress Disorder, Traumatic
C0038441|Traumatic Stress Disorder
C0038441|Traumatic Stress Disorders
C0038441|disorder; stress
C0038441|stress; disorder
C0003469|Anxiety Disorder
C0003469|Anxiety Disorders
C0003469|Disorder, Anxiety
C0003469|Disorders, Anxiety
C0003469|Anxiety disorder, unspecified
C0003469|ANXIETY DIS
C0003469|anxiety disorder (diagnosis)
C0003469|Anxiety NOS
C0003469|Anxiety Disorders [Disease/Finding]
C0003469|Anxiety disorder (disorder)
C0003469|[X]Anxiety disorder, unspecified
C0003469|[X]Anxiety disorder, unspecified (disorder)
C0003469|Anxiety
C0003469|Anxiety disorder, NOS
C0003469|Anxiety disorder [Ambiguous]
C0003469|Disorder;anxiety
C0376280|Anxiety State, Neurotic
C0376280|Neurotic Anxiety State
C0376280|Neurotic Anxiety States
C0376280|State, Neurotic Anxiety
C0376280|States, Neurotic Anxiety
C0376280|Anxiety States, Neurotic
C0086769|Attacks, Panic
C0086769|Panic attack
C0086769|Attack, Panic
C0086769|Panic attacks
C0086769|Attack(s);panic
C0086769|Panic attack (finding)
C0086769|attack; panic
C0086769|panic; attack
C0236816|Acute Stress Disorder
C0236816|Acute stress reaction
C0236816|STRESS DIS ACUTE
C0236816|STRESS DIS TRAUMATIC ACUTE
C0236816|ACUTE STRESS DIS
C0236816|acute stress disorder (diagnosis)
C0236816|acute reaction to stress
C0236816|acute reaction to stress (diagnosis)
C0236816|Gross stress reaction, NOS
C0236816|Acute stress react NOS
C0236816|Acute crisis reaction
C0236816|Psychic shock
C0236816|Stress Disorders, Acute
C0236816|Stress Disorders, Traumatic, Acute
C0236816|Acute Stress Disorders
C0236816|Stress Disorders, Traumatic, Acute [Disease/Finding]
C0236816|Reaction after;acute stress
C0236816|Acute stress reaction NOS (disorder)
C0236816|Post-traumatic stress - acute
C0236816|[X]Acute reaction to stress
C0236816|Acute stress reaction NOS
C0236816|Gross stress reaction (disorder)
C0236816|Gross stress reaction
C0236816|[X]Psychic shock
C0236816|Psychic shock (disorder)
C0236816|[X]Acute crisis reaction
C0236816|(Examination fear) or (flying phobia) or (stage fright) or (acute stress reaction NOS) (disorder)
C0236816|(Examination fear) or (flying phobia) or (stage fright) or (acute stress reaction NOS)
C0236816|[X]Acute stress reaction
C0236816|Stress Disorder, Acute
C0236816|Acute reaction to stress, unspecified
C0236816|Unspecified acute reaction to stress
C0236816|Acute stress disorder (disorder)
C0236816|crisis; acute reaction
C0236816|disorder; acute stress
C0236816|acute reaction; crisis
C0236816|acute; stress disorder
C0236816|acute; stress reaction
C0236816|psychic; shock
C0236816|shock; psychic
C0236816|stress reaction; acute
C2985218|Substance-Induced Anxiety Disorder
C1279420|Anxiety neurosis
C1279420|Anxiety Neuroses
C1279420|Anxiety neurosis (finding)
C1279420|neurosis; anxiety
C1279420|anxiety; neurosis
C1279420|Neuroses, Anxiety
C0236794|panic disorder without agoraphobia (diagnosis)
C0236794|panic disorder without agoraphobia
C0236794|Panic dis w/o agorphobia
C0236794|Panic disorder [episodic paroxysmal anxiety] without agoraphobia
C0236794|[X]Agoraphobia without history of panic disorder
C0236794|Panic disorder without agoraphobia (disorder)
C0236794|Panic disorder without agoraphobia, NOS
C0236800|panic disorder with agoraphobia
C0236800|panic disorder with agoraphobia (diagnosis)
C0236800|Agoraphobia w panic dis
C0236800|Agoraphobia with panic disorder
C0236800|[X]Panic disorder with agoraphobia
C0236800|panic disorder with agoraphobia and panic attacks
C0236800|panic disorder with agoraphobia and panic attacks (diagnosis)
C0236800|Panic disorder with agoraphobia (disorder)
C0236800|disorder; panic, with agoraphobia
C0236800|panic; disorder, with agoraphobia
C0236800|Panic disorder with agoraphobia, NOS
C1387823|mixed anxiety disorder
C1387823|anxiety disorder mixed
C1387823|mixed anxiety disorder (diagnosis)
C1387823|mixed; anxiety disorder
C1387823|anxiety disorder; mixed
C0236730|Sedative, hypnotic AND/OR anxiolytic-induced anxiety disorder (disorder)
C0236730|Sedative, hypnotic AND/OR anxiolytic-induced anxiety disorder
C0236730|Sedative, hypnotic or anxiolytic-induced anxiety disorder
C0236715|cocaine induced anxiety disorder (diagnosis)
C0236715|cocaine induced anxiety disorder
C0236715|Cocaine-induced anxiety disorder
C0236715|Cocaine-induced anxiety disorder (disorder)
C0236715|cocaine; anxiety disorder
C0236715|anxiety disorder; due to cocaine
C0236801|Specific (isolated) phobias
C0236801|PHOBIA, SPECIFIC
C0236801|Specific phobias
C0236801|Phobia, Simple
C0236801|[X]Specific (isolated) phobias
C0236801|[X]Simple phobia
C0236801|Specific Phobia
C0236801|simple phobia
C0236801|specific phobia (diagnosis)
C0236801|simple (specific) phobia
C0236801|Isolated phobia
C0236801|Simple phobia (disorder)
C0236801|phobia; simple
C0236801|phobia; specific
C0236801|simple; phobia
C0236801|specific; phobia
C0031572|Social phobia
C0031572|Phobias, Social
C0031572|Social Phobias
C0031572|social phobia (diagnosis)
C0031572|Social phobia, unspecified
C0031572|Social neurosis
C0031572|Social phobia (disorder)
C0031572|Social phobic disorders
C0031572|Social Anxiety Disorder
C0031572|-- Social Phobia
C0031572|neurosis; social
C0031572|phobia; social
C0031572|social; neurosis
C0031572|social; phobia
C0031572|anxiety disorder; social
C0031572|Social phobia, NOS
C0031572|Phobia, Social
C0003477|Separation Anxiety Disorder
C0003477|Separation anxiety
C0003477|anxiety separation
C0003477|separation anxiety (diagnosis)
C0003477|Separation anxiety (disorder)
C0003477|disorder; separation anxiety
C0003477|separation anxiety; disorder
C0003471|Anxiety disorder of childhood OR adolescence
C0003471|anxiety disorder of childhood or adolescence (diagnosis)
C0003471|Anxiety disorder of childhood OR adolescence (disorder)
C0003471|Anxiety disorder of childhood or adolescence, NOS
C0270590|anxiety hyperventilation (diagnosis)
C0270590|Anxiety hyperventilation
C0270590|Anxiety hyperventilation (disorder)
C0236748|Organic anxiety disorder
C0236748|Anxiety Disorder Due to Specified Medical Condition
C0236748|Anxiety disorder due to a general medical condition
C0236748|anxiety disorder due to general medical condition
C0236748|anxiety disorder due to general medical condition (diagnosis)
C0236748|Anxiety disorder due to medical disorder
C0236748|Organic anxiety disorder (disorder)
C0236748|anxiety disorder organic
C0236748|Organic anxiety disorder (diagnosis)
C0236748|Organic anxiety syndrome
C0236748|Anxiety disorder due to a general medical condition (disorder)
C0236748|disorder; anxiety, organic
C0236748|disorder; organic, anxiety
C0236748|medical condition; causing anxiety disorder
C0236748|organic; anxiety disorder
C0236748|organic; disorder, anxiety
C0236748|anxiety disorder; due to general medical condition
C0236748|anxiety disorder; organic
C1842981|NEUROTICISM
C3840205|Anxiety in childbirth
C3840205|Anxiety disorder in mother complicating childbirth (disorder)
C3840205|Anxiety disorder in mother complicating childbirth
C0027932|Neurosis
C0027932|Disorders, Neurotic
C0027932|Neurotic Disorder
C0027932|Neurotic Disorders
C0027932|Disorder, Neurotic
C0027932|Psychoneurosis
C0027932|Neurotic disorder, unspecified
C0027932|NEUROTIC DIS
C0027932|Neurosis NOS
C0027932|Neuroses
C0027932|Psychoneuroses
C0027932|Neurotic Disorders [Disease/Finding]
C0027932|[X]Neurotic disorder, unspecified (disorder)
C0027932|[X] Neurosis NOS
C0027932|[X]Neurosis NOS
C0027932|[X]Neurotic disorder, unspecified
C0027932|Neurotic disorder NOS (disorder)
C0027932|Neurotic disorder NOS
C0027932|Neurotic disorder (disorder)
C0027932|psychiatric disorders neurosis
C0027932|neurosis (diagnosis)
C0027932|Unspecified neurotic disorder
C0027932|Neurosis (disorder)
C0027932|Nonpsychotic mental disorder
C0027932|disease (or disorder); neurotic
C0027932|disorder; mental, neurotic
C0027932|disorder; neurotic
C0027932|mental; disorder, neurotic
C0027932|neurosis; state
C0027932|neurotic; disorder
C0027932|neurotic; state
C0027932|state; neurosis
C0027932|state; neurotic
C0027932|Neurosis, NOS
C0027932|Nonpsychotic mental disorder, NOS
C0027932|Psychoneurosis NOS
C0027932|Disorder;neurotic
C0027932|Neurotic
C1527281|Anxiety, Separation
C1527281|Separation Anxiety
C1527281|Separation anxiety disorder of childhood
C1527281|separation anxiety disorder of childhood (diagnosis)
C1527281|Anxiety Disorder, Separation
C1527281|SEPARATION ANXIETY DIS
C1527281|Anxiety, Separation [Disease/Finding]
C1527281|Separation Anxiety Disorder
C1527281|[X]Separation anxiety disorder of childhood (disorder)
C1527281|[X]Separation anxiety disorder of childhood
C1527281|Separation anxiety disorder of childhood (disorder)
C4042925|Trauma and Stressor Related Disorders
C4042925|Trauma and Stressor Related Disorders [Disease/Finding]
C4042925|trauma and stressor-related disorder
C4042925|other psychiatric disorders trauma and stressor-related
C4042925|trauma and stressor-related disorder (diagnosis)
C3887605|nightmare disorder
C3887605|nightmare disorder (diagnosis)
C3887605|Dream anxiety disorder
C3887605|[X]Dream anxiety disorder
C3887605|[X] Nightmares or dream anxiety disorder
C3887605|[X] Nightmares or dream anxiety disorder (disorder)
C3887605|Paroniria
C3887605|Nightmare
C3887605|Dream anxiety disorder (disorder)
C3887605|Nightmare, NOS
C3887605|Nightmares
C3887605|Nightmares NOS
C0338908|Mixed anxiety and depressive disorder
C0338908|depression with anxiety
C0338908|depression with anxiety (diagnosis)
C0338908|Anxiety/depression
C0338908|Anxiety with depression
C0338908|Mixed anxiety and depressive disorder (disorder)
C0338908|[X]Mixed anxiety and depressive disorder
C0338908|Anxiety depression
C0338908|Anxious depression
C0338908|Mixed anxiety & depressive
C0338908|depression; anxiety
C0338908|disorder; mixed, anxiety and depressive
C0338908|mixed; disorder, anxiety and depressive
C0338908|anxiety; depression
C0236708|amphetamine-induced anxiety disorder (diagnosis)
C0236708|amphetamine-induced anxiety disorder
C0236708|Amphetamine induced anxiety disorder
C0236708|Amphetamine-induced anxiety disorder (disorder)
C0520683|Occupation-related stress disorder
C0520683|occupation-related stress disorder (diagnosis)
C0520683|Occupation-related stress disorder (disorder)
C0520683|Work-related stress disorder
C0520683|Occupation-related stress disorder, NOS
C0520683|Work-related stress disorder, NOS
C0476644|Physical and emotional exhaustion state
C0476644|Burnout
C0476644|Burnt out
C0476644|Burnt out (qualifier value)
C0476644|Physical AND emotional exhaustion state (disorder)
C0476644|burn-out
C0302832|Obsessional neurosis
C0302832|Neurosis;obsessive
C0302832|obsessional neurosis (diagnosis)
C0302832|Obsessional neurosis (disorder)
C0302832|Obsessive reaction
C0302832|neurosis; obsessional
C0302832|neurosis; obsession
C0302832|obsession; neurosis
C0302832|obsessional; neurosis
C0302832|Obsessive Neurosis
C1879354|Separation anxiety
C1879354|Separation anxiety (finding)
C1879354|separation; anxiety
C1879354|anxiety; separation
C1879354|Anxiety;separation
C1387810|fear; reaction
C1387810|reaction; fear
C1408583|apprehensiveness; abnormal
C0850602|Chronic stress disorder
C0850602|Chronic stress disorder (disorder)
C0850602|chronic stress disorder (diagnosis)
C0850602|Disorder;chronic stress
C2063171|anxiety disorder of unknown (Axis III) etiology (diagnosis)
C2063171|anxiety disorder of unknown (Axis III) etiology
C0085631|Agitation
C0085631|Agitated (& symptom) (finding)
C0085631|Agitated behaviour
C0085631|Agitated (& symptom)
C0085631|Excessive overactivity
C0085631|Agitated behavior (finding)
C0085631|Agitated
C0085631|Feeling agitated
C0085631|Agitated - symptom
C0085631|Feeling agitated (finding)
C0085631|Increased purposeless goalless activity
C0085631|Agitated behavior
C0085631|Excitement abnormal
C0085631|Unable to keep still
C0085631|Excessive overactivity, NOS
C0085631|Increased purposeless goalless activity, NOS
C0235844|Agitation neonatal
C0235844|Neonatal agitation
C0235844|Neonatal agitation (disorder)
C0392156|Akathisia
C0392156|Akithisia
C0392156|feeling an alien urge to be in motion (akathisia)
C0392156|feeling an alien urge to be in motion (akathisia) (symptom)
C0392156|akathisia (diagnosis)
C0392156|Akathisia (disorder)
C0392156|Akathisia (finding)
C0392156|Acathisia
C0392156|Acathesia
C0027769|Nervousness
C0027769|Nervous tension
C0027769|[D]Nervousness (context-dependent category)
C0027769|Nervous
C0027769|Nervy
C0027769|Feeling of Nervousness
C0027769|Tension - nervous
C0027769|"Nerves" - nervousness
C0027769|[D]Nervous tension
C0027769|Nervously anxious
C0027769|"Nerves"
C0027769|[D]Nervousness (situation)
C0027769|["Nerves"] or [nervousness] or [nervous tension] (finding)
C0027769|["Nerves"] or [nervousness] or [nervous tension]
C0027769|Nervousness (finding)
C0027769|[D]Nervousness
C0027769|[D]Nerves
C0027769|Tension nervous
C0027769|nervous; tension
C0027769|tension; nervous
C0038435|Stress
C0038435|State of stress
C0038435|Stress (finding)
C0038435|Stress (qualifier value)
C0038435|Stress - value
C0038435|state; stress
C0038435|stress; state
C0038435|Pressure, NOS
C0038435|Stress, NOS
C0233494|Tension
C0233494|Tense Feeling
C0233494|Tense
C0233494|Mental tension
C0233494|Tension (finding)
C0233494|mental; tension
C0233494|state; tension state
C0233494|tension; mental
C0919572|Agitation postoperative
C1112506|Pseudoangina
C1112506|Angina pectoris falsa
C1868709|Activation syndrome
C2128829|anxiety relieved by medication (symptom)
C2128829|anxiety relieved by medication
C2128830|anxiety with fear of going crazy (symptom)
C2128830|anxiety with fear of going crazy
C2128830|anxiety with a fear of going crazy
C2128831|anxiety with fear of losing self-control (symptom)
C2128831|anxiety with fear of losing self-control
C2128831|anxiety with a fear of losing self-control
C2219852|anxiety with persistent worry (symptom)
C2219852|anxiety with a persistent worry
C2219852|anxiety with persistent worry
C2219854|anxiety with anticipation of misfortune
C2219854|anxiety with anticipation of misfortune (symptom)
C2219854|anxiety with an anticipation of misfortune to self or others
C2219856|anxiety with difficulty breathing (symptom)
C2219856|anxiety with difficulty breathing
C2219857|anxiety with chest pain or discomfort (symptom)
C2219857|anxiety with chest pain or discomfort
C2219858|anxiety with rapid heartbeat (symptom)
C2219858|anxiety with rapid heartbeat
C2219859|anxiety with choking or smothering sensations
C2219859|anxiety with choking or smothering sensations (symptom)
C2219862|anxiety with tingling in hands and feet (symptom)
C2219862|anxiety with tingling in hands and feet
C2219863|anxiety with muscle tension, jitters (symptom)
C2219863|anxiety with muscle tension, jitters
C2219864|anxiety with stomach discomfort
C2219864|anxiety with stomach discomfort (symptom)
C2219865|anxiety with frequent urination or diarrhea
C2219865|anxiety with frequent urination or diarrhea (symptom)
C2219866|anxiety with hot and cold flashes
C2219866|anxiety with hot and cold flashes (symptom)
C2219867|anxiety with excessive sweating
C2219867|anxiety with excessive sweating (symptom)
C2219869|anxiety unrelated to exertion or dangerous situation
C2219869|anxiety unrelated to exertion or dangerous situation (symptom)
C2219869|anxiety unrelated to exertion or danger situation
C2219871|continuous anxiety for a month or more
C2219871|anxiety continuously for a month or more
C2219871|anxiety continuously for a month or more (symptom)
C2219905|anxiety with unrealistic fear of disease (symptom)
C2219905|anxiety with unrealistic fear of disease
C2219939|anxiety from anticipation of separation (symptom)
C2219939|anxiety from anticipation of separation
C2219951|anxiety which interferes with social activities (symptom)
C2219951|anxiety which interferes with social activities
C2219951|anxiety interferes with social activities
C2219952|anxiety which interferes with work (symptom)
C2219952|anxiety which interferes with work
C2219952|anxiety interferes with work
C2219955|anxiety relieved by checking (symptom)
C2219955|anxiety relieved by checking
C2219956|anxiety relieved by washing
C2219956|anxiety relieved by washing (symptom)
C2219957|anxiety relieved by a ritual (symptom)
C2219957|anxiety relieved by a ritual
C3162298|anxiety about medical condition (symptom)
C3162298|anxiety about medical condition
C3162299|anxiety about medical regimen
C3162299|anxiety about medical regimen (symptom)
C3854439|Procedural anxiety
C3854440|Immunisation anxiety related reaction
C3854440|Immunization anxiety related reaction
C3864091|anxiety about planned surgery
C3864091|anxiety about planned surgery (symptom)
C1561362|CTCAE Grade 2 Anxiety
C1561362|Grade 2 Anxiety
C1561364|CTCAE Grade 4 Anxiety
C1561364|Grade 4 Anxiety
C1561361|CTCAE Grade 1 Anxiety
C1561361|Grade 1 Anxiety
C1561365|CTCAE Grade 5 Anxiety
C1561365|Grade 5 Anxiety
C1561363|CTCAE Grade 3 Anxiety
C1561363|Grade 3 Anxiety
