C0003289|Antidepressive Agents
C0003289|Antidepressive Drugs
C0003289|Antidepressive Medications
C0360105|Selective Serotonin Reuptake Inhibitors
C0360105|SSRI
C0719199|Celexa
C0162373|Prozac
C0376414|Paxil
C0284660|Zoloft
C0678176|Neurontin
C0657912|pregabalin
C1570232|Lyrica
C0074393|sertraline
C0074393|1-Naphthalenamine,1,2,3,4-tetrahydro-4-(3,4-dichlorophenyl)-N-methyl-, (1S-cis)-
C0074393|Sertraline [Chemical/Ingredient]
C0074393|Sertraline (product)
C0074393|Sertraline (substance)
C0078569|venlafaxine
C0078569|antidepressants venlafaxine
C0078569|venlafaxine (medication)
C0078569|1-(2-(dimethylamino)-1-(4-methoxyphenyl)ethyl)cyclohexanol
C0078569|Venlafaxine [Chemical/Ingredient]
C0078569|Venlafaxine (product)
C0078569|Venlafaxine (substance)
C0078569|VNF
C0003290|Agents, Tricyclic Antidepressive
C0003290|Antidepressive Agents, Tricyclic
C0003290|tricyclic antidepressant
C0003290|Tricyclic Antidepressants
C0003290|Drugs, Tricyclic Antidepressant
C0003290|Tricyclic Antidepressant Drugs
C0003290|tricyclic antidepressants (medication)
C0003290|[CN601] TRICYCLIC ANTIDEPRESSANTS
C0003290|Tricyclic Antidepressive Agents
C0003290|Tricyclic antidepressant drug
C0003290|Tricyclic antidepressant drug (substance)
C0003290|Antidepressants, Tricyclic
C0003290|Antidepressant Drugs, Tricyclic
C0003290|Tricyclic antidepressant (product)
C0003290|Tricyclic antidepressant (substance)
C0003290|Tricyclic antidepressant, NOS
C0016365|Fluoxetine
C0016365|Benzenepropanamine, N-methyl-gamma-(4-(trifluoromethyl)phenoxy)-, (+-)-
C0016365|N-methyl-gamma-(4-(trifluoromethyl) -phenoxy)-benzenepropanamine
C0016365|Fluoxetin
C0016365|N-Methyl-gamma-(4-(trifluoromethyl)phenoxy)benzenepropanamine
C0016365|Fluoxetine [Chemical/Ingredient]
C0016365|Fluoxetine (product)
C0016365|Fluoxetine (substance)
C0016365|FLUOX
C0031392|2 Phenethylhydrazine
C0031392|Phenelzine
C0031392|beta Phenylethylhydrazine
C0031392|Hydrazine, (2-phenylethyl)-
C0031392|Fenelzin
C0031392|beta-Phenylethylhydrazine
C0031392|Phenethylhydrazine
C0031392|Phenelzine [Chemical/Ingredient]
C0031392|2-Phenethylhydrazine
C0031392|antidepressants phenelzine
C0031392|phenelzine (medication)
C0031392|MAOI - Phenelzine
C0031392|Phenelzine (product)
C0031392|Phenelzine (substance)
C0085208|Bupropion
C0085208|1-Propanone, 1-(3-chlorophenyl)-2-((1,1-dimethylethyl)amino)-
C0085208|Amfebutamone
C0085208|bupropion (medication)
C0085208|(+-)-1-(3-Chlorophenyl)-2-((1,1-dimethylethyl)amino)-1-propanone
C0085208|Bupropion [Chemical/Ingredient]
C0085208|Amfebutamon
C0085208|Bupropion (substance)
C0085208|Bupropion (product)
C0085208|BUP
C0085208|Bupropion [dup] (substance)
C0070122|Paroxetine
C0070122|Piperidine, 3-((1,3-benzodioxol-5-yloxy)methyl)-4-(4-fluorophenyl)-, (3S-trans)-
C0070122|(-)-trans-4-(p-fluorophenyl)-3-((3,4-(methylenedioxy)phenoxy)methyl)piperidine
C0070122|(-)-(3S,4R)-4-(p-Fluorophenyl)-3-((3,4-(methylenedioxy)phenoxy)methyl)piperidine
C0070122|Paroxetine [Chemical/Ingredient]
C0070122|Paroxetine (product)
C0070122|Paroxetine (substance)
C0008845|Citalopram
C0008845|5-Isobenzofurancarbonitrile, 1-(3-(dimethylamino)propyl)-1-(4-fluorophenyl)-1,3-dihydro-
C0008845|Cytalopram
C0008845|Citalopram [Chemical/Ingredient]
C0008845|Nitalapram
C0008845|1,3-Dihydro-1-(3-(dimethylamino)propyl)-1-(4-fluorophenyl)-5-isobenzofurancarbonitrile
C0008845|Citalopram (product)
C0008845|Citalopram (substance)
C0085228|Fluvoxamine
C0085228|1-Pentanone, 5-methoxy-1-(4-(trifluoromethyl)phenyl)-, O-(2-aminoethyl)oxime, (E)-
C0085228|Fluvoxamine [Chemical/Ingredient]
C0085228|Fluvoxamine (product)
C0085228|Fluvoxamine (substance)
C0085228|Fluoxamine
C0004962|Benactyzine
C0004962|Benzeneacetic acid, alpha-hydroxy-alpha-phenyl-, 2-(diethylamino)ethyl ester
C0004962|Benactyzine [Chemical/Ingredient]
C0004962|Benactyzine (substance)
C0009035|Clorgyline
C0009035|2-Propyn-1-amine, N-(3-(2,4-dichlorophenoxy)propyl)-N-methyl-
C0009035|Clorgiline
C0009035|Clorgyline [Chemical/Ingredient]
C0009035|Clorgilin
C0009035|Chlorgyline
C0011064|Deanol
C0011064|Ethanol, 2-(dimethylamino)-
C0011064|N,N Dimethyl 2 hydroxyethylamine
C0011064|Dimethylethanolamine
C0011064|Dimethyl ethanolamine
C0011064|parasympathomimetics deanol
C0011064|deanol (medication)
C0011064|N,N-Dimethyl-N-(2-hydroxyethyl)amine
C0011064|2-Dimethylaminoethanol
C0011064|Dimethylaminoethanol
C0011064|Demanyl
C0011064|Demanol
C0011064|N,N-Dimethyl-2-hydroxyethylamine
C0011064|N,N-Dimethylethanolamine
C0011064|Deanol [Chemical/Ingredient]
C0011064|Dimethyl ethanolamine (substance)
C0011064|Deanol (substance)
C0011064|2 Dimethylaminoethanol
C0022059|Iproniazid
C0022059|4-Pyridinecarboxylic acid, 2-(1-methylethyl)hydrazide
C0022059|Iprazid
C0022059|Iproniazid [Chemical/Ingredient]
C0022059|1-Isonicotinoyl-2-isopropylhydrazine
C0022059|Iproniazid (product)
C0022059|Iproniazid (substance)
C0022154|Isocarboxazid
C0022154|3-Isoxazolecarboxylic acid, 5-methyl-, 2-(phenylmethyl)hydrazide
C0022154|Ro 5-0831
C0022154|isocarboxazid (medication)
C0022154|Isocarboxazid [Chemical/Ingredient]
C0022154|MAOI - Isocarboxazid
C0022154|Isocarboxazid (product)
C0022154|Isocarboxazid (substance)
C0027999|Nialamide
C0027999|4-Pyridinecarboxylic acid, 2-(3-oxo-3-((phenylmethyl)amino)propyl)hydrazide
C0027999|1-(2-(Benzylcarbamoyl)ethyl)-2-isonicotinoylhydrazine
C0027999|Nialamide [Chemical/Ingredient]
C0027999|Nialamide (substance)
C0032036|Pizotyline
C0032036|Piperidine, 4-(9,10-dihydro-4H-benzo(4,5)cyclohepta(1,2-b)thien-4-ylidene)-1-methyl-
C0032036|Pizotyline product
C0032036|Pizotifen
C0032036|Pizotyline [Chemical/Ingredient]
C0032036|4-(9,10-Dihydro-4H-Benzo(4,5)Cyclohepta(1,2-B)Thien-4-ylidene)-1-Methylpiperidine
C0032036|Pizotifen product (substance)
C0032036|Pizotifen product
C0032036|Pizotifen (product)
C0032036|Pizotifen (substance)
C0040778|Tranylcypromine
C0040778|trans 2 Phenylcyclopropylamine
C0040778|Cyclopropanamine, 2-phenyl-, trans-(+-)-
C0040778|Tranylcypromine [Chemical/Ingredient]
C0040778|trans-2-Phenylcyclopropylamine
C0040778|antidepressants tranylcypromine
C0040778|tranylcypromine (medication)
C0040778|MAOI - Tranylcypromine
C0040778|Tranylcypromine (product)
C0040778|Tranylcypromine (substance)
C0206486|Lithium Compounds
C0206486|Compounds, Lithium
C0206486|LITHIUM CPDS
C0206486|Lithium Compounds [Chemical/Ingredient]
C0206486|Lithium compound (substance)
C0206486|Lithium compound
C0206486|Lithium compound, NOS
C0073561|Rolipram
C0073561|Pyrrolidone, 4-(3-cyclopentyloxy-4-methoxyphenyl)-2-
C0073561|Rolipram [Chemical/Ingredient]
C0073561|(+/-)-Rolipram
C0073561|(R,S)-Rolipram
C0066673|Moclobemide
C0066673|moclobemide (medication)
C0066673|Benzamide, 4-Chloro-N-(2-(4-morpholinyl)ethyl)-
C0066673|Moclobamide
C0066673|Moclobemide [Chemical/Ingredient]
C0066673|P-Chloro-N-(2-Morpholinoethyl)Benzamide
C0066673|Moclobemide (product)
C0066673|Moclobemide (substance)
C0242905|Agents, Second-Generation Antidepressive
C0242905|Antidepressive Agents, Second Generation
C0242905|Antidepressive Agents, Second-Generation
C0242905|Antidepressive Drugs, Second Generation
C0242905|Drugs, Second-Generation Antidepressive
C0242905|Second Generation Antidepressive Agents
C0242905|Second-Generation Antidepressive Drugs
C0242905|Second-Generation Antidepressive Agents
C0242905|Antidepressants, Atypical
C0242905|Antidepressive Drugs, Second-Generation
C0242905|Atypical Antidepressants
C0085217|Carbonate, Lithium
C0085217|Lithium Carbonate
C0085217|Carbonate, Dilithium
C0085217|Carbonic acid, dilithium salt
C0085217|lithium carbonate (medication)
C0085217|Lithium Carbonate [Chemical/Ingredient]
C0085217|Dilithium Carbonate
C0085217|Lithium carbonate preparation
C0085217|Lithium carbonate (product)
C0085217|Lithium carbonate (substance)
C0003289|Agents, Antidepressive
C0003289|Antidepressive Agents
C0003289|antidepressant
C0003289|Drugs, Antidepressant
C0003289|ANTIDEPRESSANTS
C0003289|antidepressants (medication)
C0003289|Antidepressive
C0003289|Antidepressive Agent [TC]
C0003289|[CN600] ANTIDEPRESSANTS
C0003289|Antidepressive Agent
C0003289|Antidepressant drug
C0003289|Antidepressant drug (substance)
C0003289|Antidepressant Drugs
C0003289|Antidepressant (product)
C0003289|Antidepressant (substance)
C0003289|Antidepressant, NOS
C0003289|Antidepressant Agent
C1337136|l-methylfolate
C1337136|L-methylfolate (product)
C1337136|L-methylfolate (substance)
C1337136|6(S)-5-methyltetrahydrofolate
C1337136|L-methyl folic acid
C1337136|5-MTHF
C1337136|5-Methyltetrahydrofolate
C1337136|L-Glutamic Acid, N-(4-(((2-amino-1,4,5,6,7,8-hexahydro-5- methyl-4-oxo-6-pteridinyl)methyl)amino)benzoyl)-
C1337136|L-methyltetrahydrofolate
C1337136|5-Methyl terahydrofolic Acid
C2316497|Bupropion hydrobromide (substance)
C2316497|Bupropion hydrobromide
C2316497|1-Propanone, 1-(3-Chlorophenyl)-2-((1,1-dimethylethyl)amino)-, Hydrobromide
C2316497|bupropion HBr
C2316497|bupropion hydrobromide (medication)
C0215087|N,N-dimethyl-alpha-(2-(1-naphthalenyloxy)ethyl)benzenemethanamine
C0215087|dapoxetine
C0215087|Benzenemethanamine, N,N-dimethyl-alpha-(2-(1-naphthalenyloxy)ethyl)-, (+)-
C0215087|Dapoxetine (substance)
C2699580|Delfaprazine
C2699584|Delucemine Hydrochloride
C0957739|Eclanamine Maleate
C0068785|3-(2-methoxyphenoxy)-N-methyl-3-phenylpropylamine
C0068785|3-(o-methoxyphenoxy)-N-methyl-3-phenylpropylamine
C0068785|N-methyl-gamma-(2-methylphenoxy)phenylpropanolamine
C0068785|nisoxetine
C2698483|Nomelidine
C2698505|Noxiptiline
C0069709|2-(3-trifluoromethylphenyl)-4-isopropyltetrahydro-1,4-oxazine
C0069709|4-(1-methylethyl)-2-(3-(trifluoromethyl)phenyl)morpholine
C0069709|oxaflozane
C2699092|Rofelodine
C2699289|Seproxetine
C0069628|1,2,3,4-tetrahydro-2-methyl-9H-dibenzo(3,4-6,7)cyclohepta(1,2-C)pyridine
C0069628|13b,4a-carba-mianserin
C0069628|setiptiline
C2699506|Spiroxepin
C0144486|Talsupram
C2699901|Tebatizole
C0075496|sufoxazine
C0075496|teniloxazine
C2699942|Tienopramine
C0607615|tetrahydro-6-(phenoxymethyl)-2H-1,3-oxazine-2- thione
C0607615|tifemoxone
C0538554|(S)-2-(((7-fluoro-4-indanyl)oxy)methyl)morpholine monohydrochloride
C0538554|Lubazodone Hydrochloride
C0055961|(E)-1-(4- chlorophenyl)-5-methoxy-1-pentanone O-(2- aminoethyl)oxime, (E)-2-butenedioate (1:1)
C0055961|clovoxamine
C0600943|cotriptyline
C0600943|10,11-dihydro-5H-dibenzo(a,d)cycloheptenylidene-5-3-dimethylamino-2-propanone
C0663336|alpha-2-propenyl benzeneethanamine
C0663336|aletamine
C0663336|alfetadrine
C0663336|alfetamin
C0663336|alfetamine
C0663336|Alpha-Allyl-phenethylamin
C0663336|Alpha-Allylphenethylamine
C1702222|befetupitant
C2698343|Beloxepin
C0621294|clobamine mesylate
C0621294|Cilobamine Mesylate
C2699221|Cinfenine
C0047305|3-chloro-5-(3-(4-piperidino-4- carbamoylpiperidino)propyl)-10,11-dihydro-5H- dibenz(b,f)azepine dihydrochloride monohydrate
C0047305|3-chlorocarpipramine
C0047305|clocapramine
C2699359|Clodazon
C2699360|Clodazon Hydrochloride
C0615823|5H-dibenxo(a,d)cyclohepten-5-one O-(2-(methylamino)ethyl)oxime
C0615823|demexiptiline
C0044643|5-(3-(dimethylamino)propyl)-5H-dibenz- (b,f)azepine
C0044643|Depramine
C0044643|10,11-dehydroimipramine
C2699611|Deximafen
C0131796|(2-(2-dimethylamino)ethyl)-2-phenyl-3,4-dihydro-1(2H)-naphthalenone
C0131796|(S)-nafenodone
C0131796|nafenodone
C0131796|dexnafenodone
C0057877|diclofensine
C0543452|Hydrochloride, Dothiepin
C0543452|dothiepin hydrochloride (medication)
C0543452|dothiepin hydrochloride
C0543452|antidepressants dothiepin hydrochloride
C0543452|Dothiepin hydrochloride (product)
C0543452|Dothiepin hydrochloride (substance)
C0543452|Dosulepin hydrochloride
C2699861|Elanzepine
C2697947|Lubazodone
C1533126|Cyclopropanecarboxamide, 2-(aminomethyl)-N,N-diethyl-1-phenyl-, cis-(+-)-
C1533126|MILNACIPRAN
C1533126|Milnacipran (product)
C1533126|Milnacipran (substance)
C1533126|midalcipran
C1533126|milnacipran [Chemical/Ingredient]
C1533126|antidepressants snri milnacipran
C1533126|milnacipran (medication)
C0066529|milnacipran hydrochloride
C0066529|Milnacipran hydrochloride (product)
C0066529|Milnacipran hydrochloride (substance)
C0066529|milnacipran hydrochloride (medication)
C0066529|1-phenyl-1-diethylaminocarbonyl-2-aminomethylcyclopropane HCl
C2698946|Radafaxine Hydrochloride
C2699361|Clodazon Hydrochloride Anhydrous
C0052237|1,3,4,14b-tetrahydro-2-methyl-10H-pyrazino-(1,2-a)pyrrolo(2,1-c)(1,4)benzodiazepine
C0052237|aptazapine
C0052237|2H,10H-Parazino(1,2-a)pyrrolo(2,1-c)(1,4)benzodiazepine,1,3,4,14b-tetrahydro-2-methyl-
C2698177|Aptazapine Maleate
C2698177|2H,10H-Pyrazino(1,2-a)pyrrolo(2,1-c)(1,4)benzodiazepine, 1,3,4,14b-tetrahydro-2-methyl-, (+-)-, (Z)-2-butenedioate (1:1)
C2698082|2H- Indol-2-one, l,3-dihydro-3-methyl-3-[3-(methylamino)-propyl]-l-phenyl-
C2698082|Atext2phenotypein
C2607957|Benzaprinoxide
C2607957|1-Propanamine, 3-(1-chloro-5H-dibenzo(a,d)cyclohepten-5-ylidene)-N,N-dimethyl-, N-oxide
C2698511|Bipenamol
C0054270|10,11-dihydro-N,N,beta-trimethyl-5H-dibenzo(a,d) cycloheptane-5-propylamine
C0054270|butriptylene
C0054270|butriptyline
C0054270|10,11-Dihydro-N,N,beta-trimethyl-5H-dibenzo(a,d)cycloheptene-5-propylamine
C0054270|Butriptyline (product)
C0054270|Butriptyline (substance)
C1108795|butriptyline hydrochloride (medication)
C1108795|antidepressants butriptyline hydrochloride
C1108795|butriptyline hydrochloride
C1108795|5H-Dibenzo(a,d)cycloheptene-5-propylamine, 10,11-dihydro-N,N,beta-trimethyl-, Hydrochloride, DL-
C2699208|Ciclopramine
C2699208|2,3,7,8-Tetrahydro-3-methylamino-1H-chino(1,8-a,b)benzazepin
C2699343|3-(3-Chlorphenyl)-1-(dimethylamino)-3-phenyl-2-propanol
C2699343|Clemeprol
C2699343|m-Chloro-alpha-((dimethylamino)methyl)-beta-phenylphenetyl Alcohol
C0055708|ciclazindol
C0055708|Pyrimido(1,2-a)indol-10-ol, 10-(3-chlorophenyl)-2,3,4,10-tetrahydro-
C0951496|3-(2-morpholino-ethylamino)-4-methyl-6-phenyl pyridazine, dihydrochloride
C0951496|N-(4-Methyl-6-phenyl-3-pyridazinyl)-4-morpholineethanamine Dihydrochloride
C0951496|Minaprine Hydrochloride
C0951496|Morpholine, 4-(2-((4-methyl-6-phenyl-3-pyridazinyl)amino)ethyl)-, Dihydrochloride
C0951496|Minaprine Dihydrochloride
C0959897|Alpha-Allylphenethylamine Hydrochloride
C0959897|Alfetamine Hydrochloride
C0959897|Aletamine Hydrochloride
C0959897|Benzeneethanamine, alpha-2-propenyl-, Hydrochloride
C0970823|Dapoxetine Hydrochloride
C0621295|2-(3,4-dichlorophenyl)-3-((1-methylethyl)amino)bicyclo(2.2.2)octan-2-ol monomethanesulfonate
C0621295|cilobamine
C2825651|Atext2phenotypein Hydrochloride
C0953067|Indeloxazine Hydrochloride
C2825652|Dilopetine
C0635054|eclanamine
C2825653|Nuclotixene
C2825654|Adoprazine
C2825655|Caproxamine
C0063456|2-(7-indenyloxymethyl)morpholine
C0063456|indeloxazine
C0063456|Morpholine, 2-((1H-inden-7-yloxy)methyl)-
C0054826|5-(3-(4-piperidino-4-carbamoylpiperidino)propyl)- 10,11-dihydro-5(h)-dibenz(b,f)azepine
C0054826|carbadipimidine
C0054826|carpipramine
C2825656|Fenmetozole Hydrochloride
C0060175|fenmetazole
C0060175|fenmetozole
C0060175|2-((3,4-dichlorophenoxy)methyl)-2-imidazoline
C0056704|2,3,4,9-tetrahydro-N,N-dimethyl-1H-carbazol-3- amine
C0056704|2,3,4,9-tetrahydro-N,N-dimethyl-1H-carbazole-3-amine
C0056704|3-(dimethylamino)-1,2,3,4-tetrahydrocarbazole
C0056704|cyclindole
C2825657|Losindole
C0058199|dimetacrine
C0058199|dimethacrine
C0058199|isotonil
C0058199|istonil
C2825658|Lomevactone
C2825659|Fenmetramide
C2826066|Mariptiline
C2826066|1a,10b-Dihydrodibenzo(a,e)cyclopropa(c)cyclohepten-6(1H)-one O-(2-aminoethyl)oxime
C0886642|PAROXETINE HYDROCHLORIDE HEMIHYDRATE
C0886642|Paroxetine Hydrochloride, Hemihydrate
C0886642|Hemihydrate, Paroxetine Hydrochloride
C0886642|Hydrochloride Hemihydrate, Paroxetine
C0886642|Hydrochloride, Hemihydrate Paroxetine
C0886642|Hemihydrate Paroxetine Hydrochloride
C0886642|(3s-trans)-3-[(1,3-benzodioxol-5-yloxy)methyl]-4-(4-fluorophenyl)piperidine hydrochloride Hemihydrate
C2827083|Azepindole
C2827119|Cutamesine
C2827119|1-(2-(3,4-Dimethoxyphenyl)Ethyl)-4-(3-Phenylpropyl)Piperazine
C2827129|Dazadrol
C2827129|2-Pyridinemethanol, alpha-(4-Chlorophenyl)-alpha-(4,5-Dihydro-1H-Imidazol-2-yl)-
C2827129|alpha-(P-Chlorophenyl)-alpha-2-Imidazolin-2-yl-2-Pyridinemethanol
C2827130|Dazadrol Maleate
C2827154|Fantridone
C0963192|(+-)-trans-3-(3,4-Dichlorophenyl)-N-methyl-1-indanamine
C0963192|Indatraline
C0611882|5-(3-(dimethylamino)propyl)-5,11-dihydro-10H-dibenz(b,f)azepin-10-one
C0611882|ketimipramine
C0611882|ketipramine
C0611882|1-Alpha-4,5-Alpha-H-Tropanium, 3-Alpha-Hydroxy-8-(P-Phenylphenacyl)-, (-)-Tropate
C2827221|Ketipramine Fumarate
C0125662|levoprotiline
C0125662|hydroxymaprotilin, (+R)-isomer
C1565971|Talopram
C1565971|1,3-dihydro-N,3,3-trimethyl-1-phenylbenzo(c)furan-1-propanamine
C0025912|Mianserin
C0025912|Dibenzo(c,f)pyrazino(1,2-a)azepine, 1,2,3,4,10,14b-hexahydro-2-methyl-
C0025912|Mianserin [Chemical/Ingredient]
C0025912|1,2,3,4,10,14B-Hexahydro-2-Methyldibenzo(C,F)-Pyrazino(1,2-A)Azepine
C0025912|antidepressants mianserin
C0025912|mianserin (medication)
C0025912|Mianserin (product)
C0025912|Mianserin (substance)
C0700456|Hydrochloride, Mianserin
C0700456|mianserin hydrochloride (medication)
C0700456|mianserin hydrochloride
C0700456|antidepressants mianserin hydrochloride
C0700456|Dibenzo(C,F)Pyrazino(1,2-A)Azepine, 1,2,3,4,10,14B-Hexahydro-2-Methyl-, Monohydrochloride
C0700456|1,2,3,4,10,14B-Hexahydro-2-Methyldibenzo(C,F)-Pyrazino(1,2-A)Azepine Monohydrochloride
C0700456|Monohydrochloride, Mianserin
C0700456|Mianserin Monohydrochloride
C0700456|Mianserin hydrochloride (product)
C0700456|Mianserin hydrochloride (substance)
C0031974|pipradrol
C0031974|pyridrol
C0031974|pipradol
C0031974|Pipradrol (substance)
C0020934|Imipramine
C0020934|5H-Dibenz(b,f)azepine-5-propanamine, 10,11-dihydro-N,N-dimethyl-
C0020934|Imidobenzyle
C0020934|Imipramine [Chemical/Ingredient]
C0020934|Imizin
C0020934|Norchlorimipramine
C0020934|Imipramine (product)
C0020934|Imipramine (substance)
C0026388|Molindone
C0026388|4H-Indol-4-one, 3-ethyl-1,5,6,7-tetrahydro-2-methyl-5-(4-morpholinylmethyl)-
C0026388|Molindone [Chemical/Ingredient]
C0026388|Molindone (product)
C0026388|Molindone (substance)
C0040805|Trazodone
C0040805|1,2,4-Triazolo(4,3-a)pyridin-3(2H)-one, 2-(3-(4-(3-chlorophenyl)-1-piperazinyl)propyl)-
C0040805|Tradozone
C0040805|Searle Brand of Trazodone Hydrochloride
C0040805|Trazodone [Chemical/Ingredient]
C0040805|trazodone (medication)
C0040805|antidepressants trazodone
C0040805|Trazodone (product)
C0040805|Trazodone (substance)
C0038803|Sulpiride
C0038803|Benzamide, 5-(aminosulfonyl)-N-((1-ethyl-2-pyrrolidinyl)methyl)-2-methoxy-
C0038803|Sulpiride [Chemical/Ingredient]
C0038803|Sulperide
C0038803|N-((1-Ethyl-2-Pyrrolidinyl)Methyl)-5-Sulfamoyl-O-Anisamide
C0038803|antidepressants sulpiride
C0038803|sulpiride (medication)
C0038803|Sulpiride (product)
C0038803|Sulpiride (substance)
C0043479|Zimeldine
C0043479|2-Propen-1-amine, 3-(4-bromophenyl)-N,N-dimethyl-3-(3-pyridinyl)-, (Z)-
C0043479|Zimeldine [Chemical/Ingredient]
C0043479|Zimelidin
C0043479|Zimelidine
C0043479|Zimeldine (substance)
C0028420|Nortriptyline
C0028420|1-Propanamine, 3-(10,11-dihydro-5H-dibenzo(a,d)cyclohepten-5-ylidene)-N-methyl-
C0028420|Desitriptyline
C0028420|Nortriptyline [Chemical/Ingredient]
C0028420|Desmethylamitriptylin
C0028420|Nortriptyline (substance)
C0028420|Nortryptyline
C0028420|Nortriptyline (product)
C0028420|NTPL
C0025810|Methylphenidate
C0025810|2-Piperidineacetic acid, alpha-phenyl-, methyl ester
C0025810|alpha-Phenyl-2-piperidineacetic Acid Methyl Ester
C0025810|Methylphenidate [Chemical/Ingredient]
C0025810|methylphenidate (medication)
C0025810|cns stimulants methylphenidate
C0025810|Methylphenidate (product)
C0025810|Methylphenidate (substance)
C0025810|d-methylphenidate
C0031407|beta-phenylisopropylhydrazine
C0031407|pheniprazine
C0031407|Hydrazine, (1-methyl-2-phenylethyl)-
C0013085|Doxepin
C0013085|1-Propanamine, 3-dibenz(b,e)oxepin-11(6H)-ylidene-N,N-dimethyl-
C0013085|Doxepin [Chemical/Ingredient]
C0013085|Doxepin (product)
C0013085|Doxepin (substance)
C0024778|Maprotiline
C0024778|9,10-Ethanoanthracene-9(10H)-propanamine, N-methyl-
C0024778|Maprotilin
C0024778|N-Methyl-9,10-ethanoanthracene-9(10H)-propylamine
C0024778|Dibencycladine
C0024778|Maprotiline [Chemical/Ingredient]
C0024778|Maprotiline (product)
C0024778|Maprotiline (substance)
C0011685|Desipramine
C0011685|5H-Dibenz(b,f)azepine-5-propanamine, 10,11-dihydro-N-methyl-
C0011685|Desmethylimipramine
C0011685|Demethylimipramine
C0011685|Desipramine [Chemical/Ingredient]
C0011685|antidepressants desipramine
C0011685|desipramine (medication)
C0011685|Desipramine (product)
C0011685|Desipramine (substance)
C0009010|Clomipramine
C0009010|5H-Dibenz(b,f)azepine-5-propanamine, 3-chloro-10,11-dihydro-N,N-dimethyl-
C0009010|3-Chloro-5-(3-(dimethylamino)propyl)-10,11-dihydro-5H-dibenz(b,f)azepine
C0009010|Chlomipramine
C0009010|Clomipramine [Chemical/Ingredient]
C0009010|Chlorimipramine
C0009010|Clomipramine (substance)
C0009010|Clomipramine (product)
C0028277|Nomifensine
C0028277|8-Isoquinolinamine, 1,2,3,4-tetrahydro-2-methyl-4-phenyl-
C0028277|Nomifensin
C0028277|Linamiphen
C0028277|Nomifensine [Chemical/Ingredient]
C0009170|Cocaine
C0009170|8-Azabicyclo(3.2.1)octane-2-carboxylic acid, 3-(benzoyloxy)-8-methyl-, methyl ester, (1R-(exo,exo))-
C0009170|(1R,2R,3S,5S)-2-Methoxycarbonyltropan-3-yl Benzoate
C0009170|Cocaine [Chemical/Ingredient]
C0009170|cocaine (Schedule I substance)
C0009170|Blow
C0009170|C
C0009170|Snow
C0009170|Coke
C0009170|Coca
C0009170|Cocaine product
C0009170|Cocaine (product)
C0009170|Cocaine (substance)
C0355303|Compound antidepressants
C0355303|Compound antidepressants (product)
C0355303|Compound antidepressants (substance)
C0771200|Venlafaxine Hydrochloride
C0771200|venlafaxine hydrochloride (medication)
C0771200|antidepressants venlafaxine hydrochloride
C0771200|Hydrochloride, Venlafaxine
C0771200|Cyclohexanol, 1-(2-(dimethylamino)-1-(4-methoxyphenyl)ethyl)-, hydrochloride
C0771200|Venlafaxine Hydrochloride [Chemical/Ingredient]
C0771200|1-(2-(dimethylamino)-1-(4-methoxyphenyl)ethyl)cyclohexanol HCl
C0771200|Venlafaxine hydrochloride (substance)
C0771200|Venlafaxine hydrochloride (product)
C0600356|H 102 09
C0600356|H10209
C0600356|H-102-09
C0002600|Amitriptyline
C0002600|1-Propanamine, 3-(10,11-dihydro-5H-dibenzo(a,d)cyclohepten-5-ylidene)-N,N-dimethyl-
C0002600|Amitriptyline [Chemical/Ingredient]
C0002600|Amitriptyline (product)
C0002600|Amitriptyline (substance)
C0678139|Seroxat
C0591911|Optimax
C0591911|Merck Brand of Tryptophan
C0360105|selective serotonin reuptake inhibitors (medication)
C0360105|serotonin reuptake inhibitors
C0360105|selective serotonin reuptake inhibitors (SSRIs)
C0360105|selective serotonin reuptake inhibitors
C0360105|Selective Serotonin Reuptake Inhibitor
C0360105|SSRIs
C0360105|SSRI
C0360105|SSRI - Selective serotonin re-uptake inhibitor
C0360105|Selective serotonin re-uptake inhibitor
C0360105|Selective serotonin re-uptake inhibitor (product)
C0360105|Selective serotonin re-uptake inhibitor (substance)
C0543469|viloxazine hydrochloride (medication)
C0543469|antidepressants viloxazine hydrochloride
C0543469|viloxazine hydrochloride
C0543469|Viloxazine hydrochloride (product)
C0543469|Viloxazine hydrochloride (substance)
C1529955|antidepressants dibenzepin hydrochloride
C1529955|dibenzepin hydrochloride
C1529955|dibenzepin hydrochloride (medication)
C0877847|Maleate, Nomifensine
C0877847|nomifensine maleate (medication)
C0877847|nomifensine maleate
C0877847|Nomifensine Maleate (1:1)
C2079567|perphenazine + nortriptyline (medication)
C2079567|perphenazine + nortriptyline
C2079567|Nortriptyline / Perphenazine
C2189302|veralipride + bromazepam
C2189302|veralipride + bromazepam (medication)
C2189302|Bromazepam / veralipride
C0041056|Trimipramine
C0041056|5H-Dibenz(b,f)azepine-5-propanamine, 10,11-dihydro-N,N,beta-trimethyl-
C0041056|trimipramine (medication)
C0041056|Trimeprimine
C0041056|10,11 Dihydro-N,N,beta-trimethyl-5H-dibenz(b,f)azepine-5-propanamine
C0041056|Trimipramine [Chemical/Ingredient]
C0041056|Trimipramine (product)
C0041056|Trimipramine (substance)
C0036579|Selegiline
C0036579|Benzeneethanamine, N,alpha-dimethyl-N-2-propynyl-, (R)-
C0036579|selegiline (medication)
C0036579|(-)-Deprenil
C0036579|(-)-Phenylisopropylmethylpropynylamine
C0036579|L-Deprenyl
C0036579|Selegiline [Chemical/Ingredient]
C0036579|Selegyline
C0036579|Selegiline, (R)-Isomer
C0036579|(-)-Selegiline
C0036579|Selegiline (product)
C0036579|Selegiline (substance)
C1579361|SNRI antidepressants
C1579361|Serotonin and Norepinephrine Reuptake Inhibitors (SNRIs)
C1579361|serotonin and norepinephrine reuptake inhibitors (medication)
C1579361|antidepressants serotonin and norepinephrine reuptake inhibitors
C1579361|serotonin and norepinephrine reuptake inhibitors
C1579361|Serotonin and Noradrenaline Reuptake Inhibitors
C1579361|NRIs and SSRIs
C1579361|Serotonin and Norepinephrine Uptake Inhibitors
C1579361|SSRIs and NRIs
C1579361|Serotonin and Noradrenaline Uptake Inhibitors
C1579361|SNRIs
C2064901|benactyzine hydrochloride + meprobamate
C2064901|benactyzine hydrochloride + meprobamate (medication)
C1616289|hydrogenated ergot alkaloids (medication)
C1616289|hydrogenated ergot alkaloids
C1616289|Ergot Alkaloids, Hydrogenated
C1616289|Hydrogenated ergot alkaloid
C1616289|Alkaloids, Hydrogenated Ergot
C0026457|Inhibitor, Monoamine Oxidase
C0026457|Inhibitors, Monoamine Oxidase
C0026457|Monoamine Oxidase Inhibitors
C0026457|MAO inhibitor
C0026457|Inhibitors, MAO
C0026457|MAO INHIB
C0026457|MONOAMINE OXIDASE INHIB
C0026457|monoamine oxidase inhibitor
C0026457|monoamine oxidase inhibitors (medication)
C0026457|MAO inhibitors
C0026457|monoamine oxidase inhibitors (MAOI)
C0026457|MAOI
C0026457|Monoamine oxidase--Inhibitors
C0026457|MAOI - Monoamine-oxidase inhibitor
C0026457|Monoamine-oxidase inhibitor
C0026457|Monoamine oxidase inhibitor (product)
C0026457|Monoamine oxidase inhibitor (substance)
C0026457|Monoamine oxidase inhibitor, NOS
C0026457|Amine Oxidase Inhibitors
C1302097|perphenazine + amitriptyline hydrochloride (medication)
C1302097|perphenazine + amitriptyline hydrochloride
C1302097|antidepressants perphenazine + amitriptyline HCl
C1302097|Amitriptyline hydrochloride + perphenazine
C1302097|Amitriptyline hydrochloride + perphenazine (product)
C0002644|Amoxapine
C0002644|Dibenz(b,f)(1,4)oxazepine, 2-chloro-11-(1-piperazinyl)-
C0002644|amoxapine (medication)
C0002644|Amoxapine [Chemical/Ingredient]
C0002644|Desmethylloxapine
C0002644|2-Chloro-11-(1-piperazinyl)dibenz(b,f)(1,4)oxazepine
C0002644|Amoxapine - chemical
C0002644|Amoxapine - chemical (substance)
C0002644|Amoxapine (product)
C0002644|Amoxapine (substance)
C0049506|6-azamianserin
C0049506|Pyrazino(2,1-a)pyrido(2,3-c)(2)benzazepine, 1,2,3,4,10,14b-hexahydro-2-methyl-
C0049506|mirtazapine
C0049506|mirtazapine (medication)
C0049506|mirtazapine [Chemical/Ingredient]
C0049506|Mirtazapine (product)
C0049506|Mirtazapine (substance)
C1875508|MONAMINE OXIDASE INHIBITOR ANTIDEPRESSANTS
C1875508|[CN602] MONAMINE OXIDASE INHIBITOR ANTIDEPRESSANTS
C1579362|ANTIDEPRESSANTS,OTHER
C1579362|[CN609] ANTIDEPRESSANTS,OTHER
C2981302|MO-1255
C2981302|Encyprate
C2981302|Carbamic Acid, Cyclopropyl(Phenylmethyl)-, Ethyl Ester
C2981302|Ethyl N-Benzylcyclopropanecarbamate
C2981302|A-19757
C2981303|Esreboxetine Succinate
C2981304|Fantridone Hydrochloride Anhydrous
C2981304|5-(3-(Dimethylamino)Propyl)-6(5H)-Phenanthridinone Monohydrochloride
C2981304|6(5H)-Phenanthridinone, 5-(3-(Dimethylamino)Propyl)-, Monohydrochloride
C0023961|Lofepramine
C0023961|Ethanone, 1-(4-chlorophenyl)-2-((3-(10,11-dihydro-5H-dibenz(b,f)azepin-5-yl)propyl)methylamino)-
C0023961|Lofepramine [Chemical/Ingredient]
C0023961|Lopramine
C0023961|4'-Chloro-2-((3-(10,11-Dihydro-5H-Dibenz(b,f)azepin-5-yl)Propyl)Methylamino)Acetophenone
C0023961|Lofepramine (product)
C0023961|Lofepramine (substance)
C0023330|Hydrochloride, Lofepramine
C0023330|antidepressants lofepramine hydrochloride
C0023330|lofepramine hydrochloride
C0023330|lofepramine hydrochloride (medication)
C0023330|Lofepramine hydrochloride (substance)
C0023330|4'-Chloro-2-((3-(10,11-Dihydro-5H-Dibenz(b, f)azepin-5-yl)Propyl)Methylamino)acetophenone Monohydrochloride
C0023330|Ethanone, 1-(4-Chlorophenyl)-2-((3-(10,11-Dihydro-5H-Dibenz(b, f)azepin-5-yl)Propyl)Methylamino)-, Monohydrochloride
C0066057|15-methyl-10-methylamino-10,11- dihydrodibenzo(b,f)-azepine
C0066057|metapramine
C0066057|15-methyl-10-methylamino-10,11-dihydrodibenzo(b,f)- azepine
C0066057|10,11-Dihydro-5-Methyl-10-(Methylamino)-5H-Dibenz(B,F)Azepine
C0029105|Opipramol
C0029105|1-Piperazineethanol, 4-(3-(5H-dibenz(b,f)azepin-5-yl)propyl)-
C0029105|Opipramol [Chemical/Ingredient]
C2983799|Orvepitant
C2983799|1-Piperidinecarboxamide, N-[(1R)-1-[3,5-bis(trifluoromethyl)phenyl]ethyl]-2-(4-fluoro-2-methylphenyl)-4-[(8aS)-hexahydro-6-oxopyrrolo[1,2-a]pyrazin-2(1H)-yl]-N-methyl-, (2R,4S)-
C2983800|GW823296B
C2983800|Orvepitant Maleate
C2983846|Melitracen Hydrochloride
C2983846|U 24,973A
C2983847|Modaline Sulfate
C2983847|W 3207B
C2983848|Naprodoxime
C2983849|Nemifitide
C2983850|Nitrafudam
C2983851|Omiloxetine
C1530072|vilazodone
C1530072|5-{4-[4-(5-cyano-1H-indol-3-yl)butyl]piperazin-1-yl}benzofuran-2-carboxamide
C1530072|Vilazodone (substance)
C1530072|5-(4-(4-(5-cyano-3-indolyl)butyl)-1-piperazinyl)benzofuran-2-carboxamide
C2962546|vilazodone hydrochloride
C2962546|5-{4-[4-(5-cyano-1H-indol-3-yl)butyl]piperazin-1-yl}benzofuran-2-carboxamide Hydrochloride
C2962546|antidepressants vilazodone
C2962546|vilazodone HCl (medication)
C2962546|vilazodone HCl
C2962546|Vilazodone hydrochloride (substance)
C2962546|HCl, Vilazodone
C2962546|Hydrochloride, Vilazodone
C2962546|2-benzofurancarboxamide, 5-(4-(4-(5-cyano-1H-indol-3-yl)butyl)-1-piperazinyl)-, hydrochloride (1:1)
C2962546|Vilazodone Hydrochloride [Chemical/Ingredient]
C2698285|Azaloxan
C0282270|Hydrochloride, Opipramol
C0282270|Opipramol Hydrochloride
C0282270|Opipramol Dihydrochloride
C0282270|4-(3-(5H-Dibenz(b,f)azepin-5-yl)Propyl)-1-Piperazineethanol Dihydrochloride
C0282270|1-Piperazineethanol, 4-(3-(5H-Dibenz(B,F)Azepin-5-yl)Propyl)-, Dihydrochloride
C0732706|lithium succinate 80 MG/ML Topical Cream
C0732706|lithium succinate 8 % Topical Cream
C0732706|Lithium succinate 8% cream
C0732706|Lithium succinate 8% cream (product)
C0732706|Lithium succinate 8% cream (substance)
C0013065|Dothiepin
C0013065|1-Propanamine, 3-dibenzo(b,e)thiepin-11(6H)-ylidene-N,N-dimethyl-
C0013065|Dothiepin [Chemical/Ingredient]
C0013065|Dosulepin
C0013065|Dothiepin (product)
C0013065|Dothiepin (substance)
C0013065|Dosulepin (substance)
C0973506|Other antidepressant drugs (product)
C0973506|Other antidepressant drugs
C0973506|Other antidepressant drugs (substance)
C0693279|BUPROPION HCL 100MG SA TAB
C0693279|BUPROPION HCL 100MG TAB,SA
C0693279|BUPROPION HCL 100MG TAB,SA [VA Product]
C0693279|buPROPion Hydrochloride 100 MG Extended Release Oral Tablet
C0693279|Bupropion hydrochloride 100mg m/r tablet (product)
C0693279|Bupropion hydrochloride 100mg m/r tablet
C0162758|Serotonin Uptake Inhibitors
C0162758|5 HT Uptake Inhibitors
C0162758|5 Hydroxytryptamine Uptake Inhibitors
C0162758|Inhibitors, 5 HT Uptake
C0162758|Inhibitors, 5 Hydroxytryptamine Uptake
C0162758|Uptake Inhibitors, 5 HT
C0162758|Uptake Inhibitors, 5 Hydroxytryptamine
C0162758|serotonin inhibitor
C0162758|HT 05 UPTAKE INHIBITORS
C0162758|SEROTONIN UPTAKE INHIB
C0162758|5 HT UPTAKE INHIB
C0162758|SEROTONIN REUPTAKE INHIB
C0162758|INHIB 5 HYDROXYTRYPTAMINE UPTAKE
C0162758|HYDROXYTRYPTAMINE UPTAKE INHIBITORS 05
C0162758|UPTAKE INHIB SEROTONIN
C0162758|INHIB 5 HT UPTAKE
C0162758|UPTAKE INHIB 5 HT
C0162758|5 HYDROXYTRYPTAMINE UPTAKE INHIB
C0162758|REUPTAKE INHIB SEROTONIN
C0162758|INHIB SREOTONIN REUPTAKE
C0162758|UPTAKE INHIB 5 HYDROXYTRYPTAMINE
C0162758|INHIB SEROTONIN UPTAKE
C0162758|serotonin reuptake inhibitor
C0162758|Serotonin uptake inhibitor (substance)
C0162758|Serotonin uptake inhibitor
C0162758|Serotonin uptake inhibitor (product)
C0162758|Uptake Inhibitors, 5-HT
C0162758|Serotonin Reuptake Inhibitors
C0162758|Uptake Inhibitors, 5-Hydroxytryptamine
C0162758|Uptake Inhibitors, Serotonin
C0162758|Inhibitors, 5-Hydroxytryptamine Uptake
C0162758|Inhibitors, 5-HT Uptake
C0162758|5-Hydroxytryptamine Uptake Inhibitors
C0162758|Inhibitors, Serotonin Reuptake
C0162758|Reuptake Inhibitors, Serotonin
C0162758|5-HT Uptake Inhibitors
C0162758|Inhibitors, Serotonin Uptake
C0162758|Serotonin uptake inhibitor, NOS
C0486980|Hydroxybupropion
C0486980|4-hydroxy bupropion
C0486980|Hydroxybupropion (substance)
C0068485|nefazodone
C0068485|nefazodone [Chemical/Ingredient]
C0068485|Nefazodone (product)
C0068485|Nefazodone (substance)
C0358139|lithium succinate 0.08 MG/MG Topical Ointment
C0358139|lithium succinate 8 % Topical Ointment
C0358139|Lithium succinate 8% ointment
C0358139|Lithium succinate 8% ointment (product)
C0358139|Lithium succinate 8% ointment (substance)
C0245561|duloxetine
C0245561|selective norepinephrine reuptake inhibitors duloxetine
C0245561|duloxetine (medication)
C0245561|N-methyl-3-(1-naphthalenyloxy)-3-(2-thiophene)propanamide
C0245561|N-methyl-3-(1-naphthalenyloxy)-2-thiophenepropanamine
C0245561|Duloxetine (product)
C0245561|Duloxetine (substance)
C0304364|Bicyclic antidepressant (substance)
C0304364|Bicyclic antidepressant
C0304364|Bicyclic antidepressant, NOS
C0700535|Doxepin Hydrochloride
C0700535|Hydrochloride, Doxepin
C0700535|Doxepin Hydrochloride [Chemical/Ingredient]
C0700535|Doxepin Hydrochloride, Cis-Trans Isomer Mixture (approximately 1:5)
C0700535|Doxepin hydrochloride [antipruritic] (product)
C0700535|Doxepin hydrochloride (product)
C0700535|Doxepin hydrochloride [antipruritic]
C0700535|antidepressants doxepin hydrochloride
C0700535|antipruritics doxepin hydrochloride
C0700535|antipruritics doxepin hydrochloride (medication)
C0700535|antidepressants doxepin hydrochloride (medication)
C0700535|Doxepin hydrochloride (substance)
C0700535|Doxepin hydrochloride [antipruritic] (substance)
C1289960|O-Desmethyvenlafaxine (substance)
C1289960|O-Desmethyvenlafaxine
C3650301|antidepressants maprotiline (medication)
C3650301|antidepressants maprotiline
C3650306|antidepressants escitalopram
C3650306|antidepressants escitalopram (medication)
C2936679|flupentixol, melitracen drug combination
C2936679|flupentixol - melitracen
C2936679|flupentixol + melitracen (medication)
C2936679|flupentixol + melitracen
C2936679|antidepressants flupentixol + melitracen
C3650307|antidepressants dothiepin
C3650307|antidepressants dothiepin (medication)
C0971637|Agomelatine
C0971637|Agomelatine (substance)
C0971637|Agomelatine (product)
C1993532|Nomifensine &#x7C; bld-ser-plas
C1099456|Escitalopram
C1099456|S(+)-Citalopram
C1099456|(S)-Citalopram
C1099456|Escitalopram (product)
C1099456|Escitalopram (substance)
C0074493|sibutramine
C0074493|sibutramine [Chemical/Ingredient]
C0074493|Sibutramine product (product)
C0074493|Sibutramine product
C0074493|Sibutramine (product)
C0074493|Sibutramine (substance)
C1981553|Antidepressants &#x7C; gastric fluid
C1972481|Reboxetine &#x7C; Bld-Ser-Plas
C1981554|Antidepressants &#x7C; urine
C1975864|Zimelidine &#x7C; bld-ser-plas
C1992738|Moclobemide &#x7C; bld-ser-plas
C1994490|Phenelzine &#x7C; bld-ser-plas
C1981552|Antidepressants &#x7C; bld-ser-plas
C0072127|1-(alpha-propylphenethyl)pyrrolidine
C0072127|phenylpyrrolidinylpentan
C0072127|prolintane
C0072127|Prolintane (product)
C0072127|Prolintane (substance)
C0076652|(3-chloro-6-methyl-5,5-dioxo-6,11-dihydrodibenzo(c,f)(1,2)thiazepin-11-yl)-7-aminoheptanoic acid
C0076652|tianeptine
C0076652|Tianeptine (substance)
C3847513|Vilazodone &#x7C; Urine
C0040098|Thymoleptics
C0040094|Thymoanaleptics
C0771509|tianeptine sodium
C0771509|tianeptine sodium (medication)
C0771509|Tianeptine sodium (substance)
C4038278|Citalopram+Escitalopram &#x7C; Urine
C3661282|vortioxetine
C3661282|1-(2-(2,4-dimethylphenylsulfanyl)phenyl)piperazine
C3661282|antidepressants vortioxetine
C3661282|vortioxetine (medication)
C3661282|Vortioxetine (substance)
C1742884|Desvenlafaxine Succinate
C1742884|Desvenlafaxine succinate (substance)
C1742884|desvenlafaxine succinate (medication)
C1742884|Butanedioic Acid, Compound With 4-(2-(Dimethylamino)-1-(1-Hydroxycyclohexyl)Ethyl)Phenol (1:1), Monohydrate
C1742884|Succinate Monohydrate, O-desmethylvenlafaxine
C1742884|Monohydrate, O-desmethylvenlafaxine Succinate
C1742884|O desmethylvenlafaxine Succinate Monohydrate
C1742884|Succinate, Desvenlafaxine
C1742884|O desmethylvenlafaxine Succinate
C1742884|Succinate, O-desmethylvenlafaxine
C1742884|O-desmethylvenlafaxine Succinate Monohydrate
C1742884|O-desmethylvenlafaxine Succinate
C1742884|Desvenlafaxine Succinate [Chemical/Ingredient]
C1742884|2-(1-hydroxycyclohexyl)-2-((4-hydroxyphenyl)ethyl)dimethylammonium 3-carboxypropanoate monohydrate
C1505020|Duloxetine hydrochloride
C1505020|Duloxetine hydrochloride (substance)
C1505020|duloxetine hydrochloride (medication)
C1505020|Hydrochloride, Duloxetine
C1505020|HCl, Duloxetine
C1505020|Duloxetine Hydrochloride [Chemical/Ingredient]
C1505020|Duloxetine HCl
C2980164|Gaboxetine KIT
C2980164|Gaboxetine Convenience Pack
C2980164|Acetylcarnitine/Choline Bitartrate/Cocoa Extract/Gamma Aminobutyric Acid/Ginkgo Biloba Leaf/Glutamic Acid/Grape Seed Extract/Griffonia Seed Extract/Valerian Root Extract/Whey Protein Hydrolysate;Fluoxetine Hydrochloride 62.5 MG; 10 MG Oral Capsule [GABOXETINE]
C0041249|L Tryptophan
C0041249|Tryptophan
C0041249|L-Tryptophan
C0041249|L-tryptophan (medication)
C0041249|Levotryptophan
C0041249|Tryptophan [Chemical/Ingredient]
C0041249|L-Tryptophan (substance)
C0041249|Trp
C0041249|(S)-2-Amino-3-(1H-indol-3-yl)-propanoic acid
C0041249|Tryptophan product
C0041249|L-Tryptophan (product)
C0041249|Tryptophan (substance)
C0023870|Lithium
C0023870|Lithium product
C0023870|lithium (medication)
C0023870|Lithium [Chemical/Ingredient]
C0023870|Lithium Metallicum
C0023870|Li
C0023870|Li element
C0023870|Li+ element
C0023870|Li - Lithium
C0023870|Lithium (product)
C0023870|Lithium (substance)
C0023870|Lithium, NOS
C0023870|Lithium product (product)
C0023870|Lithium product (substance)
C0042665|Viloxazine
C0042665|Morpholine, 2-((2-ethoxyphenoxy)methyl)-
C0042665|Viloxazine [Chemical/Ingredient]
C0042665|Viloxazine (product)
C0042665|Viloxazine (substance)
C0168388|reboxetine
C0168388|reboxetine [Chemical/Ingredient]
C0168388|selective norepinephrine reuptake inhibitors reboxetine
C0168388|reboxetine (medication)
C0168388|Reboxetine (product)
C0168388|Reboxetine (substance)
C0360108|Tetracyclic antidepressant
C0360108|Tetracyclic antidepressant drug
C0360108|Tetracyclic antidepressant (product)
C0360108|Tetracyclic antidepressant (substance)
C0360108|Tetracyclic antidepressant, NOS
C1271027|Triazolopyridine
C1271027|Triazolopyridine (substance)
C1271027|Triazolopyridine (product)
C0012035|Dibenzothiepins
C0012035|Dibenzothiepins [Chemical/Ingredient]
C0012035|Dibenzothiepin
C0012035|Dibenzothiepin (substance)
C0063220|1,3,4,6,8,13-hexahydroxy-10,11-dimethylphenanthro(1,10,9,8-opqra)perylene-7,14-dione
C0063220|hypericin
C0063220|4,5,7,4',5',7'-Hexahydroxy-2,2'-dimethyl-mesonapthtodianthron
C0063220|Hypericin (substance)
C0066561|3-(morpholinoethyl)amino-4-methyl-6-phenylpyridazine
C0066561|minaprine
C0066561|N-(4-methyl-6-phenyl-3-pyridazinyl)-4-morpholineethanamine
C0066561|4-Morpholineethanamine, N-(4-methyl-6-phenyl-3-pyridazinyl)-
C0074500|mesocarb
C0074500|N-phenylcarbamoyl-3-(beta-phenylisopropyl)sydnonimine
C0074500|sidnocarb
C0074500|sydnocarb
C0071143|1,10-trimethylene-8-methyl-1,2,3,4-tetrahydropyrazino(1,2-a)indole
C0071143|1H-Pyrazino(3,2,1-jk)carbazole, 2,3,3a,4,5,6-hexahydro-8-methyl-, monohydrochloride
C0071143|pirlindol
C0071143|pirlindole
C0071143|pyrlindole
C0060145|femoxetine
C0060145|femoxitine
C0060145|Piperidine, 3-((4-methoxyphenoxy)methyl)-1-methyl-4-phenyl-, (3R-trans)-
C0060145|trans-(+)-3-((4-methoxyphenoxy)methyl)-1-methyl-4-phenylpiperidine
C0060145|trans-3-((4-methoxyphenoxy)methyl)-1-methyl-4-phenylpiperidine
C0076804|(3-methyl)-3-phenyl-5-hydroxymethyl-2-oxazolidinone
C0076804|5-(hydroxymethyl)-3-(3-methylphenyl)-2- oxazolidinone
C0076804|toloxatone
C0076804|5-(Hydroxymethyl)-3-(3-methylphenyl)-2-oxazolidinone
C0076804|5-Hydroxymethyl-3-(m-tolyl)-2-oxazolidinone
C0076784|1-(3,4-dimethoxyphenyl)-5-ethyl-7,8-dimethoxy- 4-methyl-5H-2,3-benzodiazepine
C0076784|tofisopam
C0076784|tofizopam
C0076784|1-(3,4-dimethoxyphenyl)-5-ethyl-7,8-dimethoxy-4-methyl-5H-2,3-benzodiazepine
C0069039|3-(4-bromophenyl)-N-methyl-(3-pyiidyl)allylamine oxalate
C0069039|norzimeldine
C0069039|norzimelidine
C0072076|Butanamide, 4-(((4-chlorophenyl)(5-fluoro-2-hydroxyphenyl)methylene)amino)-
C0072076|progabide
C0063448|(3-indolyl-2-ethyl)piperidine
C0063448|1H-Indole, 3-(2-(4-piperidinyl)ethyl)-
C0063448|4-(2-(3-indolyl)ethyl)piperidine
C0063448|indalpine
C0043636|(des-Tyr(1))-gamma-endorphin
C0043636|1-de-Tyr-gamma-endorphin
C0043636|beta-lipotropin(62-77)
C0043636|beta-LPH(62-77)
C0043636|DTgammaE
C0043636|gamma-endorphin, des-Tyr(1)-
C0043636|gamma-endorphin, des-tyrosine(1)-
C0139500|pyro(l-alpha-aminoadipyl)-L-histidyl-L-thiazolidine-4-carboxamide
C0139500|pyro-Aad-His-Tzl-NH2
C0139500|pyro-2-aminoadipylhistidylthiazolidine-4-carboxyamide
C0139500|(2S)-N-((2S)-1-((4S)-4-Carbamoyl-1,3-thiazolidin-3-yl)-3-(1H-imidazol-5-yl)-1-oxo-2-propanyl)-6-oxo-2-piperidinecarboxamide
C0075784|2-amino-6-allyl-5,6,7,8-tetrahydro-4H-thiazolo-(5,4-d)azepin-dihydrochloride
C0075784|4H-Thiazolo(4,5-d)azepin-2-amine, 5,6,7,8-tetrahydro-6-(2-propenyl)-, dihydrochloride
C0075784|talipexole
C0075784|6-allyl-2-amino-5,6,7,8-tetrahydro-4H-thiazolo(4,5-d)azepin dihydrochloride
C0051086|alaproclate
C0051086|DL-Alanine, 2-(4-chlorophenyl)-1,1-dimethylethyl ester
C0063159|hydroxymaprotilin
C0063159|oxaprotiline
C0106291|1-Butanamine, N-methyl-4-(2-(phenylmethyl)phenoxy)-, hydrochloride
C0106291|2-(4-methylaminobutoxy)diphenylmethane
C0106291|4-(2-benzylphenoxy)-N-methylbutylamine
C0106291|bifemelane
C0051917|1-(4-methoxybenzoyl)-2-pyrrolidinone
C0051917|1-anisoyl-2-pyrrolidinone
C0051917|aniracetam
C0050844|adinazolam
C0066624|4,4-dimethyl-1-(4-(4-(2-pyrimidinyl)-1-piperazinyl)butyl)-2,6-piperidinedione
C0066624|gepirone
C0075591|sulforidazine
C0060454|flesinoxan
C0060454|p-fluoro-N-(2-(4-(2-(hydroxymethyl)-1,4-benzodioxan-5-yl)-1-piperazinyl)ethyl)benzamide
C0299772|L 701,324
C0299772|L 701324
C0299772|L-701,324
C0299772|L-701324
C1445647|Phenylpiperazine antidepressant (substance)
C1445647|Phenylpiperazine antidepressant
C0303506|Lithium and its derivatives
C0303506|Lithium AND/OR lithium compound (substance)
C0303506|Lithium AND/OR lithium compound
C1881039|Hepzidine
C1880846|Fosenazide
C0123216|ifoxetine
C0600526|Sertraline Hydrochloride
C0600526|Hydrochloride, Sertraline
C0600526|sertraline hydrochloride (medication)
C0600526|antidepressants sertraline hydrochloride
C0600526|Sertraline Hydrochloride (1S-cis)-Isomer
C0600526|Sertraline Hydrochloride [Chemical/Ingredient]
C0600526|Sertraline hydrochloride (substance)
C0600526|Sertraline hydrochloride (product)
C1881247|Intriptyline
C1831797|casopitant mesylate
C0060394|fipexide
C0733380|fluoxetine hydrochloride
C0733380|antidepressants fluoxetine hydrochloride
C0733380|fluoxetine hydrochloride (medication)
C0733380|Fluoxetine Hydrochloride [Chemical/Ingredient]
C0733380|FLUoxetine HCl
C0733380|Fluoxetine hydrochloride (substance)
C0733380|Fluoxetine hydrochloride [dup] (substance)
C1880764|Feprosidnine
C1881816|Mezepine
C0526501|4-amino-5-chloro-2-ethoxy-N-((4-(4-fluorobenzyl)-2-morpholinyl)methyl)benzamide
C0526501|Benzamide, 4-amino-5-chloro-2-ethoxy-N-((4-((4-fluorophenyl)methyl)-2-morpholinyl)methyl)-, 2-hydroxy-1,2,3-propanetricarboxylate (1:1)
C0526501|mosapride
C1881248|Intriptyline Hydrochloride
C1873234|Tesofensine
C1881896|Monometacrine
C1880560|Etacepride
C1881131|Imafen Hydrochloride
C1880288|Desvenlafaxine
C1880288|Desvenlafaxine (product)
C1880288|Desvenlafaxine (substance)
C1880288|O desmethylvenlafaxine
C1880288|4-(2-(dimethylamino)-1-(1-hydroxycyclohexyl)ethyl)phenol
C1880288|O-desmethylvenlafaxine
C1880733|Fantridone Hydrochloride
C0065963|mepiprazole
C0070047|1-benzoyl-3-(1-(2-naphthylmethyl)-4-piperidyl)urea
C0070047|panuramine
C1881414|Litracen
C1880857|Ftorpropazine
C0165077|4-(2-naphthalenylmethoxy)piperidine
C0165077|litoxetine
C1881811|Metoxepin
C0066473|1H-3,4,6a-triazafluoranthene, 2,4,5,6-tetrahydro-9-methoxy-4-methyl-
C0066473|3-methyl-8-methoxy-(3H)-1,2,5,6-tetrahydropyrazino(1,2,3-ab)-beta-carboline
C0066473|metralindole
C0117861|flerobuterol
C1365510|Paroxetine Mesylate
C1365510|Paroxetine Methanesulfonate
C1365510|Piperidine, 3-((1,3-benzodioxol-5-yloxy)methyl)-4-(4-fluorophenyl)-,(3S,4R)-, Methanesulfonate
C1365510|Paroxetine mesylate (substance)
C1365510|paroxetine mesylate (medication)
C1365510|(-)-(3S,4R)-4-(p-Fluorophenyl)-3-((3,4-(methylenedioxy)phenoxy)methyl)piperidine Mesylate
C1365510|Paroxetine mesilate
C1882438|Prazepine
C1881288|Ivoqualine
C0078842|4-(3-chlorophenyl)-1,6,7,8-tetrahydro-1,3-dimethylpyrazolo(3,4-e)(1,4)diazepine
C0078842|zometapine
C0700563|Bupropion Hydrochloride
C0700563|(+-)-1-(3-Chlorophenyl)-2-[(1,1-dimethylethyl)amino]-1-propanone Hydrochloride
C0700563|antidepressants bupropion hydrochloride
C0700563|bupropion hydrochloride (medication)
C0700563|Bupropion Hydrochloride [Chemical/Ingredient]
C0700563|Bupropion hydrochloride (substance)
C0700563|Bupropion hydrochloride (product)
C1170741|Atomoxetine Hydrochloride
C1170741|(-)-N -Methyl-3-phenyl-3-(o-tolyloxy)-propylamine Hydrochloride
C1170741|(-)-N-methyl-gamma(2-methylphenoxy)benzenepropamine Hydrochloride
C1170741|ATOMOXETINE HCL
C1170741|atomoxetine HCl (medication)
C1170741|HCl, Atomoxetine
C1170741|Hydrochloride, Atomoxetine
C1170741|Atomoxetine Hydrochloride [Chemical/Ingredient]
C1170741|N-methyl-gamma-(2-methylphenoxy)benzenepropanamine hydrochloride
C1170741|Atomoxetine hydrochloride (substance)
C0771310|Nefazodone Hydrochloride
C0771310|antidepressants nefazodone hydrochloride
C0771310|nefazodone hydrochloride (medication)
C0771310|Nefazodone hydrochloride (substance)
C0771310|Nefazodone hydrochloride (product)
C0771310|Nefazadone HCl
C1881066|Homopipramol
C1881066|2-(4-(3-(5H-Dibenz(b,f)azepin-5-yl)propyl)-1,4-diazepin-1-yl)ethanol
C1881066|4-(3-(5H-Dibenz(b,f)azepin-5-yl)propyl)hexahydro-1H-1,4-diazepine-1-ethanol
C0071001|eptastigmine
C0071001|heptyl physostigmine
C0071001|physostigmine heptyl
C0071001|pyrrolo(2,3-b)indol-5-ol-1,2,3,3a,8,8a-hexahydro-1,3a,8-trimethyl heptylcarbamate ester
C0071001|heptastigmine
C0071001|heptylphysostigmine
C0071001|heptyl-physostigmine
C0724555|citalopram (as citalopram hydrobromide)
C0724555|Citalopram Hydrobromide
C0724555|(![PLUS-MINUS SIGN]!)-1-(3-dimethylaminopropyl)-1- (4-fluorophenyl)-1,3 dihydroisobenzofuran-5-carbonitrile, HBr
C0724555|(±)-1-(3-dimethylaminopropyl)-1- (4-fluorophenyl)-1,3 dihydroisobenzofuran-5-carbonitrile, HBr
C0724555|citalopram hydrobromide (medication)
C0724555|1-[3-(Dimethylamino)propyl]-1-(4-fluorophenyl)-1,3-dihydro-5-isobenzofurancarbonitrile Monohydrobromide
C0724555|Citalopram hydrobromide (substance)
C1880541|Eprobemide
C1881269|Irolapride
C0771019|Paroxetine hydrochloride
C0771019|paroxetine hydrochloride (medication)
C0771019|(-)-(3S,4R)-4-(p-Fluorophenyl)-3-((3,4-(methylenedioxy)phenoxy)methyl)piperidine Hydrochloride
C0771019|Paroxetine Hydrochloride [Chemical/Ingredient]
C0771019|Hydrochloride, Paroxetine
C0771019|Paroxetine hydrochloride (product)
C0771019|Paroxetine hydrochloride (substance)
C0282369|Trazodone Hydrochloride
C0282369|2-(3-(4-(3-Chlorophenyl)piperazin-1-y)propyl)-1,2,4-triazolo(4,3-a)pyridine-3(2H)-one Hydrochloride
C0282369|1,2,4-Triazolo(4,3-a)pyridin-3(2H)-one, 2-(3-(4-(3-chlorophenyl)-1-piperazinyl)propyl)-, Monohydrochloride
C0282369|trazodone hydrochloride (medication)
C0282369|antidepressants trazodone hydrochloride
C0282369|Trazodone Hydrochloride [Chemical/Ingredient]
C0282369|Trazodone hydrochloride (substance)
C0282369|Trazodone hydrochloride [dup] (substance)
C0208216|3-chloro-5-(3-(2-oxo-1,2,3,5,6,7,8,8a-octahydroimidazo(1,2-a)pyridine-3-spiro-4'-piperidino)propyl)-10,11-dihydro-5H-dibenz(b,f)azepine
C0208216|Mosapramine
C0208216|Spiro(imidazo(1,2-a)pyridine-3(2H),4'-piperidin)-2-one, 1'-(3-(3-chloro-10,11-dihydro-5H-dibenz(b,f)azepin-5-yl)propyl)hexahydro-, dihydrochloride
C0700473|Fluvoxamine maleate
C0700473|fluvoxamine maleate (medication)
C0700473|Fluvoxamine Maleate [Chemical/Ingredient]
C0700473|Fluvoxamine maleate (substance)
C0700473|Fluvoxamine Maleate, (E)-Isomer
C0700473|Fluvoxamine maleate [dup] (substance)
C1880815|Fluoxetine Hydrochloride, (R)-
C1880815|Fluoxetine Hydrochloride, R-
C1880815|Benzenepropanamine, N-methyl-gamma-(4-(trifluoromethyl)phenoxy)-, Hydrochloride (1:1), (gamma R)-
C0074710|2,6-Benzothiazolediamine, 4,5,6,7-tetrahydro-N6-propyl-, (S)-
C0074710|2-amino-4,5,6,7-tetrahydro-6-propylaminobenzothiazole
C0074710|pramipexole
C0074710|2-amino-6-propylaminotetrahydrobenzothiazole
C0074710|4,5,6,7-tetrahydro-N6-propyl-2,6-benzothiazole-diamine
C0074710|pramipexol
C0074710|Pramipexole (product)
C0074710|Pramipexole (substance)
C1882243|Oxitriptyline
C0127034|maroxepin
C0127034|maroxepine
C1882439|Prazitone
C1880799|Flubepride
C0125988|Cyclobenzaprine Hydrochloride
C0125988|Cloben
C0125988|3-(5H-Dibenzo(a,d)cyclohepten-5-ylidene)propyl(dimethyl)ammonium Chloride
C0125988|Cycloflex
C0125988|FR2100873
C0125988|Flexiban
C0125988|1-Propanamine, 3-(5H-dibenzo(a,d)cyclohepten-5-ylidene)-N,N-dimethyl-, Hydrochloride
C0125988|10,11delta-Amitriptyline Hydrochloride
C0125988|muscle relaxants skeletal cyclobenzaprine hydrochloride
C0125988|cyclobenzaprine hydrochloride (medication)
C0125988|Cyclobenzaprine hydrochloride (substance)
C0125988|Cyclobenzaprine hydrochloride (product)
C0063841|(4-chlorophenoxy)acetic acid 2-(1-methylethyl)hydrazide
C0063841|iproclozide
C0063841|p-(chlorophenoxy)acetic acid 2-isopropylhydrazide
C0606667|Pirolazamide
C0606667|hexahydro-alpha,alpha-diphenylpyrrolo-(1,2-alpha)pyrazine-2(1H)-butyramide
C1170746|Escitalopram Oxalate
C1170746|5-Isobenzofurancarbonitrile, 1-(3-(dimethylamino)propyl)-1-(4-fluorophenyl)-1,3-dihydro-,(1S)-, ethanedioate(1:1)
C1170746|escitalopram oxalate (medication)
C1170746|Escitalopram oxalate (substance)
C0060188|2-(4-chlorophenyl)-4-methyl-2,4-pentanediol
C0060188|fenpentadiol
C1881130|Imafen
C1882389|Pipofezine
C1881138|Imipraminoxide
C1880856|Ftormetazine
C0088224|1,3,4,9-tetrahydro-N,N,1-trimethylindeno(1,2-c)- pyran-1,ethylamine.HCl
C0088224|Pirandamine Hydrochloride
C1883593|Zafuleptine
C1883384|Trazolopride
C2347566|casopitant
C2349098|Valdipromide
C0608826|aceprometazine
C0608826|1-(10-(2-(dimethylamino)propyl)-10H-phenothiazin- 2-yl)ethanone
C0050721|2-(1-adamantylamino)ethyl(p-chlorophenoxy)acetate
C0050721|adafenoxate
C2347998|Afalanine
C2347998|Acetylphenylalanine
C0051694|amitriptyline N-oxide
C0051694|Amitriptylinoxide
C2346789|Ansoxetine
C2346868|Atibeprone
C2346892|Azaloxan Fumarate
C2346896|Azipramine
C2346971|Bazinaprine
C0053072|befuraline
C0053072|N-benzo(b)furan-2-ylcarbonyl-N'-benzylpiperazine.HCl
C0053611|1,2-Ethanediamine, N,N-dimethyl-N'-((3-phenyl-1H-indol-1-yl)methyl)-
C0053611|binedaline
C0053611|binodaline
C0054820|2,3-dihydro-4H-1,3-benzoxazin-2-one-3-acetamide
C0054820|2H-1,3-benzoxazine-3(4H)-acetamide, 2-oxo-
C0054820|4H-3-methylcarboxamide-1,3-benzoxazin-2-one
C0054820|caroxazone
C2348381|Efetozole
C2348443|Enefexine
C2348450|Enprazepine
C0060170|2-(N-butyl-o-chlorobenzimidoyl)-4-chlorophenyl
C0060170|fengabine
C0060305|fezolamine
C0956920|Fezolamine Fumarate
C0537150|3alpha-hydroxy-3beta-methyl-5alpha-pregnan-20-one
C0537150|ganaxolone
C2347511|Piberaline
C0072207|propizepin
C0072207|propizepine
C0072207|pyridobenzodiazepine
C0076671|9-ethyl-4-fluoro-1-methyl-7,8,9,10-tetrahydrothieno(3,2e)pyrido(4,3b)indole lactate
C0076671|tiflucarbine
C2348815|Trazium Esilate
C0132764|7-(1,2-dimethylheptyl)-2,2-dimethyl-4-(4-pyridinyl)-2H-1-benzopyran-5-ol
C0132764|nonabine
C2347355|Nitrafudam Hydrochloride
C2348183|Seproxetine Hydrochloride
C2348647|Talopram Hydrochloride
C0076823|atomoxetine
C0076823|Tomoxetine
C0076823|Atomoxetine (product)
C0076823|Atomoxetine (substance)
C0051607|10,11-dihydrodibenzo(a,d)cyclohept-5-enyl-7-aminoheptanoic acid
C0051607|7-((10,11-dihydro-5H-dibenzo(a,d)cyclohepten-5-yl)amino)heptanoic acid
C0051607|amineptin
C0051607|amineptine
C2168874|pyritinol + cyproheptadine + vitamins (medication)
C2168874|pyritinol + cyproheptadine + vitamins
C0071125|pirandamine
C0600985|1-naphthalenamine, 8-chloro-1,2,3,4-tetrahydro-5-methoxy-N,N-dimethyl-
C0600985|N,N-dimethyl-5-methoxy-8-chloro-1,2,3,4-tetrahydro-1-naphthylamine
C0600985|lometraline
C0888036|Lometraline Hydrochloride
C0113211|N-desmethylsertraline
C0113211|N-demethylsertraline
C0113211|desmethylsertraline
C0113211|Desmethylsertraline (substance)
C3650305|antidepressants fluoxetine
C3650305|antidepressants fluoxetine (medication)
C3650304|antidepressants fluvoxamine
C3650304|antidepressants fluvoxamine (medication)
C3650297|antidepressants paroxetine (medication)
C3650297|antidepressants paroxetine
C3650299|antidepressants nefazodone
C3650299|antidepressants nefazodone (medication)
C0068987|desmethylfluoxetine
C0068987|norfluoxetin
C0068987|norfluoxetine
C0068987|Norfluoxetine (substance)
C0719199|Celexa
C0719199|citalopram hydrobromide (Celexa)
C0162373|Prozac
C0376414|Paxil
C0709644|Sertraline 50 MG Oral Tablet [Zoloft]
C0709644|Zoloft 50 MG Oral Tablet
C0709644|Zoloft 50mg Tablet
C0709644|Zoloft, 50 mg oral tablet
C0709644|Zoloft (as sertraline hydrochloride) 50 MG Oral Tablet
C0709644|SERTRALINE HYDROCHLORIDE 50 mg ORAL TABLET, FILM COATED [ZOLOFT]
C0709644|Sertraline Hydrochloride 50 MG Oral Tablet [ZOLOFT]
C0709632|Sertraline 100 MG Oral Tablet [Zoloft]
C0709632|Zoloft 100mg Tablet
C0709632|Zoloft, 100 mg oral tablet
C0709632|Zoloft (as sertraline hydrochloride) 100 MG Oral Tablet
C0709632|SERTRALINE HYDROCHLORIDE 100 mg ORAL TABLET, FILM COATED [ZOLOFT]
C0709632|Sertraline Hydrochloride 100 MG Oral Tablet [ZOLOFT]
C0709632|Zoloft 100 MG Oral Tablet
C0284660|Zoloft
C0284660|Altruline
C0284660|Parke Davis Brand of Sertraline Hydrochloride
C0284660|Lustral
C0284660|Roerig Brand of Sertraline Hydrochloride
C0284660|Pfizer Brand of Sertraline Hydrochloride
C0060926|1-(aminomethyl)cyclohexaneacetic acid
C0060926|gabapentin
C0060926|gabapentin (medication)
C0060926|gabapentin [Chemical/Ingredient]
C0060926|Convalis
C0060926|Gabapentin (product)
C0060926|Gabapentin (substance)
C0678176|Neurontin
C0657912|pregabalin
C0657912|3-(Aminomethyl)-5-methyl-hexanoic Acid
C0657912|3-Isobutyl GABA
C0657912|pregabalin (medication)
C0657912|(S+)-3-isobutyl GABA
C0657912|(R-)-3-isobutyl GABA
C0657912|3-(aminomethyl)-5-methylhexanoic acid
C0657912|(S)-3-(aminomethyl)-5-methylhexanoic acid
C0657912|GABA, 3-isobutyl
C0657912|3 isobutyl GABA
C0657912|Pregabalin [Chemical/Ingredient]
C0657912|Pregabalin (product)
C0657912|Pregabalin (substance)
C2740401|pregabalin 20 MG/ML Oral Solution
C2740401|Pregabalin 20mg/mL oral solution
C2740401|Pregabalin 20mg/mL oral solution (product)
C2740401|Pregabalin Soln 20 MG/ML
C2740401|Pregabalin 20mg Oral solution
C2740401|PREGABALIN 20MG/ML SOLN,ORAL
C2740401|PREGABALIN 20MG/ML ORAL SOLN
C2740401|PREGABALIN 20MG/ML SOLN,ORAL [VA Product]
C1532848|pregabalin 200 MG Oral Capsule
C1532848|Pregabalin Cap 200 MG
C1532848|PREGABALIN 200MG CAP,ORAL
C1532848|PREGABALIN 200MG ORAL CAP
C1532848|PREGABALIN 200MG CAP,ORAL [VA Product]
C1532848|Pregabalin 200mg Oral capsule
C1532848|Pregabalin 200mg capsule (product)
C1532848|Pregabalin 200mg capsule
C1532851|pregabalin 50 MG Oral Capsule
C1532851|Pregabalin Cap 50 MG
C1532851|PREGABALIN 50MG CAP,ORAL
C1532851|PREGABALIN 50MG ORAL CAP
C1532851|PREGABALIN 50MG CAP,UD
C1532851|PREGABALIN 50MG CAP UD
C1532851|PREGABALIN 50MG CAP,ORAL [VA Product]
C1532851|PREGABALIN 50MG CAP,UD [VA Product]
C1532851|Pregabalin 50mg Oral capsule
C1532851|Pregabalin 50mg capsule (product)
C1532851|Pregabalin 50mg capsule
C1532852|pregabalin 75 MG Oral Capsule
C1532852|Pregabalin Cap 75 MG
C1532852|PREGABALIN 75MG CAP,ORAL
C1532852|PREGABALIN 75MG CAP,UD
C1532852|PREGABALIN 75MG ORAL CAP
C1532852|PREGABALIN 75MG CAP UD
C1532852|PREGABALIN 75MG CAP,ORAL [VA Product]
C1532852|PREGABALIN 75MG CAP,UD [VA Product]
C1532852|Pregabalin 75mg Oral capsule
C1532852|Pregabalin 75mg capsule (product)
C1532852|Pregabalin 75mg capsule
C1532849|pregabalin 25 MG Oral Capsule
C1532849|Pregabalin Cap 25 MG
C1532849|PREGABALIN 25MG CAP,ORAL
C1532849|PREGABALIN 25MG ORAL CAP
C1532849|PREGABALIN 25MG CAP,ORAL [VA Product]
C1532849|Pregabalin 25mg Oral capsule
C1532849|Pregabalin 25mg capsule (product)
C1532849|Pregabalin 25mg capsule
C1532847|pregabalin 150 MG Oral Capsule
C1532847|Pregabalin Cap 150 MG
C1532847|PREGABALIN 150MG CAP,ORAL
C1532847|PREGABALIN 150MG CAP UD
C1532847|PREGABALIN 150MG ORAL CAP
C1532847|PREGABALIN 150MG CAP,UD
C1532847|PREGABALIN 150MG CAP,ORAL [VA Product]
C1532847|PREGABALIN 150MG CAP,UD [VA Product]
C1532847|Pregabalin 150mg Oral capsule
C1532847|Pregabalin 150mg capsule (product)
C1532847|Pregabalin 150mg capsule
C0388352|CI 1008
C0388352|CI1008
C0388352|1008, CI
C0388352|CI-1008
C1972026|Pregabalin &#x7C; Bld-Ser-Plas
C3170841|Pregabalin &#x7C; Urine
C1570232|Lyrica
C1532846|pregabalin 100 MG Oral Capsule
C1532846|Pregabalin Cap 100 MG
C1532846|PREGABALIN 100MG CAP,ORAL
C1532846|PREGABALIN 100MG CAP,UD
C1532846|PREGABALIN 100MG ORAL CAP
C1532846|PREGABALIN 100MG CAP UD
C1532846|PREGABALIN 100MG CAP,UD [VA Product]
C1532846|PREGABALIN 100MG CAP,ORAL [VA Product]
C1532846|Pregabalin 100mg Oral capsule
C1532846|Pregabalin 100mg capsule (product)
C1532846|Pregabalin 100mg capsule
C1532850|pregabalin 300 MG Oral Capsule
C1532850|Pregabalin Cap 300 MG
C1532850|PREGABALIN 300MG CAP,ORAL
C1532850|PREGABALIN 300MG ORAL CAP
C1532850|PREGABALIN 300MG CAP,ORAL [VA Product]
C1532850|Pregabalin 300mg Oral capsule
C1532850|Pregabalin 300mg capsule (product)
C1532850|Pregabalin 300mg capsule
C1613977|pregabalin 225 MG Oral Capsule
C1613977|Pregabalin Cap 225 MG
C1613977|Pregabalin 225mg capsule (product)
C1613977|Pregabalin 225mg capsule
C1613977|PREGABALIN 225MG CAP,ORAL
C1613977|PREGABALIN 225MG ORAL CAP
C1613977|PREGABALIN 225MG CAP,ORAL [VA Product]
C1613977|Pregabalin 225mg Oral capsule
C1955823|PD 144723
