C1255280|25-Oh D Vitamin Test
C1255280|Vit D 25-OH
C1255280|Vitamin D 25-OH
C1255280|Vitamin D 25-OH
