C0085178|Needlestick Injuries
C0582072|Sharps Injuries
C0561474|Needle stick injury of nose
C0561474|Needle stick injury of nose (disorder)
C0085178|Injuries, Needle-Stick
C0085178|Injury, Needle-Stick
C0085178|Injury, Needlestick
C0085178|Needle Stick Injuries
C0085178|Needle Sticks
C0085178|Needle-Stick
C0085178|Needle-Stick Injury
C0085178|Needlestick
C0085178|Needlestick Injuries
C0085178|Needlestick Injury
C0085178|NEEDLESTICK INJ
C0085178|INJ NEEDLESTICK
C0085178|Needlesticks
C0085178|Needle-Stick Injuries
C0085178|Needle-Sticks
C0085178|Injuries, Needlestick
C0085178|Needlestick Injuries [Disease/Finding]
C0085178|Injury;needle stick
C0085178|Needle stick
C0085178|Needle prick injury
C0085178|Needle stick injury
C0085178|Needle stick injury (disorder)
C2116782|puncture by needle
C2116782|puncture by needle (physical finding)
C0582070|Needle stick injury with clean needle
C0582070|Needle stick injury with clean needle (disorder)
C0582071|Needle stick injury with contaminated needle
C0582071|Needle stick injury with dirty needle
C0582071|Needle stick injury with contaminated needle (disorder)
C0561467|Needle stick injury of head and neck
C0561467|Needle stick injury of head and neck (disorder)
C0561500|Needle stick injury of lower limb
C0561500|Needle stick injury of lower limb (disorder)
C0561479|Needle stick injury of upper limb
C0561479|Needle stick injury of upper limb (disorder)
C0561491|Needle stick injury of trunk
C0561491|Needle stick injury of trunk (disorder)
C0582072|Sharps injury
C0582072|Sharps injury (disorder)
C0582072|Injuries, Sharps
C0582072|Injury, Sharps
C0582072|Sharps Injuries
