C0003962|Ascites
C0741240|ASCITES FLUID INFECTION
C0741242|ASCITES NEW ONSET
C0741245|ASCITES UNKNOWN ORIGIN
C0003964|Peritoneal Fluid (body substance)
C0401037|Hepatic ascites
C0003962|Ascites
C0003962|[D]Ascites (context-dependent category)
C0003962|[D]Ascites NOS (context-dependent category)
C0003962|abdominal dropsy
C0003962|hydrops abdominis
C0003962|peritoneal dropsy
C0003962|peritoneal exudate
C0003962|hydroperitonia
C0003962|abdominal ascites
C0003962|ascites (physical finding)
C0003962|ascites (diagnosis)
C0003962|abdomen ascites
C0003962|ascites was discovered
C0003962|Ascites NOS
C0003962|Ascites [Disease/Finding]
C0003962|[D]Ascites (situation)
C0003962|[D]Ascites NOS (situation)
C0003962|Ascites (disorder)
C0003962|[D]Ascites NOS
C0003962|[D]Ascites
C0003962|Hydroperitoneum
C0003962|INCREASING ABDOMINAL DISTENTION OR ASCITES
C0003962|abdominis; hydrops
C0003962|hydrops; abdominis
C0003962|Ascites, NOS
C2227708|abdominal x-ray, AP view: ascites (procedure)
C2227708|abdominal x-ray, AP view: ascites
C0220656|malignant ascites
C0220656|malignant ascites (diagnosis)
C0220656|Ascites, Malignant
C0220656|Malignant ascites (disorder)
C0220656|Malignant ascites, NOS
C0220656|Malignant peritoneal effusion
C0220656|ascites; malignant
C0220656|malignant; ascites
C1955521|Other ascites
C1955521|Ascites NEC
C2142846|pseudochylous ascites
C2142846|pseudochylous ascites (diagnosis)
C0426682|Fluid wave
C0426682|abdominal fluid wave
C0426682|ascites fluid wave
C0426682|abdominal fluid wave (physical finding)
C0426682|Finding of fluid thrill of abdomen (finding)
C0426682|Finding of fluid thrill of abdomen
C0426682|Fluid thrill
C0426682|Fluid thrill in abdomen
C0426682|Observation of fluid thrill of abdomen
C0426682|Fluid thrill in abdomen (finding)
C0277979|Shifting abdominal dullness finding
C0277979|ascites shifting dullness
C0277979|abdominal shifting dullness
C0277979|shifting dullness of abdomen
C0277979|abdominal shifting dullness (physical finding)
C0277979|ascites with shifting dullness was discovered
C0277979|Shifting dullness (finding)
C0277979|Shifting dullness
C0277979|Shifting abdominal dullness
C0277979|Shifting abdominal dullness (observable entity)
C0277979|Shifting abdominal dullness finding (finding)
C0426679|abdominal puddle sign
C0426679|abdominal puddle sign (physical finding)
C0426679|ascites puddle sign
C0426679|Puddle sign
C0426679|Puddle sign (finding)
C0741244|ascites tense
C0741244|tense abdomen (physical finding)
C0741244|tense abdomen
C0741244|tense ascites was discovered
C0741244|Tense ascites
C0741244|Tense ascites (disorder)
C2022430|echocardiography: ascites (procedure)
C2022430|echocardiography: ascites
C2321829|sample template ascites (diagnosis)
C2321829|sample template ascites
C3532188|Refractory ascites
C3532188|Refractory ascites (disorder)
C0269720|disproportion at birth due to fetal ascites (diagnosis)
C0269720|disproportion at birth due to fetal ascites
C0269720|disproportion (at birth) due to fetal ascites
C0269720|Foetal ascites causing disproportion
C0269720|Fetal ascites causing disproportion
C0269720|Fetal ascites causing disproportion (disorder)
C0269720|disproportion; fetal ascites
C0269720|fetal; ascites, disproportion
C0585187|Infected ascites
C0585187|Infected ascites (disorder)
C0267773|Biliary ascites
C0267773|Bile ascites
C0267773|Bile ascites (disorder)
C0267774|Urine ascites
C0267774|Urine ascites (disorder)
C0267774|Uroabdomen
C0019086|Haemorrhagic ascites
C0019086|Hemorrhagic peritoneal effusion
C0019086|Hemorrhagic ascites
C0019086|Hemorrhagic ascites (disorder)
C0031144|Chronic peritoneal effusion (disorder)
C0031144|chronic peritoneal effusion
C0031144|chronic peritoneal effusion (diagnosis)
C0031144|Peritoneal effusion
C0031144|Peritoneal effusion (chronic)
C0008732|Chylous ascites
C0008732|ASCITES, CHYLOUS
C0008732|chyloperitoneum
C0008732|chylous ascites (diagnosis)
C0008732|Chylous Ascites [Disease/Finding]
C0008732|Ascites chylous
C0008732|Chylous ascites (disorder)
C0008732|ascites; chylous
C0008732|chylous; ascites
C0341525|Cardiac ascites
C0341525|Cardiac ascites (disorder)
C0267772|Pancreatic ascites
C0267772|Pancreatic ascites (disorder)
C0025184|Meig Syndrome
C0025184|Meig's Syndrome
C0025184|Meigs' syndrome
C0025184|Meigs Syndrome
C0025184|Meig's syndrome (diagnosis)
C0025184|Meigs Syndrome [Disease/Finding]
C0025184|Demons-Meigs syndrome
C0025184|Ovarian-ascites-pleural effusion syndrome
C0025184|Meigs-Cass syndrome
C0025184|Meigs' syndrome (disorder)
C0267776|Dialysis-associated ascites
C0267776|Dialysis-associated ascites (disorder)
C0401038|Hypoalbuminaemic ascites
C0401038|Metabolic ascites
C0401038|Hypoalbuminemic ascites
C0401038|Metabolic ascites (disorder)
C0401037|Hepatic ascites
C0401037|Hepatic ascites (disorder)
C3670559|Fibrinous peritoneal effusion
C3670559|Fibrinous ascites
C3670559|Fibrinous ascites (disorder)
C3670560|Modified transudative peritoneal effusion
C3670560|Modified transudative ascites (disorder)
C3670560|Modified transudative ascites
C3670560|Modified transudate ascites
C0519092|Transudate ascites
C0519092|Transudative peritoneal effusion
C0519092|Transudative ascites (disorder)
C0519092|Transudative ascites
C1285291|Fetal ascites
C1285291|Fetal ascities
C1285291|Foetal ascites
C1285291|fetus; ascites
C1285291|Fetal ascites (disorder)
C1285291|Fetal ascities (disorder)
C4038874|Ascites due to alcoholic cirrhosis (disorder)
C4038874|Ascites due to alcoholic cirrhosis
C4038944|Ascites due to alcoholic hepatitis
C4038944|Ascites due to alcoholic hepatitis (disorder)
C0275919|Tuberculous ascites
C0275919|Tuberculous ascites (disorder)
C0275919|ascites; tuberculous
C3665480|[D]Fluid in peritoneal cavity (context-dependent category)
C3665480|fluid in peritoneal cavity
C3665480|[D]Fluid in peritoneal cavity (situation)
C3665480|[D]Fluid in peritoneal cavity
C3665480|Fluid in peritoneal cavity (finding)
C1385680|effusion; abdomen
C1385680|abdomen; effusion
C1390873|abdomen; upset, fluid
C1390873|upset; abdomen, fluid
C1390876|distension; abdomen, fluid
C1390876|abdomen; distension, fluid
C1390885|effusion; peritoneal cavity
C1390885|peritoneal cavity; effusion
C0003964|Ascitic Fluid
C0003964|Ascitic Fluids
C0003964|Effusion, Peritoneal
C0003964|Effusions, Peritoneal
C0003964|Fluid, Ascitic
C0003964|Fluid, Peritoneal
C0003964|Fluids, Ascitic
C0003964|Fluids, Peritoneal
C0003964|Peritoneal Effusions
C0003964|Peritoneal Fluids
C0003964|peritoneal fluid
C0003964|Peritoneal Fluid (body substance)
C0003964|Peritoneal fluid (substance)
C0003964|Peritoneal effusion
C0003964|Fluid, Ascites
C0003964|effusion; peritoneal
C0003964|peritoneal; effusion
C0003964|Ascitic fluid (substance)
C0437001|On examination - ascites
C0437001|O/E - ascites
C0437001|O/E - ascites NOS (finding)
C0437001|On examination - ascites NOS
C0437001|O/E - ascites NOS
C0437001|On examination - ascites NOS (disorder)
C0437001|O/E - ascites (finding)
C0437001|On examination - ascites (context-dependent category)
C0437001|On examination - ascites NOS (context-dependent category)
C0437001|On examination - ascites (disorder)
C4038684|Hepatic ascites co-occurrent with chronic active hepatitis due to toxic liver disease
C4038684|Hepatic ascites co-occurrent with chronic active hepatitis due to toxic liver disease (disorder)
C4040413|Hepatic ascites due to chronic alcoholic hepatitis (disorder)
C4040413|Hepatic ascites due to chronic alcoholic hepatitis
