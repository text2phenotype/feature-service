C0024808|Smokes weed
C0024808|Weed smoker
C0024808|Marijuana smoker
C0024808|Smokes marijuana
C0024808|Marihuana
C0024809|Marijuana Abuse
C0678449|Cannabis substance
C0700268|Cannabis sativa plant
C0936079|Cannabis
C0936079|Cannabis smoker
C0936079|Smokes cannabis
C1547291|Marijuana Recreational Drug Use Code
C0024808|Marihuana
C0024808|MARIJUANA
C0024808|Cannabis
C0024808|Marijuanas
C0024808|Marihuanas
C0024808|MARIJUANA [VA Product]
C0024809|Abuse, Marihuana
C0024809|Abuse, Marijuana
C0024809|Marijuana Abuse
C0024809|marijuana
C0024809|Marihuana Abuse
C0024809|Marijuana Abuse [Disease/Finding]
C0024809|Abuse;drug(s);marijuana
C0024809|Cannabis
C0024809|Hash
C0024809|Weed
C0024809|Pot
C0024809|abuse; marihuana
C0024809|marihuana; abuse
C0018614|Abuse, Hashish
C0018614|hashish; abuse
C0018614|abuse; hashish
C0018614|Hashish Abuse
C0017089|Ganjas
C0017089|Ganja
C0018210|Gramineae
C0018210|Poaceae
C0018210|Grass
C0018210|Grasses
C0018210|Family Gramineae
C0018210|Family Poaceae (organism)
C0018210|Family Poaceae
C0018210|Family poaceae - gramineae
C0018210|Grass (organism)
C0018210|Family poaceae - gramineae (organism)
C0018210|grass family
C0006863|Cannabidiol
C0006863|1,3-Benzenediol, 2-(3-methyl-6-(1-methylethenyl)-2-cyclohexen-1-yl)-5-pentyl-, (1R-trans)-
C0006863|Cannabidiol [Chemical/Ingredient]
C0006863|CBD
C0006863|Cannabidiol (substance)
C0006865|Cannabinol
C0006865|6H-Dibenzo(b,d)pyran-1-ol, 6,6,9-trimethyl-3-pentyl-
C0006865|3-Amyl-1-hydroxy-6,6,9-trimethyl-6H-dibenzo(b,d)pyran
C0006865|Cannabinol [Chemical/Ingredient]
C0006865|6,6,9-Trimethyl-3-pentyl-6H-dibenzo(b,d)pyran-1-ol
C0006865|CBN
C0006865|Cannabinol (substance)
C0556618|Cannabis grass - non-pharmaceutical
C0556618|Marijuana grass
C0556618|Marihuana grass
C0556618|Cannabis grass - non-pharmaceutical (substance)
C0700258|Marijuana leaf
C0700258|Cannabis leaves - non-pharmaceutical
C0700258|Marihuana leaf
C0700258|Cannabis leaves - non-pharmaceutical (substance)
C0556617|Cannabis oil - non-pharmaceutical
C0556617|Marijuana oil
C0556617|Marihuana oil
C0556617|Cannabis oil - non-pharmaceutical (substance)
C0018613|hashish
C0018613|Hashishs
C0018613|Cannabis resin - non-pharmaceutical
C0018613|Marijuana resin
C0018613|Marihuana resin
C0018613|Cannabis resin - non-pharmaceutical (substance)
C0005337|Bhangs
C0005337|Bhang
C0700268|marijuana
C0700268|Cannabis sativa
C0700268|Cannabis sativa plant
C0700268|sativas, Cannabis
C0700268|Cannabis sativas
C0700268|sativa, Cannabis
C0700268|Cannabis sativa L.
C0700268|Cannabis
C0700268|CANNABIS SATIVA WHOLE
C0700268|Marihuana
C0700268|Indian hemp
C0700268|Cannabis sativa (organism)
C0162335|Hemp
C0162335|Hemps
C0162335|Hemp (physical object)
C0949248|indica, Cannabis
C0949248|indicas, Cannabis
C0949248|Cannabis indicas
C0949248|Cannabis indica
C0936079|Cannabis
C0936079|Plant, Hemp
C0936079|Hemp Plants
C0936079|Plants, Hemp
C0936079|Cannabi
C0936079|Cannabis L., 1753
C0936079|Hemp Plant
C0936079|Cannabis (organism)
C0936079|Cannabis, NOS
C0936079|Hemp (Cannabis)
