C0199967|Transfusion of coagulation factors
C0199967|Blood Transfusion
C0852255|Blood and blood product treatment
C0481253|Contaminated substance transfused or infused (finding)
C0481253|Contaminated substance transfused or infused
C0730400|Solid organ transplant
C0857825|Infection in solid organ transplant recipients
C0199967|Clotting factor transfusion
C0199967|Coag factor transfusion
C0199967|Transfusion of coagulation factors
C0199967|Transfusion of coagulation factor
C0199967|Transfusion of coagulation factors (procedure)
C0199968|Antihaemophilic factor transfusion (procedure)
C0199968|Antihemophilic factor transfusion
C0199968|Transfusion of antihemophilic factor
C0199968|Transfusion of antihaemophilic factor
C0199968|Antihaemophilic factor transfusion
C0199968|Transfusion of antihemophilic factor (procedure)
C0199968|Antihemophilic factor transfusion (procedure)
C2242940|plasma fractions, human (treatment)
C2242940|plasma fractions, human
C3161607|plasma fractions, human factor xiii concentrate (human)
C3161607|plasma fractions, human factor xiii concentrate (human) (treatment)
C2064859|plasma fractions, human factor VIII (AHF, AHG)
C2064859|plasma fractions, human factor VIII (AHF, AHG) (treatment)
C2064857|plasma fractions, human albumin, normal serum (treatment)
C2064857|plasma fractions, human albumin, normal serum
C2064858|plasma fractions, factor IX complex (human)
C2064858|human factor IX complex (human)
C2064858|human factor IX complex (human) (treatment)
C2194217|factor VIIa transfusion (treatment)
C2194217|factor VIIa
C2194217|factor VIIa (treatment)
C2069055|plasma fractions, human albumin + globulin (treatment)
C2069055|plasma fractions, human albumin + globulin
C2069056|plasma fractions, antithrombin III (human) (treatment)
C2069056|plasma fractions, antithrombin III (human)
C4064322|plasma fractions, coagulation factor X (human) (treatment)
C4064322|plasma fractions, coagulation factor X (human)
C4064322|plasma fractions, human factor x
C1293889|Coagulation factor IX product administration by intravascular infusion
C1293889|Transfusion of factor IX (procedure)
C1293889|Transfusion of factor IX
C1293888|Coagulation factor VII product administration by intravascular infusion
C1293888|Transfusion of factor VII (procedure)
C1293888|Transfusion of factor VII
C1960763|Transfusion antithrombin III factor (procedure)
C1960763|Transfusion antithrombin III factor
C0854629|Allogenic bone marrow transplantation therapy
C0854630|Autologous bone marrow transplantation therapy
C0005842|Autotransfusion
C0005842|Autotransfusions
C0005842|Blood Transfusion, Autologous
C0005842|Autotransfusion Procedure
C0005842|TRANSFUSION AUTOL BLOOD
C0005842|BLOOD TRANSFUSIONS AUTOL
C0005842|AUTOL BLOOD TRANSFUSIONS
C0005842|TRANSFUSIONS AUTOL BLOOD
C0005842|BLOOD TRANSFUSION AUTOL
C0005842|AUTOL BLOOD TRANSFUSION
C0005842|autotransfusion (treatment)
C0005842|Blood--Transfusion, Autologous
C0005842|Autologous blood transfusion
C0005842|Blood Transfusions, Autologous
C0005842|Autologous Blood Transfusions
C0005842|Transfusion, Autologous Blood
C0005842|Transfusions, Autologous Blood
C0005842|Abt - autologous blood transfusion
C0005842|Autotransfusion (procedure)
C0005842|Autotransfusion, NOS
C0005842|Intravenous autotransfusion each treatment
C0005842|IV autotransfusion ea.Tx
C0854631|Cord blood transplant therapy
C0015236|Exchange Transfusion, Whole Blood
C0015236|blood exchange transfusion
C0015236|Exchange blood transfusion
C0015236|EXCHANGE TRANSFUSION
C0015236|exchange transfusion (treatment)
C0015236|Exchange transfusion of blood
C0015236|Exchange blood transfusion NOS
C0015236|Exchange blood transfusion NOS (procedure)
C0015236|Exchange transfusion, blood
C0015236|Transfusion replacement, total
C0015236|Exsanguination transfusion
C0015236|EBT - Exchange blood transfusion
C0015236|Exchange transfusion (procedure)
C0015236|Transfusion, exsanguination
C0854634|Mismatched donor bone marrow transplantation therapy
C0371803|Exchange transfusion, blood; newborn
C0371803|Neonatal exchange blood transfusion
C0371803|exchange transfusion of newborn (treatment)
C0371803|exchange transfusion of newborn
C0371803|Neonatal exchange transfusion
C0371803|BL EXCHANGE/TRANSFUSE NB
C0371803|EXCHNG TRANSFUSION BLOOD NEWBORN
C0371803|Exchange blood transfusion, newborn
C0371803|Exchange blood transfusion (neonatal)
C0371803|Neonatal exchange transfusion (procedure)
C0199962|packed red blood cell transfusion
C0199962|Transfusion of packed red blood cells
C0199962|Red Blood Cell Transfusion
C0199962|Transfusion of PRBC
C0199962|Intravenous blood transfusion of packed cells
C0199962|Intravenous blood transfusion of packed cells (procedure)
C0199962|Transfusion of packed red blood cells (procedure)
C0199962|PRBC Transfusion
C0199964|Plasma expander transfusion
C0199964|Blood expander transfus
C0199964|Blood expander transfusion
C0199964|Transfusion of blood expander
C0199964|Plasma expander transfusion (procedure)
C0199964|Transfusion of blood expander (procedure)
C0199964|Transfusion of plasma expander
C0199964|Transfusion of blood expander, NOS
C0199964|Transfusion of plasma expander, NOS
C0032134|Plasmaphereses
C0032134|Plasmapheresis
C0032134|Therapeu plasmapheresis
C0032134|Plasmaphoresis
C0032134|Plasma Exchange
C0032134|Plasmapheresis (procedure)
C0032134|therapeutic plasmapheresis
C0032134|Therapeutic Plasma Exchange
C0086818|Platelet Transfusion
C0086818|Platelet Transfusions
C0086818|Transfusion, Platelet
C0086818|Transfusions, Platelet
C0086818|Blood Platelet Transfusions
C0086818|Platelet Transfusion, Blood
C0086818|Platelet Transfusions, Blood
C0086818|Transfusion, Blood Platelet
C0086818|Transfusions, Blood Platelet
C0086818|transfusion of platelets (treatment)
C0086818|transfusion of platelets
C0086818|Platelet transfusion (procedure)
C0086818|Blood platelets--Transfusion
C0086818|Blood Platelet Transfusion
C0086818|Transfusion of thrombocytes
C0086818|Intravenous blood transfusion of platelets
C0086818|Intravenous blood transfusion of platelets (procedure)
C0854635|Unrelated donor bone marrow transplantation therapy
C0677960|T lymphocyte depletion therapy
C0677960|T-cell depletion
C0677960|T-Lymphocyte Depletion Therapy
C0677960|T-Cell Depletion Therapy
C0919689|Donor leukocyte infusion
C0194015|Bone marrow harvest
C0194015|aspiration of bone marrow from donor for transplant
C0194015|aspiration of bone marrow from donor for transplant (treatment)
C0194015|bone marrow collection for transplant (treatment)
C0194015|bone marrow collection for transplant
C0194015|Donor marrow aspiration
C0194015|Bone marrow harvesting
C0194015|Harvest of bone marrow
C0194015|Aspiration of bone marrow from donor for transplant (procedure)
C0023416|Leukaphereses
C0023416|Leukapheresis
C0023416|Leukocytaphereses
C0023416|Leukocytophereses
C0023416|Leukophereses
C0023416|therapeutic leukopheresis (treatment)
C0023416|therapeutic leukopheresis
C0023416|Therapeutc leukopheresis
C0023416|Leukopheresis
C0023416|Leukocytapheresis
C0023416|Leukocytopheresis
C0023416|Leucapheresis
C0023416|Leukopheresis (procedure)
C0023416|Therapeutic leukocytapheresis
C0079186|Cytaphereses
C0079186|Cytapheresis
C0411265|Blood stem cell harvest
C0411265|Stem cell harvesting
C0411265|Harvest of stem cells
C0411265|Harvest of stem cells (procedure)
C0411265|Harvesting of stem cells (procedure)
C0411265|Harvesting of stem cells
C0948144|Peripheral blood stem cell apheresis
C0948145|Erythrocytapheresis
C0948145|Erythrocytapheresis (procedure)
C0949035|Low density lipoprotein apheresis (procedure)
C0949035|Low density lipoprotein apheresis
C0949035|LDL apheresis
C0032202|Blood Plateletphereses
C0032202|Plateletphereses
C0032202|Plateletphereses, Blood
C0032202|Plateletpheresis
C0032202|Plateletpheresis, Blood
C0032202|Thrombocytaphereses
C0032202|Thrombocytophereses
C0032202|Therapeutic plateletpheresis
C0032202|cellular apheresis for platelets (treatment)
C0032202|therapeutic plateletpheresis (treatment)
C0032202|cellular apheresis for platelets
C0032202|apheresis for platelets
C0032202|Therapeu plateltpheresis
C0032202|THERAPEUTIC APHERESIS PLATELETS
C0032202|Mechanical separation of platelet cells from blood
C0032202|Therapeutic apheresis for platelets
C0032202|Therapeutic apheresis; for platelets
C0032202|Blood Plateletpheresis
C0032202|Thrombocytapheresis
C0032202|Thrombocytopheresis
C0032202|Platelet apheresis
C0032202|Plateletpheresis (procedure)
C0032202|APHERESIS PLATELETS
C0948460|Vascular catheter specimen collection
C0524864|Hematopoietic Stem Cell Mobilization
C0524864|Mobilization, Stem Cell
C0524864|Haematopoietic stem cell mobilisation
C0524864|Hematopoietic stem cell mobilisation
C0524864|Stem cell mobilisation
C0524864|Stem cell mobilization
C0005791|Aphereses
C0005791|Blood Component Removal
C0005791|Blood Component Removals
C0005791|Component Removal, Blood
C0005791|Component Removals, Blood
C0005791|Phereses
C0005791|Removal, Blood Component
C0005791|Removals, Blood Component
C0005791|Apheresis (procedure)
C0005791|Apheresis
C0005791|Apheresis.therapeutic
C0005791|Therapeutic apheresis (procedure)
C0005791|Therapeutic apheresis
C0005791|Pheresis
C0005791|Collection, Apheresis/Leukapheresis
C0005791|Apheresis NOS
C0005791|Hemapheresis
C0005791|Apheresis procedure
C0005791|Apheresis - action (qualifier value)
C0005791|Apheresis - action
C0005791|Therapeutic apheresis, NOS
C0206373|Photopheresis
C0206373|Extracorporeal Photochemotherapies
C0206373|Photochemotherapies, Extracorporeal
C0206373|Photopheresis, Extracorporeal
C0206373|extracorporeal photophoresis
C0206373|EXTRACORPOREAL PHOTOCHEMOTHER
C0206373|PHOTOCHEMOTHER EXTRACORPOREAL
C0206373|Extracorporeal Photopheresis
C0206373|photopheresis (treatment)
C0206373|Photophoresis
C0206373|Therapeutc photopheresis
C0206373|PHOTOPHERESIS EXTRACORPOREAL
C0206373|Extracorporeal Photochemotherapy
C0206373|Photochemotherapy, Extracorporeal
C0206373|Extracorporeal photopheresis (procedure)
C0206373|Therapeutic photopheresis
C1879316|Transfusion
C1879316|Transfusion (procedure)
C1879316|transfusions
C1879316|transfusions (treatment)
C1879316|Transfusion, NOS
C0852255|Blood and blood product treatment
C4049189|Immunoadsorption therapy
C0481253|Contaminated transfusion
C0481253|Contaminated substance transfused or infused (event)
C0481253|Contaminated substance transfused or infused NOS (event)
C0481253|Contaminated substance transfused or infused
C0481253|Contaminated substance transfused or infused NOS
C0481253|Contaminated substance transfused or infused (finding)
C0481253|Contaminated substance transfused or infused NOS (finding)
C1261338|Contaminated medical or biological substance, transfused or infused
C1261338|Injury due to contaminated medical or biological substance, transfused or infused
C1261338|Contaminated med/biolog sub, transfused or infused
C1261338|[X]Contaminated medical or biological substances, transfused or infused (disorder)
C1261338|[X]Contaminated medical or biological substances, transfused or infused
C1261338|[X]Contaminated medical or biological substances, transfused or infused (finding)
C2108022|contamination during transfusion or infusion with bacteria (treatment)
C2108022|contamination during transfusion or infusion with bacteria
C2108032|contamination during transfusion or infusion with endotoxin-producing bacteria (treatment)
C2108032|contamination during transfusion or infusion with endotoxin-producing bacteria
C2108026|contamination during transfusion or infusion with virus (treatment)
C2108026|contamination during transfusion or infusion with virus
C2108013|contaminated blood, fluid, or drug during transfusion or infusion (treatment)
C2108013|contaminated blood, fluid, or drug during transfusion or infusion
C2108023|contamination during transfusion or infusion with bacterial pyogens (treatment)
C2108023|contamination during transfusion or infusion with bacterial pyogens
C2108024|contamination during transfusion or infusion with hepatotoxic substance
C2108024|contamination during transfusion or infusion with hepatotoxic substance (treatment)
C2108025|contamination during transfusion or infusion with viral hepatitis (treatment)
C2108025|contamination during transfusion or infusion with viral hepatitis
C0030275|Graftings, Pancreas
C0030275|Pancreas Grafting
C0030275|Pancreas Graftings
C0030275|Pancreas Transplantation
C0030275|Pancreas Transplantations
C0030275|Transplantations, Pancreas
C0030275|PANCREAS TRANSPL
C0030275|TRANSPL PANCREAS
C0030275|pancreatic transplantation
C0030275|pancreatic transplantation (treatment)
C0030275|Pancreat transplant NOS
C0030275|Pancreas transplant
C0030275|Transplantation of pancreas NOS
C0030275|Transplantation of pancreas NOS (procedure)
C0030275|Pancreatic transplant
C0030275|Pancreatic transplant (procedure)
C0030275|Pancreas Transplantation Procedures
C0030275|Grafting, Pancreas
C0030275|Transplantation, Pancreas
C0030275|Transplantation of pancreas
C0030275|Transplantation of pancreas (procedure)
C0030275|Transplantation of pancreas, NOS
C0030275|Pancreatic transplant, not otherwise specified
C0030275|Transplant of pancreas
C0024128|Graftings, Lung
C0024128|Lung Grafting
C0024128|Lung Graftings
C0024128|Lung Transplantation
C0024128|Lung Transplantations
C0024128|Transplantations, Lung
C0024128|Lung transplant
C0024128|LUNG TRANSPL
C0024128|TRANSPL LUNG
C0024128|lung transplant (treatment)
C0024128|surgery lung transplant
C0024128|Lung transplant NOS
C0024128|Transplant of lung
C0024128|Transplantation of lung NOS
C0024128|Transplantation of lung NOS (procedure)
C0024128|Lung transplant (procedure)
C0024128|Lung Transplantation Procedures
C0024128|Lungs--Transplantation
C0024128|Cardio/pulm: Lung transplant
C0024128|Grafting, Lung
C0024128|Transplantation, Lung
C0024128|LTx - Lung transplant
C0024128|Transplant of lung (procedure)
C0024128|Transplant of lung, NOS
C0024128|Lung transplantation, not otherwise specified
C0024128|En bloc lung transplantation
C0024128|Transplant;lung
C0018833|Grafting, Heart Lung
C0018833|Graftings, Heart-Lung
C0018833|Heart Lung Transplantation
C0018833|Heart-Lung Grafting
C0018833|Heart-Lung Graftings
C0018833|Heart-Lung Transplantation
C0018833|Heart-Lung Transplantations
C0018833|Transplantation, Heart Lung
C0018833|Transplantations, Heart-Lung
C0018833|Heart and lung transplant
C0018833|TRANSPL HEART LUNG
C0018833|HEART LUNG TRANSPL
C0018833|heart-lung transplant
C0018833|heart-lung transplant (treatment)
C0018833|Heart & lung transplant
C0018833|Comb heart/lung transpla
C0018833|Heart and heart-lung transplant
C0018833|Heart and heart-lung transplant (procedure)
C0018833|Transplantation of heart and lung NOS (procedure)
C0018833|Transplantation of heart and lung NOS
C0018833|Heart and heart-lung transplantation
C0018833|Heart/Lung Transplantation Procedures
C0018833|Grafting, Heart-Lung
C0018833|Transplantation, Heart-Lung
C0018833|HLTx - Heart lung transplant
C0018833|Heart Lung Grafting
C0018833|Heart and Lung Transplantation
C0018833|Combined heart-lung transplantation
C0730400|solid organ transplant (treatment)
C0730400|Solid organ transplant
C0730400|Solid organ transplant (procedure)
C0401176|renal transplant cadaveric donor
C0401176|cadaveric donor renal transplant (treatment)
C0401176|cadaveric donor renal transplant
C0401176|Cadaver renal allograft
C0401176|Cadaver renal allotransplant
C0401176|Cadaveric renal transplant
C0401176|Cadaveric renal transplant (procedure)
C0194034|spleen transplantation
C0194034|Spleen transplant
C0194034|Spleen transplant (procedure)
C0194034|Transplantation of spleen
C0194034|Transplantation of spleen (procedure)
C0022671|Kidney Grafting
C0022671|Kidney Transplantation
C0022671|Kidney Transplantations
C0022671|Renal Transplantations
C0022671|Transplantations, Kidney
C0022671|Transplantations, Renal
C0022671|Kidney transplant
C0022671|Renal transplant
C0022671|KIDNEY TRANSPL
C0022671|RENAL TRANSPL
C0022671|TRANSPL RENAL
C0022671|TRANSPL KIDNEY
C0022671|renal transplantation
C0022671|renal transplant (treatment)
C0022671|Transplantation of kidney NOS (procedure)
C0022671|Transplantation of kidney NOS
C0022671|Renal transplant (procedure)
C0022671|Renal Transplantation Procedures
C0022671|Kidneys--Transplantation
C0022671|Transplantation, Kidney
C0022671|Transplantation, Renal
C0022671|Grafting, Kidney
C0022671|Transplant of kidney
C0022671|Renal graft
C0022671|Transplantation of kidney
C0022671|Tx - Kidney transplantation
C0022671|Tx - Renal transplantation
C0022671|Transplant of kidney (procedure)
C0022671|Transplant of kidney, NOS
C0022671|Kidney transplantation, NOS
C0022671|Renal transplant, NOS
C0022671|Kidney Transplants
C0022671|Transplant;renal
C0023911|Graftings, Liver
C0023911|Hepatic Transplantations
C0023911|Liver Grafting
C0023911|Liver Graftings
C0023911|Liver Transplantation
C0023911|Liver Transplantations
C0023911|Transplantations, Hepatic
C0023911|Transplantations, Liver
C0023911|Liver transplant
C0023911|Hepatic Transplantation
C0023911|Transplantation of Liver
C0023911|TRANSPL HEPATIC
C0023911|HEPATIC TRANSPL
C0023911|TRANSPL LIVER
C0023911|LIVER TRANSPL
C0023911|liver transplant (treatment)
C0023911|Transplantation of liver NOS
C0023911|Transplantation of liver NOS (procedure)
C0023911|Liver transplant (procedure)
C0023911|Liver Transplantation Procedures
C0023911|Liver--Transplantation
C0023911|Grafting, Liver
C0023911|Transplantation, Liver
C0023911|Transplantation, Hepatic
C0023911|Tx - Liver transplantation
C0023911|LTx - Liver transplant
C0023911|Transplantation of liver (procedure)
C0023911|Transplantation of liver, NOS
C0023911|Transplant;liver
C0018823|Cardiac Transplantations
C0018823|Graftings, Heart
C0018823|Heart Grafting
C0018823|Heart Graftings
C0018823|Heart Transplantation
C0018823|Heart Transplantations
C0018823|Transplantations, Cardiac
C0018823|Transplantations, Heart
C0018823|Heart transplant
C0018823|TRANSPL CARDIAC
C0018823|CARDIAC TRANSPL
C0018823|TRANSPL HEART
C0018823|HEART TRANSPL
C0018823|transplantation of heart
C0018823|transplantation of heart (treatment)
C0018823|Cardiac Transplantation
C0018823|Transplant;cardiac
C0018823|Heart transplant (procedure)
C0018823|Heart--Transplantation
C0018823|CARDIAC TRANSPLANT
C0018823|Cardio/pulm: Heart transplant
C0018823|Grafting, Heart
C0018823|Transplantation, Heart
C0018823|Transplantation, Cardiac
C0018823|CTx - Cardiac transplant
C0018823|HTx - Heart transplant
C0018823|HtTx - Heart transplant
C0018823|Transplantation of heart (procedure)
C0018823|Transplantation of heart, NOS
C0018823|Heart Transplants
C0857825|Infection in solid organ transplant recipients
