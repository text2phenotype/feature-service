C0019029|Hemoglobin concentration result
C0019046|Hemoglobin
C0518015|Hemoglobin measurement
C0019018|Glycosylated hemoglobin A
C0202054|Glucohemoglobin measurement
C0373638|GLYCATED HEMOGLOBIN TEST
C0019018|Glycosylated hemoglobin A
C0202054|Glucohemoglobin measurement
C0373638|GLYCATED HEMOGLOBIN TEST
C3829717|Hemoglobin A1C to Hemoglobin Ratio Measurement
C0239940|Glycosylated haemoglobin increased
C0366781|Hemoglobin A1c/Hemoglobin total
C0366782|Hemoglobin A1c/Hemoglobin total
C0474680|Hemoglobin A1c measurement
C0800962|Hemoglobin A1c/Hemoglobin total
C0800963|Hemoglobin A1c/Hemoglobin total
C0806334|Hemoglobin A1c/Hemoglobin total
C1261236|Hemoglobin A1c level result
C1318607|HBA1c target
C1869903|hemoglobin A1c protein, human
C2114346|hemoglobin A1C level less than 7.0%
C2114374|hemoglobin A1C results documented and reviewed - hemoglobin A1C level greater 9.0%
C2707530|Hemoglobin A1c:-:Pt:Bld:-
C2733523|Ordinal level of hemoglobin A1c (observable entity)
C2919483|High hemoglobin A1c level
C2923665|Hemoglobin A1c/Hemoglobin total
C2973266|Hemoglobin A1c/Hemoglobin total
C3484089|Hemoglobin A1c/Hemoglobin total
C4073162|Elevated hemoglobin A1c
C4274658|Hemoglobin A1C test not done
C4315035|Elevated hemoglobin A1c (HbA1c)
C4325149|home hemoglobin A1C monitor
C4505389|Glycated Hemoglobin A1c
C0555792|Hemoglobin A1C - diabetic control interpretation
C1287394|Hemoglobin A1C - diabetic control finding
C1624104|Hemoglobin A1c:MCnc:Pt:Bld:Qn
C1624124|HbA1c measurement device panel
C2012263|hemoglobin A1C measurement using home device
C2114347|hemoglobin A1C level 7.0-9.0%
C2114373|hemoglobin A1C results documented and reviewed
C3838427|blood hemoglobin A1c/total ratio
C1737720|Most recent hemoglobin A1c level > 9.0% (DM)
C1964112|Most recent hemoglobin A1c (HbA1c) level less than 7.0% (DM)
C2732640|Calculation of estimated average glucose based on hemoglobin A1c
C2925136|Hemoglobin A1c 
C3838424|blood hemoglobin A1c/total ratio by HPLC
C3838425|blood hemoglobin A1c/total ratio by electrophoresis
C3838426|blood hemoglobin A1c/total ratio by calculation
C4028083|patient goals - keep hemoglobin a1c levels under ___
C4325143|HOME HEMOGLOBIN A1C MONITOR MISCELL EACH
C0438276|Hemoglobin A1c less than 7% indicating good diabetic control
C0438277|Hemoglobin A1c between 7%-10% indicating borderline diabetic control
C0438278|Hemoglobin A1c greater than 10% indicating poor diabetic control
C1277712|HbA1c measurement (DCCT aligned)
C1611204|Hemoglobin; glycosylated (A1C) by device cleared by FDA for home us
C1964113|Most recent hemoglobin A1c (HbA1c) level 7.0-9.0% (DM)
C4281023|Hemoglobin A1c greater than 9% indicating poor diabetic control
C4281024|Hemoglobin A1c between 7%-9% indicating borderline diabetic control
C4304316|Provision of written information about diabetes and high hemoglobin A1c level
C2960128|Hemoglobin A1c target value using International Federation of Clinical Chemistry and Laboratory Medicine standardized metho
C0007061|Carboxyhemoglobin
C0007061|Hemoglobins, carbonyl-
C0007061|Carbonyl hemoglobin
C0007061|Carbonyl haemoglobin
C0007061|Carbomonoxyhemoglobin
C0007061|Carbonmonoxyhemoglobin
C0007061|Carbonylhemoglobin
C0007061|Carboxyhemoglobin [Chemical/Ingredient]
C0007061|Carbonyl hemoglobin (substance)
C0007061|COHb
C0007061|Carbon monoxide hemoglobin
C0007061|Carbon monoxide haemoglobin
C0007061|Carboxyhaemoglobin
C0007061|HbCO - Carboxyhaemoglobin
C0007061|HbCO - Carboxyhemoglobin
C0007061|Carboxyhemoglobin (substance)
C0007061|COHbon monoxide hemoglobin
C0019016|A, Hemoglobin
C0019016|Hemoglobin A
C0019016|Hb alpha2 beta2
C0019016|Hb alpha<sub>2</sub> beta<sub>2</sub>
C0019016|HBA
C0019016|Hemoglobin A [Chemical/Ingredient]
C0019016|Hb A
C0019016|Haemoglobin A
C0019016|Hb A - Haemoglobin A
C0019016|Hb A - Hemoglobin A
C0019016|Hb alpha>2< beta>2<
C0019016|Hemoglobin A (substance)
C0019020|C, Hemoglobin
C0019020|Hemoglobin C
C0019020|HBC
C0019020|Hemoglobin C [Chemical/Ingredient]
C0019020|Haemoglobin C
C0019020|Hb C - Haemoglobin C
C0019020|Hb C - Hemoglobin C
C0019020|Hb 6 (A3), Glu-lys, beta chain
C0019020|Hemoglobin C (substance)
C0019020|Hb 6(A3), Glu-lys, beta chain
C0019020|Hb 6(A3), Glu-lys
C0015936|Fetal Hemoglobin
C0015936|Hemoglobin F
C0015936|Hemoglobin, Fetal
C0015936|Hb alpha2 gamma2
C0015936|Hb alpha<sub>2</sub> gamma<sub>2</sub>
C0015936|HBF
C0015936|Foetal haemoglobin
C0015936|Fetal Hemoglobin [Chemical/Ingredient]
C0015936|Hb F
C0015936|Haemoglobin F
C0015936|Hemoglobin.fetal
C0015936|Hb F - Haemoglobin F
C0015936|Hb F - Hemoglobin F
C0015936|Hb alpha>2< gamma>2<
C0015936|Fetal haemoglobin
C0015936|Hemoglobin F (substance)
C0019026|H, Hemoglobin
C0019026|Hemoglobin H
C0019026|Hb beta4
C0019026|Hb beta<sub>4</sub>
C0019026|HBH
C0019026|Hemoglobin H [Chemical/Ingredient]
C0019026|Haemoglobin H
C0019026|Hb beta>4<
C0019026|Hemoglobin H (substance)
C0019043|Hemoglobin, Sickle
C0019043|S, Hemoglobin
C0019043|Sickle Hemoglobin
C0019043|hemoglobin S
C0019043|HBS
C0019043|Haemoglobin S -RETIRED-
C0019043|Hemoglobin S -RETIRED-
C0019043|Hemoglobin, Sickle [Chemical/Ingredient]
C0019043|Haemoglobin S
C0019043|Hemoglobin S (substance)
C0019043|Haemoglobin S (substance)
C0019043|Hb S
C0019043|HbS hemoglobin
C0019043|Hb S - Haemoglobin S
C0019043|Hb S - Hemoglobin S
C0019043|Sickle haemoglobin
C0019043|Hb 6 (A3), Glu-val
C0019043|Hb 6(A3), Glu-val
C0025635|Methemoglobin
C0025635|Hemoglobins, met-
C0025635|Methemoglobin [Chemical/Ingredient]
C0025635|Ferrihemoglobin
C0025635|Methaemoglobin
C0025635|Methemoglobin (substance)
C0030069|Oxyhemoglobins
C0030069|oxyhemoglobin
C0030069|O2 Hb
C0030069|O<sub>2</sub>Hb
C0030069|Oxyhemoglobins [Chemical/Ingredient]
C0030069|Oxyhaemoglobin
C0030069|HbO2 - Oxyhaemoglobin
C0030069|HbO2 - Oxyhemoglobin
C0030069|O>2<Hb
C0030069|Oxyhemoglobin (substance)
C2353985|OxyVita
C2350441|Subunits, Hemoglobin
C2350441|Hemoglobin Subunits
C2350441|Hemoglobin Subunits [Chemical/Ingredient]
C0014764|Erythrocruorins
C0014764|Erythrocruorins [Chemical/Ingredient]
C0019047|Hemoglobins, Abnormal
C0019047|ABNORM HEMOGLOBINS
C0019047|HEMOGLOBINS ABNORM
C0019047|Abnormal hemoglobin NOS
C0019047|Hemoglobins, Abnormal [Chemical/Ingredient]
C0019047|Abnormal Hemoglobins
C0019047|Abnormal haemoglobin
C0019047|Abnormal hemoglobin
C0019047|Abnormal hemoglobin (substance)
C0019047|Abnormal hemoglobin, NOS
C0038731|Sulfhemoglobin
C0038731|Hemoglobins, sulf-
C0038731|Sulfhemoglobin [Chemical/Ingredient]
C0038731|Sulphaemoglobin
C0038731|Sulfemoglobin
C0038731|Sulfhemoglobin (substance)
C0038731|SulfHb
C0038731|SulphHb
C0038731|Sulfhaemoglobin
C0038731|Sulfhemoglobin [dup] (substance)
C0019046|Hemoglobin
C0019046|Hemoglobins
C0019046|Hemoglobins [Chemical/Ingredient]
C0019046|Hgb
C0019046|Hb
C0019046|Haemoglobin
C0019046|Hb - Haemoglobin
C0019046|Hb - Hemoglobin
C0019046|HGB - Haemoglobin
C0019046|HGB - Hemoglobin
C0019046|Hemoglobin (substance)
C0019046|Hemoglobin, NOS
C0019046|Haemoglobin, NOS
C1956056|Truncated Hemoglobins
C1956056|Hemoglobin, Truncated
C1956056|Hemoglobins, TrHb
C1956056|TrHb Hemoglobins
C1956056|Truncated Hemoglobins [Chemical/Ingredient]
C1956056|Truncated Hemoglobin
C1956056|Hemoglobins, Truncated
C0015891|Hemoglobin, Ferrous
C0015891|Ferrous Hemoglobin
C2935533|non-symbiotic hemoglobin 1 protein, rice
C2935533|non-symbiotic hemoglobin 1 protein, Oryza sativa
C2935621|HBOC-205LL.LT.MW600
C0057437|deoxyhemoglobin
C0057437|Hb(T)
C0057437|T-state hemoglobin
C0057437|HHb
C0057437|MetHb
C0057437|Reduced hemoglobin
C0057437|Deoxyhaemoglobin
C0057437|Reduced haemoglobin
C0057437|Deoxyhemoglobin (substance)
C0019035|SS, Hemoglobin
C0019035|Hemoglobin SS
C0052175|apohemoglobin
C0062119|haptoglobin-hemoglobin complex
C0062119|hemoglobin-haptoglobin complex
C0062418|Hb P
C0062418|hemoglobin P
C0063048|hybrid hemoglobins
C0121409|hemorphin 6
C0121409|hemorphin-6
C0534165|S-nitrosohemoglobin
C0534165|S-Nitrosated Hemoglobin
C0534165|S-Nitroso-Hemoglobin
C0534165|S-nitrosylhemoglobin
C0056041|cobalt hemoglobin
C0056041|coboglobin
C0068873|Hb X
C0068873|nitrosyl hemoglobin
C0068873|nitrosylhemoglobin
C0068873|nitrosylferrohemoglobin
C0056649|cyanhemoglobin
C0056649|cyanohemoglobin
C0056649|hemoglobin cyanide
C0062478|hemoglobin, stroma free
C0062478|SFHb
C0062478|stroma-free hemoglobin
C0062248|Hb B
C0062248|hemoglobin B
C0071588|PLP-Hb
C0071588|poly Hb-PLP
C0071588|polyhemoglobin-pyridoxal-5-phosphate
C0071588|pyridoxal phosphate modified hemoglobin
C0071588|pyridoxalated polymerized hemoglobin
C0071588|p-polyHb
C0071588|polymerized pyridoxylated hemoglobin
C0142130|poly SFH-P
C0142130|SFH-PLP
C0142130|SFHB-PP
C0142130|pyridoxalated polymerized stroma-free hemoglobin
C0056024|cobalt deoxyhemoglobin
C0056024|deoxycobalthemoglobin
C0056024|Hemoglobin A, cobalto-
C0071587|poly Hb
C0071587|polyhemoglobin
C0057619|dextran-hemoglobin
C0057619|dextran-hemoglobin complex (deoxygenated)
C0057619|DHCDO
C0108535|carp-human hybrid hemoglobin
C0065652|manganese-iron hybrid hemoglobin
C0065652|Mn-Fe(II) hybrid Hb
C0123968|Co-Fe(II) hybrid Hb
C0123968|cobalt-iron hybrid hemoglobin
C0123968|iron-cobalt hybrid hemoglobin
C0062487|hemorphin 4
C0062487|hemorphin-4
C0062487|L-Threonine, N-(N-(1-L-tyrosyl-L-prolyl)-L-tryptophyl)-
C0062487|Tyr-Pro-Trp-Thr
C0062487|tyrosyl-prolyl-tryptophyl-threonine
C0072711|PLP-Hb-PEG
C0072711|POE conjugated pyridoxalated hemoglobin
C0072711|polyoxyethylene conjugated pyridoxalate hemoglobin
C0072711|pyridoxalated-hemoglobin-polyethylene glycol conjugate
C0072711|pyridoxalated-hemoglobin-polyoxyethylene conjugate
C0072711|pyridoxylated hemoglobin-polyoxyethylene conjugated solution
C0072711|PHP conjugate
C0072711|pyridoxylated haemoglobin-polyoxyethylene conjugate
C0377989|PHP44 conjugate
C0377990|PHP88 conjugate
C0050784|adenosine triphosphate-stroma-free hemoglobin
C0050784|ATP-Hb
C0050784|ATP-SFH
C0078783|zinc hemoglobin
C0078783|Zn-Hb
C0052777|azidohemoglobin
C0052777|Hb N3
C0052777|hemoglobin azide
C0285562|Ni(II)-Fe(II) hybrid Hb
C0285562|alpha(Fe)(II)-beta(Ni)(II) hybrid Hb
C0285562|alpha(Ni)(II)-beta(Fe)(II) hybrid Hb
C0285562|nickel-iron hybrid hemoglobin
C0082846|alpha, alpha-Hb
C0082846|Hb-XL99alpha
C0082846|HbXL99alpha
C0082846|hemoglobin XL99alpha
C0082846|XLHb hemoglobin
C0082846|bis(3,5-dibromosalicyl)fumarate-cross-linked hemoglobin
C0121105|HbBv-FMDA
C0209012|Hb acetylated
C0209012|acetylated Hb
C0209012|acetylated hemoglobin
C0062476|4-aminobiphenylhemoglobin adduct
C0062476|4ABP-Hb
C0062476|hemoglobin, 4-aminobiphenyl-
C0245921|globin compound IV
C0245921|hemoglobin IV
C0102331|alpha(A) globin
C0102331|alpha(A) hemoglobin
C0109312|Chi t I allergen
C0109312|Chironomus thummi hemoglobin
C0109312|hemoglobin protein, Chironomus thummi
C0167672|Leu-Val-Val-Tyr-Pro-Trp-Thr-Gln-Arg-Phe
C0167672|LVV-hemorphin-7
C0167672|leucyl-valyl-valyl-tyrosyl-prolyl-tryptophyl-threonyl-glutaminyl-arginyl-phenylalanine
C0167672|LVV-H7
C0212463|Hb (64-76)
C0212463|hemoglobin (64-76)
C0215199|upbHb
C0215199|polymerized bovine hemoglobin
C0217022|HbBv-DVS
C0217022|bovine hemoglobin-divinyl sulfone
C0217024|poly HbBv-DVS
C0217024|polymerized bovine hemoglobin-divinyl sulfone
C0219010|Vitreoscilla hemoglobin
C0219010|VHb protein, Vitreoscilla
C0219010|hemoglobin protein, Vitreoscilla
C0219880|HbI, S. inaequivalvis
C0219880|homodimeric Hb, S. inaequivalvis
C0219880|dimeric hemoglobin, Scapharca inaequivalvis
C0247389|DCLHb
C0247389|diaspirin-cross-linked hemoglobin
C0250445|L-Phenylalanine, N-(N2-(N2-(N-(N-(1-L-tyrosyl-L-prolyl)-L-tryptophyl)-L-threonyl)-L-glutaminyl)-L-arginyl)-
C0250445|Tyr-Pro-Trp-Thr-Gln-Arg-Phe
C0250445|hemorphin 7
C0250445|hemorphin-7
C0250445|tyrosyl-prolyl-tryptophyl-threonyl-glutaminyl-arginyl-phenylalanine
C0251387|Hb18 peptide
C0251387|hemoglobin 18 peptide
C0251389|Hba11 peptide
C0251389|hemoglobin a11 peptide
C0252834|Urechis caupo Hb
C0252834|Urechis caupo hemoglobin
C0252834|hemoglobin, Urechis caupo
C0254489|LI410 protein, Chlamydomonas eugametos
C0254491|LI637 protein, Chlamydomonas eugametos
C0299241|VV-hemorphin-7
C0299241|Val-Val-Tyr-Pro-Trp-Thr-Gln-Arg-Phe
C0299241|valyl-valyl-tyrosyl-prolyl-tryptophyl-threonyl-glutaminyl-arginyl-phenylalanine
C0300427|Hb, T. heterochaetus
C0300427|hemoglobin, Tylorrhynchus
C0381552|Dex-BTC-Hb
C0381552|Hb-dex-BTC
C0381552|dextran 10-benzene-tetracarboxylate-hemoglobin
C0381552|dextran-benzene-tetra-carboxylate hemoglobin
C0381552|hemoglobin-dextran 10-benzene-tetracarboxylate
C0381551|benzene tetracarboxylate substituted dextran
C0384641|O-raffinose cross-linked human hemoglobin
C0384641|O-raffinose cross-linked oligomeric hemoglobin
C0384641|o-R-poly-Hb
C0384641|hemoglobin-raffimer
C0388973|fumaryl beta,beta-CLHb
C0388973|fumaryl beta,beta-crosslinked hemoglobin
C0389721|MgII-FeII Hb
C0389721|MgII-FeII hemoglobin
C0389721|magnesium-iron hemoglobin
C0389849|deoxy-des-alpha-Arg(141)-Hb
C0389849|deoxy-des-alpha-arginine(141) hemoglobin
C0535034|HBII B SI
C0535035|HbII A SI
C0535038|HbII, S. inaequivalvis
C0535038|tetrameric Hb, S. inaequivalvis
C0535038|tetrameric hemoglobin, Scapharca inaequivalvis
C0082471|erythrocruorin
C0017853|Glycosylated Hemoglobin
C0017853|Hemoglobin, Glycosylated
C0017853|Hemoglobins, Glycated
C0017853|Glycosylated Hb
C0017853|Glycated hemoglobin
C0017853|Glycated haemoglobin
C0017853|Hemoglobin.glycated
C0017853|Glycated Hemoglobins
C0017853|Glycosylated haemoglobin
C0017853|Glycosylated hemoglobin (substance)
C0018927|Hematin
C0018927|Haematin
C0018927|Ferriporphyrin hydroxide
C0018927|Ferriprotoporphyrin basic
C0018927|Hematin (substance)
C0018927|Hydroxyhemin
C0018988|Chloride, Ferriheme
C0018988|Chloride, Ferriprotoporphyrin IX
C0018988|Hemin
C0018988|Ferrate(2-), chloro(7,12-diethenyl-3,8,13,17-tetramethyl-21H,23H-porphine-2,18-dipropanoato(4-)-N21,N22,N23,N24)-, dihydrogen, (SP-5-13)-
C0018988|Hemin (product)
C0018988|Hemin agent
C0018988|Haemin agent
C0018988|Haemin
C0018988|enzyme inhibitors hemin
C0018988|hemin (medication)
C0018988|Protohemin
C0018988|Ferriheme Chloride
C0018988|Hemin [Chemical/Ingredient]
C0018988|Chlorohemin
C0018988|Protohemin IX
C0018988|Ferriprotoporphyrin IX Chloride
C0018988|Haemin preparation
C0018988|Hemin (substance)
C0018988|Hemin agent (substance)
C0018988|Hemin preparation
C0018988|Hemin preparation (substance)
C0055513|choleglobin
C0055513|Verdoglobin
C0055513|Verdoglobin (substance)
C0055513|Verdohemoglobin
C0055513|Verdohaemoglobin
C0055513|Verdohemoglobin (substance)
C0018966|Heme
C0018966|Ferrate(2-), (7,12-diethenyl-3,8,13,17-tetramethyl-21H,23H-porphine-2,18-dipropanoato(4-)-N21,N22,N23,N24)-, dihydrogen, (SP-4-2)-
C0018966|ferroheme
C0018966|Ferroprotoporphyrin
C0018966|Protoheme IX
C0018966|Heme [Chemical/Ingredient]
C0018966|Haem
C0018966|Heme b
C0018966|Protoheme
C0018966|Hemes
C0018966|Reduced Hematin
C0018966|Hematein
C0018966|Benz(b)indeno(1,2-d)pyran-9(6h)-one, 6a,7-dihydro-3,4,6a,10-tetrahydroxy-
C0018966|Hematin
C0018966|Heme Group
C0018966|Haeme
C0018966|Heme (substance)
C0018966|Hem
C0019024|E, Hemoglobin
C0019024|Hemoglobin E
C0019024|HBE
C0019024|Hemoglobin E [Chemical/Ingredient]
C0019024|Hemoglobin E (substance)
C0019024|HbE - Haemoglobin E
C0019024|HbE - Hemoglobin E
C0019024|Haemoglobin E
C0019024|Hb E - Hemoglobin E
C0019024|Hb E - Haemoglobin E
C0019024|Hb 26 (B8), Glu-lys, beta chain
C0019024|Hb 26(B8), Glu-lys, beta chain
C0019024|Hemoglobin E [dup] (substance)
C3687697|Hemoglobin glutamer-200 (bovine) (substance)
C3687697|Hemoglobin glutamer-200 (bovine)
C3478324|Hemoglobin &#x7C; Pericardial fluid
C1988924|Hemoglobin &#x7C; reticulocytes
C1988928|Hemoglobin &#x7C; XXX
C2736165|Hgb Ur Ql Strip.auto
C2736165|Hemoglobin:ACnc:Pt:Urine:Ord:Test strip.automated
C2736165|Hemoglobin [Presence] in Urine by Automated test strip
C2736165|Hemoglobin:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip.automated
C2965248|Hemoglobin &#x7C; fetus &#x7C; Bld-Ser-Plas
C1988917|Hemoglobin &#x7C; blood venous
C1988926|Hemoglobin &#x7C; synovial fluid
C3854324|Hemoglobin.free
C3854324|Free hemoglobin (substance)
C3854324|Free hemoglobin
C3854324|Free haemoglobin
C0362931|Hemoglobin:MCnc:Pt:Urine:Qn
C0362931|Hemoglobin [Mass/volume] in Urine
C0362931|Hgb Ur-mCnc
C0362931|Hemoglobin:Mass Concentration:Point in time:Urine:Quantitative
C0368020|Hemoglobin:ACnc:Pt:Urine:Ord:Test strip
C0368020|Hgb Ur Ql Strip
C0368020|Hemoglobin [Presence] in Urine by Test strip
C0368020|Hemoglobin:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C1988919|Hemoglobin &#x7C; cerebral spinal fluid
C1988914|Hemoglobin &#x7C; blood cord arterial
C1988913|Hemoglobin &#x7C; blood cord
C2587436|Hemoglobin &#x7C; Blood product unit &#x7C; Bld-Ser-Plas
C1988915|Hemoglobin &#x7C; blood cord venous
C1988910|Hemoglobin &#x7C; bld-ser-plas
C1988927|Hemoglobin &#x7C; urine
C1988922|Hemoglobin &#x7C; pleural fluid
C1988911|Hemoglobin &#x7C; blood arterial
C1988921|Hemoglobin &#124; peritoneal fluid
C1988921|Hemoglobin &#x7C; peritoneal fluid
C1988916|Hemoglobin &#x7C; blood mixed venous
C1988912|Hemoglobin &#x7C; blood capillary
C1988918|Hemoglobin &#x7C; body fluid
C1978486|Hemoglobin [Mass/volume] in Urine by Automated test strip
C1978486|Hgb Ur Strip.auto-mCnc
C1978486|Hemoglobin:MCnc:Pt:Urine:Qn:Test strip.automated
C1978486|Hemoglobin:Mass Concentration:Point in time:Urine:Quantitative:Test strip.automated
C1954901|Hemoglobin [Mass/volume] in Urine by Test strip
C1954901|Hgb Ur Strip-mCnc
C1954901|Hemoglobin:MCnc:Pt:Urine:Qn:Test strip
C1954901|Hemoglobin:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C3657113|polyhemoglobin-superoxide dismutase-catalase-carbonic anhydrase
C3657113|PolySFHb-SOD-CAT-CA
C3529748|Hb 98-114, bovine
C3529748|hemoglobin (98-114), bovine
C3490724|polypeptide-Fe
C3180469|polynitroxylated pegylated hemoglobin
C3883879|RVDPVNFKLLSH
C3883879|Arg-Val-Asp-Pro-Val-Asn-Phe-Lys-Leu-Leu-Cys-His
C3883879|RVD-hemopressin, human
C4045299|YQ23 compound
C4042582|alpha1-32 Hb, bovine
C4042582|hemoglobin alpha-chain (1-32), bovine
C0014730|Eryhem
C4078062|HbAHP-25
C0019030|Hemoglobin M
C0019030|M, Hemoglobin
C0019030|HBM
C0019030|Hemoglobin M [Chemical/Ingredient]
C0019030|Haemoglobin M
C0019030|Hb M - Haemoglobin M
C0019030|Hb M - Hemoglobin M
C0019030|Hemoglobin M (substance)
C0062251|Hb Bart's
C0062251|hemoglobin Bart's
C0062251|hemoglobin Barts
C0062251|methemoglobin Bart's
C0062251|Hemoglobin Bart
C0062251|Haemoglobin Bart
C0062251|Haemoglobin Barts
C0062251|Hb - Haemoglobin Barts
C0062251|Hb - Hemoglobin Barts
C0062251|Hemoglobin Bart (substance)
C0019018|Hemoglobin A, Glycosylated
C0019018|Glycosylated hemoglobin A
C0019018|HbA1c
C0019018|HBA GLYCOSYLATED
C0019018|HBA 01
C0019018|HEMOGLOBIN AA 01
C0019018|HB AC 01
C0019018|Haemoglobin A1c
C0019018|HbA>1c<
C0019018|Hemoglobin A1c
C0019018|HbA<sub>1c</sub>
C0019018|Hemoglobin A, Glycosylated [Chemical/Ingredient]
C0019018|Hb A1a+b
C0019018|Glycohemoglobin A
C0019018|HbA1
C0019018|Hemoglobin A(1)
C0019018|Hb A1
C0019018|Hb A1c
C0019018|HbA<sub>1c</sub> (substance)
C0019018|HbA1c (substance)
C0019018|HbA>1c< (substance)
C0019018|HbA1 - Glycated haemoglobin
C0019018|HbA1 - Glycated hemoglobin
C0019018|Glycosylated haemoglobin A
C0019018|Glycosylated hemoglobin A (substance)
C0313267|HEMOGLOBIN, ALKALI RESISTANT
C0313267|Alkali-resistant hemoglobin
C0313267|Alkali-resistant haemoglobin
C0313267|Alkali-resistant hemoglobin (substance)
C0313266|Ferri-hemoglobin
C0313266|Ferri-haemoglobin
C0313266|Ferri-hemoglobin (substance)
C0313263|Hemoglobin A,a
C0313263|Haemoglobin A,a
C0313263|Hemoglobin A,a (substance)
C0313264|Hemoglobin A,b
C0313264|Haemoglobin A,b
C0313264|Hemoglobin A,b (substance)
C0301731|hemoglobin Gower I
C0301731|Hb epsilon4
C0301731|Hb epsilon<sub>4</sub>
C0301731|Hemoglobin Gower-1
C0301731|Haemoglobin Gower-1
C0301731|Hb epsilon>4<
C0301731|Hemoglobin Gower-1 (substance)
C0301731|Hb Gower I
C0301732|hemoglobin Gower II
C0301732|Hemoglobin alpha2 epsilon2
C0301732|Haemoglobin alpha2 epsilon2
C0301732|Haemoglobin alpha<sub>2</sub> epsilon<sub>2</sub>
C0301732|Hemoglobin alpha<sub>2</sub> epsilon<sub>2</sub>
C0301732|Hemoglobin Gower-2
C0301732|Haemoglobin Gower-2
C0301732|Haemoglobin alpha>2< epsilon>2<
C0301732|Hemoglobin alpha>2< epsilon>2<
C0301732|Hemoglobin Gower-2 (substance)
C0301732|Hb Gower II
C0301809|Verdochromogen
C0301809|Verdochromogen (substance)
C0443781|Globin chain
C0443781|Globin chain (substance)
C0019019|A2, Hemoglobin
C0019019|Hemoglobin A2
C0019019|Hb alpha2 delta2
C0019019|Haemoglobin A2
C0019019|Haemoglobin A<sub>2</sub>
C0019019|Hb alpha<sub>2</sub> delta<sub>2</sub>
C0019019|Hemoglobin A2 (substance)
C0019019|Hemoglobin A<sub>2</sub> (substance)
C0019019|Hemoglobin A<sub>2</sub>
C0019019|HBA2
C0019019|HEMOGLOBIN AA 02
C0019019|Hemoglobin A2 [Chemical/Ingredient]
C0019019|Hb A2 - Haemoglobin A2
C0019019|Hb A2 - Hemoglobin A2
C0019019|Hb alpha>2< delta>2<
C0019019|Haemoglobin A>2<
C0019019|Hemoglobin A>2<
C0019019|Hemoglobin A>2< (substance)
C0369310|Haemoglobin A3
C0369310|Hemoglobin A3
C0369310|Haemoglobin A<sub>3</sub>
C0369310|Hemoglobin A3 (substance)
C0369310|Hemoglobin A<sub>3</sub> (substance)
C0369310|Hemoglobin A<sub>3</sub>
C0369310|Haemoglobin A>3<
C0369310|Hemoglobin A>3<
C0369310|Hemoglobin A>3< (substance)
C0532041|cyanoglobin protein, Nostoc
C0603512|manganese hemoglobin
C0606551|dyshaemoglobins
C0606551|dyshemoglobins
C0606551|Dyshemoglobin
C0607103|N-ethylsuccinimide hemoglobin
C0607103|NES-Hb
C1448496|hemoglobin I, non-mammalian
C0612736|nitrosyl-deoxy asymetrical hybrid hemoglobin
C0612736|NDAH hemoglobin
C0071452|PLDTHC
C0071452|poly(lysinediylterephthaloyl)microcapsules
C0071452|poly(N(alpha),N(epsilon) L-lysinediylterephthaloyl)hemolysate capsules
C0613702|dansyl-hemoglobin
C0613702|DNS-Hb
C0618939|Pyr-Hb-inulin
C0618939|pyridoxyl-hemoglobin-inulin
C0618939|pyridoxylated hemoglobin-inulin
C0620678|TFE Cys(beta93)Hb
C0620678|trifluoroethyl-cysteine-beta93 hemoglobin
C0620678|TFEC93HB
C0623643|me-apoHb
C0623643|methyl apohemoglobin
C0628391|hemorphin 5
C0628391|hemorphin-5
C0628391|Tyr-Pro-Trp-Thr-Gln
C0635222|haemoglobin L
C0635222|Hb L
C0635222|Hemoglobin L
C0636206|Hb isothiocyanate
C0636206|hemoglobin isothiocyanate
C0636692|Hb alpha-chain fragments (123-136)
C0636692|hemoglobin alpha-chain fragments (123-136)
C0636692|Hb (123-136)
C0639350|dimeric hemoglobin, Calyptogena soyoae
C0639350|Hb I, Calyptogena soyoae
C0647545|LVV hemorphin-6
C0647545|LVV-hemorphin 6
C0647886|hemoglobin II, Casuarina glauca
C0647886|HBII protein, Casuarina glauca
C0647886|Hb II protein, Casuarina glauca
C0212332|hemoglobin polymer
C0659625|hemoglobin linker chain L1 protein, Lumbricus terrestris
C0661309|deoxyHB-DPG
C0661309|deoxyhaemoglobin-2,3-diphosphoglycerate complex
C0661576|Hb III, LP
C0661576|hemoglobin III, Lucina pectinata
C0252444|polyHb-SOD-catalase
C0252444|polyhemoglobin-superoxide dismutase-catalase
C0252444|polyHb-SOD-CAT
C1611853|hemoglobin linker chain L2, Neanthes diversicolor
C0383956|HBOC 201
C0383956|HBOC-201
C0383956|hemoglobin-based oxygen carrier-201
C0383956|hemoglobin glutamer-250
C1308309|GLB2 protein, Arabidopsis
C1308309|AHB2 protein, Arabidopsis
C0669866|polyethylene glycol-hemoglobin conjugate
C0669866|PEG-Hb
C0669866|PEG-hemoglobin
C0673757|exorphin C
C0673757|Tyr-Pro-Ile-Ser-Leu
C0673757|tyrosyl-prolyl-isoleucyl-seryl-leucine
C0759385|bis(3,5-dibromosalicyl)sebacate-crosslinked hemoglobin
C0759385|DBBS-Hb
C0909600|Ascaris haemoglobin
C0909600|hemoglobin, Ascaris
C0909654|PNH-Hb
C0909654|polynitroxyl alphaalpha-hemoglobin
C0909654|polynitroxyl hemoglobin
C0911144|hemoglobin-based oxygen carrier-200
C0911144|HBOC-200
C0911144|hemoglobin glutamer-200
C0912247|glutathionyl hemoglobin
C0912247|GSH-Hb
C0912753|Hb Mermis
C0912753|hemoglobin, Mermis nigrescens
C1309473|glbN protein, Synechocystis
C1309473|slr2097 protein, Synechocystis
C0914187|Hb II, C. kaikoi
C0914187|hemoglobin II, Calyptogena
C1309669|Mhb1 protein, Medicago sativa
C1309669|non-symbiotic hemoglobin 1 protein, Medicago sativa
C0965761|3ABP-Hb
C0965761|hemoglobin, 3-aminobiphenyl-
C1120100|Hb FS hemoglobin
C1120100|alpha2gammabetaS
C1122894|erythrogen
C1173496|class 1 hemoglobin, Arabidopsis
C1173496|GLB1 protein, Arabidopsis
C1173496|AHB1 protein, Arabidopsis
C1174169|LVV-H4
C1174169|LVV-hemorphin-4
C1175813|PVNFKFLSH
C1175813|hemopressin
C1176132|MP4 PEG-Hb conjugate
C1176132|PEG-Hb conjugate, MP4
C1258934|HBOC rHB2.0, human
C1258934|hemoglobin-based oxygen carrier rHB2.0, human
C1453434|LVV-hemorphin-5
C1453434|Leu-Val-Val-Tyr-Pro-Trp-Thr-Gln
C1453434|leucyl-valyl-valyl-tyrosyl-prolyl-tryptophyl-threonyl-glutaminyl
C1453435|VV-hemorphin-5
C1453435|Val-Val-Tyr-Pro-Trp-Thr-Gln
C1453435|valyl-valyl-tyrosyl-prolyl-tryptophyl-threonyl-glutaminyl
C1504975|PolyHb-tyrosinase
C1504975|polyhemoglobin-tyrosinase
C1529786|MP4OX cpd
C1529786|MP4 (MalPEG-Hb)
C1529786|MalPEG-Hb, MP4
C1529786|maleimide-polyethylene glycol-modified hemoglobin, MP4
C1612076|Hb (107-136), bovine
C1612076|hemoglobin (107-136), bovine
C1700203|CG15180 protein, Drosophila
C1700203|Glob2 protein, Drosophila
C1701816|CG14675 protein, Drosophila
C1701816|Glob3 protein, Drosophila
C1700175|PolyHeme
C0387963|DHP I dehaloperoxidase
C0387963|dehaloperoxidase DHP I
C1872127|ferrylhemoglobin
C1872127|ferrylHb
C1872127|hemoglobin(Fe(IV)O)
C1999517|HRC 101
C2000553|PolyHb-Fg
C2000553|polyhemoglobin-fibrinogen
C0017645|Globin
C0017645|Globins
C0017645|Globins [Chemical/Ingredient]
C0518015|Haemoglobin
C0518015|Haem
C0518015|Hemoglobin Measurement
C0518015|hemoglobin
C0518015|hemoglobin measurement (lab test)
C0518015|Test;haemoglobin
C0518015|BLOOD COUNT HEMOGLOBIN
C0518015|Hemoglobin level
C0518015|Measurement of hemoglobin (Hgb)
C0518015|Hemoglobin determination (procedure)
C0518015|Hemoglobin determination
C0518015|Haemoglobin determination
C0518015|HGB
C0518015|Blood count; hemoglobin (Hgb)
C0518015|FHGB
C0518015|Free Hemoglobin
C0518015|Hemoglobin determination, NOS
C0518015|Haemoglobin determination, NOS
C0518015|Test;hemoglobin
C0518015|haemoglobin test
C0518015|hemoglobin test
C2825554|Percent Hemoglobin A
C2825554|Hemoglobin A to Total Hemoglobin Ratio Measurement
C2825555|Hemoglobin A2 to Total Hemoglobin Ratio Measurement
C2825555|Percent Hemoglobin A2
C2825556|Hemoglobin C to Total Hemoglobin Ratio Measurement
C2825556|Percent Hemoglobin C
C2825557|Percent Hemoglobin S
C2825557|Hemoglobin S to Total Hemoglobin Ratio Measurement
C2825557|Hemoglobin S Measurement
C1281911|Hemoglobin A measurement
C1281911|Hemoglobin A (& level)
C1281911|Haemoglobin A (& level)
C1281911|Haemoglobin A (& level) (procedure)
C1281911|Hemoglobin A
C1281911|HGBA
C1281911|Haemoglobin A level
C1281911|Haemoglobin A measurement
C1281911|Hemoglobin A level
C1281911|Hemoglobin A measurement (procedure)
C0474543|Hemoglobin A2 Measurement
C0474543|Hemoglobin A2 level
C0474543|Haemoglobin A2 level (procedure)
C0474543|Haemoglobin A2 level
C0474543|Hemoglobin A2
C0474543|HGBA2
C0474543|Haemoglobin A2
C0474543|Haemoglobin A2 measurement
C0474543|Hemoglobin A2 measurement (procedure)
C2984939|Hemoglobin B Measurement
C2984939|Hemoglobin B
C2984939|HGBB
C1275423|Hemoglobin C measurment
C1275423|Haemoglobin C measurement
C1275423|Measurement of haemoglobin C
C1275423|Haemoglobin C level (procedure)
C1275423|Measurement of hemoglobin C (procedure)
C1275423|Measurement of hemoglobin C
C1275423|Haemoglobin C
C1275423|Hemoglobin C Measurement
C1275423|Hemoglobin C
C1275423|HGBC
C1275423|Haemoglobin C level
C1275423|Hemoglobin C level
C0200695|Fetal hemoglobin determination
C0200695|Foetal haemoglobin
C0200695|Foetal hemoglobin determination
C0200695|Hemoglobin F Measurement
C0200695|Fetal hemoglobin level
C0200695|Hemoglobin F (& level)
C0200695|Haemoglobin F (& level) (procedure)
C0200695|Haemoglobin F (& level)
C0200695|HGBF
C0200695|Hemoglobin F
C0200695|Fetal Hemoglobin
C0200695|Haemoglobin F
C0200695|Foetal haemoglobin determination
C0200695|Haemoglobin F level
C0200695|Hemoglobin F level
C0200695|Fetal haemoglobin determination
C0200695|Fetal hemoglobin determination (procedure)
C0587341|Hb estimation
C0587341|Haemoglobin estimation
C0587341|Hemoglobin estimation
C0587341|Hemoglobin estimation NOS
C0587341|Haemoglobin estimation NOS
C0587341|Hemoglobin estimation (& level)
C0587341|Haemoglobin estimation (& level) (procedure)
C0587341|Hemoglobin estimation NOS (procedure)
C0587341|Haemoglobin estimation NOS (procedure)
C0587341|Haemoglobin estimation (& level)
C0587341|Haemoglobin estimation level
C0587341|Hemoglobin estimation level
C0587341|Haemoglobin level estimation
C0587341|Hb estimation (procedure)
C0587341|Hemoglobin level estimation (procedure)
C0587341|Hemoglobin level estimation
C3890034|Reticulocyte Hemoglobin Measurement
C3890034|Reticulocyte Hemoglobin
C3890034|Total Reticulocyte Corpuscular Hemoglobin Content Measurement
C3890034|CHr
C3890034|RETICH
C3890034|Ret. Corpuscular Hemoglobin Content
C0202133|Hemoglobin; methemoglobin, quantitative
C0202133|HEMOGLOBIN METHEMOGLOBIN QUANTITATIVE
C0202133|Methemoglobin measurement, quantitative
C0202133|Methaemoglobin measurement, quantitative
C0202133|Methemoglobin measurement, quantitative (procedure)
C0202133|BLOOD METHEMOGLOBIN ASSAY
C1611204|GLYCOSYLATED HB HOME DEVICE
C1611204|HGB GLYCOSYLATED DEVICE CLEARED FDA HOME USE
C1611204|Hemoglobin; glycosylated (A1C) by device cleared by FDA for home use
C0373637|FETAL HEMOGLOBIN ASSAY QUAL
C0373637|Hemoglobin; F (fetal), qualitative
C0373637|HEMOGLOBIN F FETAL QUALITATIVE
C0373637|Qualitative analysis of hemoglobin F (Hb F)
C0202132|Hemoglobin; methemoglobin, qualitative
C0202132|HEMOGLOBIN METHEMOGLOBIN QUALITATIVE
C0202132|Qualitative analysis of methemoglobin in hemoglobin
C0202132|Methemoglobin measurement, qualitative
C0202132|Methaemoglobin measurement, qualitative
C0202132|Methemoglobin measurement, qualitative (procedure)
C0202132|BLOOD METHEMOGLOBIN TEST
C0373638|Glycosylated haemoglobin
C0373638|GLYCATED HEMOGLOBIN TEST
C0373638|GLYCOSYLATED HEMOGLOBIN TEST
C0373638|HbA1c measurement
C0373638|hemoglobin A1C
C0373638|blood hemoglobin A1C measurement
C0373638|blood hemoglobin A1C measurement (lab test)
C0373638|blood glycosylated hemoglobin A1C measurement
C0373638|HEMOGLOBIN GLYCOSYLATED A1C
C0373638|Measurement of glycosylated hemoglobin (HbA1C)
C0373638|Glycohemoglobin
C0373638|Glycosylated hemoglobin
C0373638|Haemoglobin glycosylated
C0373638|HbA1C
C0373638|Hemoglobin glycosylated
C0373638|Glycohaemoglobin
C0373638|Glycosylated Hemoglobins Test
C0373638|Hemoglobin; glycosylated (A1C)
C0523686|Hemoglobin; thermolabile
C0523686|thermolabile hemoglobin
C0523686|thermolabile hemoglobin (lab test)
C0523686|Hemoglobin, thermolabile measurement
C0523686|thermolabile hemoglobin level
C0523686|HEMOGLOBIN THERMOLABILE
C0523686|Thermolabile (heat sensitive) hemoglobin level
C0523686|Haemoglobin, thermolabile measurement
C0523686|Hemoglobin, thermolabile measurement (procedure)
C0523686|ASSAY OF HEMOGLOBIN HEAT
C0236439|Hemoglobin; urine
C0236439|urine hemoglobin (lab test)
C0236439|urine hemoglobin
C0236439|Urine hemoglobin level
C0236439|ASSAY OF HEMOGLOBIN URINE
C0236439|Haemoglobin urine
C0236439|Urinary hemoglobin
C0236439|Urinary haemoglobin
C0236439|Hemoglobin urine
C0236439|Urine Hemoglobin Test
C0236439|ASSAY OF URINE HEMOGLOBIN
C0373636|Hemoglobin; F (fetal), chemical
C0373636|FETAL HEMOGLOBIN CHEMICAL
C0373636|HEMOGLOBIN F FETAL CHEMICAL
C0373636|Chemical analysis of hemoglobin F
C0373635|Hemoglobin; by copper sulfate method, non-automated
C0373635|HEMOGLOBIN COPPER SULFATE
C0373635|HEMOGLOBIN COPPER SULFATE METHOD NON-AUTOMATED
C0373635|Hemoglobin by copper sulfate method, non-automated
C0373635|Haemoglobin by copper sulphate method, non-automated
C0373635|Hemoglobin by copper sulfate method, non-automated (procedure)
C0474563|Hemoglobin; plasma
C0474563|Measurement of total hemoglobin concentration in plasma specimen
C0474563|Measurement of total haemoglobin concentration in plasma specimen
C0474563|Haemoglobin determination, plasma
C0474563|Hemoglobin determination, plasma (procedure)
C0474563|Measurement of total hemoglobin concentration in plasma specimen (procedure)
C0474563|Hemoglobin determination, plasma
C0474563|plasma hemoglobin measurement (lab test)
C0474563|plasma hemoglobin measurement
C0474563|Measurement of hemoglobin in plasma
C0474563|Plasma hemoglobin level
C0474563|ASSAY OF HEMOGLOBIN PLASMA
C0474563|Plasma Hemoglobins Test
C0474563|Plasma haemoglobin level
C0474563|Assay of plasma hemoglobin
C0373643|Hemoglobin; unstable, screen
C0373643|unstable hemoglobin screen
C0373643|unstable hemoglobin screen (lab test)
C0373643|HEMOGLOBIN UNSTABLE SCREEN
C0373643|Screening test for unstable hemoglobin
C0373643|Screening for unstable hemoglobin
C0373643|HEMOGLOBIN STABILITY SCREEN
C0373641|Hemoglobin; sulfhemoglobin, quantitative
C0373641|HEMOGLOBIN SULFHEMOGLOBIN QUANTITATIVE
C0373641|BLOOD SULFHEMOGLOBIN ASSAY
C3897698|Reticulocyte Mean Corpuscular Hemoglobin Measurement
C3897698|CHCMr
C3897698|Ret. Mean Corpuscular Hemoglobin
C3897698|RETIMCH
C3888302|HEMOGLOBIN S
C3888302|HEMOGLOBIN S PHENOTYPE
C3888302|HGBS
C3888302|Hemoglobin S Measurement
C3888302|Sickle Hemoglobin
C4066087|calculated hemoglobin level
C4066087|hemoglobin calculated
C4066087|calculated hemoglobin level (lab test)
C0200694|Measurement of total hemoglobin concentration and hematocrit (procedure)
C0200694|Hemoglobin and hematocrit determination
C0200694|Measurement of total hemoglobin concentration and hematocrit
C0200694|Measurement of total haemoglobin concentration and haematocrit
C0200694|Hemoglobin and hematocrit determination (procedure)
C0200694|Haemoglobin and haematocrit determination
C0200694|H & H determination
C0200694|total hemoglobin concentration and hematocrit
C0200694|total hemoglobin concentration and hematocrit (lab test)
C0200694|Haemoglobin and hematocrit determination
C0474755|Copper sulfate screening test
C0474755|Copper sulphate screening test
C0474755|Copper sulfate screening test (procedure)
C0523149|Semi-quantitative measurement of total haemoglobin in blood specimen
C0523149|Semi-quantitative measurement of total hemoglobin in blood specimen
C0523149|Haemoglobin determination, blood, semi-quantitative
C0523149|Semi-quantitative measurement of total hemoglobin in blood specimen (procedure)
C0523149|Hemoglobin determination, blood, semi-quantitative (procedure)
C0523149|Hemoglobin determination, blood, semi-quantitative
C0523151|Haemoglobin determination, urine
C0523151|Hemoglobin determination, urine (procedure)
C0523151|Measurement of total hemoglobin concentration in urine specimen (procedure)
C0523151|Measurement of total hemoglobin concentration in urine specimen
C0523151|Measurement of total haemoglobin concentration in urine specimen
C0523151|Hemoglobin determination, urine
C1314664|Haemoglobin concentration
C1314664|Dipstick assessment of hemoglobin concentration (procedure)
C1314664|Hemoglobin level
C1314664|Haemoglobin level
C1314664|Hb - Haemoglobin level
C1314664|Hb - Hemoglobin concentration
C1314664|Dipstick assessment of haemoglobin concentration
C1314664|Hb - Hemoglobin level
C1314664|Dipstick assessment of hemoglobin concentration
C1314664|Hb - Haemoglobin concentration
C1314664|Hemoglobin concentration
C0202054|Glycosylated Hemoglobin Measurement
C0202054|Glucohemoglobin measurement
C0202054|HBA1C
C0202054|Hemoglobin A1C
C0202054|Glycosylated Hemoglobin
C0202054|Glycated hemoglobin measurement
C0202054|Glycated haemoglobin measurement
C0202054|Glycosylated haemoglobin measurement
C0202054|Glucohaemoglobin measurement
C0202054|Glucohemoglobin measurement (procedure)
C0202054|Glucohemoglobin measurement, NOS
C0475357|Glycated haemoglobin-c fraction
C0475357|Glycated hemoglobin-c fraction
C0475357|Glycosylated haemoglobin-c fraction
C0475357|Glycosylated hemoglobin-c fraction
C0475357|HbA1c - Glycated haemoglobin-c fraction
C0475357|HbA1c - Glycated hemoglobin-c fraction
C0475357|HbA1c - Glycosylated haemoglobin-c fraction
C0475357|HbA1c - Glycosylated hemoglobin-c fraction
C0475357|Glycosylated hemoglobin-c fraction (substance)
C0018631|Hb A1a-2
C0019041|A1a-1 Hemoglobin, Glycosylated
C0019041|Glycosylated A1a-1 Hemoglobin
C0019041|Hemoglobin, Glycosylated A1a 1
C0019041|Hemoglobin, Glycosylated A1a-1
C0019041|Hb A1a-1
C2925136|Hemoglobin A1c &#x7C; Bld-Ser-Plas
C3181446|HbA(1c) protein, mouse
C0061430|glucosylated hemoglobin A
C0061430|hemoglobin A, glucosylated
C0019042|A1b Hemoglobin, Glycosylated
C0019042|Glycosylated A1b Hemoglobin
C0019042|Hemoglobin, Glycosylated A1b
C0019042|Hb A1b
C0071823|pre-hemoglobin A, glycosylated
C0209024|HBA(1c)-nitric oxide
C0209024|HbNO
C0209024|nitric oxide hemoglobin
C0209024|hemoglobin A, glycosylated-nitric oxide complex
C0296853|Hb A1d
C0296853|hemoglobin A1d
C1869903|hemoglobin A1c protein, human
C1869903|HbA1c protein, human
C1869903|blood HbA1c protein, human
C0585938|Hemoglobin A1 level
C0585938|Haemoglobin A1 level
C0585938|Haemoglobin A1 level (procedure)
C0585938|Haemoglobin A1 measurement
C0585938|Hemoglobin A1 measurement
C0585938|Hemoglobin A1 measurement (procedure)
C1295145|Glucose measurement estimated from glycated haemoglobin
C1295145|Glucose measurement estimated from glycated hemoglobin (procedure)
C1295145|Glucose measurement estimated from glycated hemoglobin
C0474680|Hemoglobin A1C level
C0474680|Haemoglobin A1c level
C0474680|Haemoglobin A1c level (procedure)
C0474680|Hemoglobin A1c Test
C0474680|Hemoglobin A1c measurement
C0474680|Haemoglobin A1c measurement
C0474680|HbA1c - Haemoglobin A1c level
C0474680|HbA1c - Hemoglobin A1c level
C0474680|Hemoglobin A1c measurement (procedure)
C1319284|Total glycosylated haemoglobin level (procedure)
C1319284|Total glycosylated hemoglobin level (procedure)
C1319284|Total glycosylated haemoglobin level
C1319284|Total glycosylated haemoglobin measurement
C1319284|Total glycosylated hemoglobin level
C1319284|Total glycosylated hemoglobin measurement
C1254681|Total Glycosylated Hemoglobins Test
C2012263|glycosylated hemoglobin A1C using home device
C2012263|hemoglobin A1C using home device
C2012263|hemoglobin A1C measurement using home device
C2012263|hemoglobin A1C measurement using home device (lab test)
C2012263|glycosylated hemoglobin A1C measurement using home device
C0239940|Glycosylated haemoglobin increased
C0239940|HbA1C increased
C0239940|Glycosylated hemoglobin increased
C0239940|Glycosylated haemoglobin high
C0239940|Glycohaemoglobin increased
C0239940|Glycohemoglobin increased
C0239940|Glycosylated hemoglobin high
C0239940|Hemoglobin A1C increased
C0239940|Haemoglobin A1C increased
C0239940|HgbA1c Increased
C0366781|Hemoglobin A1c/Hemoglobin.total in Blood
C0366781|Hgb A1c MFr Bld
C0366781|Hemoglobin A1c/Hemoglobin.total:MFr:Pt:Bld:Qn
C0366781|Hemoglobin A1c/Hemoglobin.total:Mass Fraction:Point in time:Whole blood:Quantitative
C0366782|Hemoglobin A1c/Hemoglobin.total in Blood by Electrophoresis
C0366782|Hgb A1c MFr Bld Elph
C0366782|Hemoglobin A1c/Hemoglobin.total:Mass Fraction:Point in time:Whole blood:Quantitative:Electrophoresis
C0366782|Hemoglobin A1c/Hemoglobin.total:MFr:Pt:Bld:Qn:Electrophoresis
C1255497|NYH Lab Procedure: Glycohgb A1c-Rogosin
C3838426|blood hemoglobin A1c/total ratio by calculation
C3838426|glycosylated hemoglobin a1c / total ratio by calculation
C3838426|blood hemoglobin A1c/total ratio by calculation (lab test)
C3838425|glycosylated hemoglobin a1c / total ratio by electrophoresis
C3838425|blood hemoglobin A1c/total ratio by electrophoresis (lab test)
C3838425|blood hemoglobin A1c/total ratio by electrophoresis
C3838424|glycosylated hemoglobin a1c / total ratio by hplc
C3838424|blood hemoglobin A1c/total ratio by HPLC
C3838424|blood hemoglobin A1c/total ratio by HPLC (lab test)
C3838427|blood hemoglobin A1c/total ratio
C3838427|blood hemoglobin A1c/total ratio (lab test)
C3838427|glycosylated hemoglobin a1c / total ratio
C1277712|Hemoglobin A1c measurement aligned to the Diabetes Control and Complications Trial (procedure)
C1277712|HbA1c measurement (DCCT aligned) (procedure)
C1277712|Hemoglobin A1c measurement aligned to the Diabetes Control and Complications Trial
C1277712|HbA1c level (DCCT aligned) (procedure)
C1277712|HbA1c level (DCCT aligned)
C1277712|HbA1c measurement (DCCT aligned)
C0800962|Hemoglobin A1c/Hemoglobin.total in Blood by calculation
C0800962|Hemoglobin A1c/Hemoglobin.total:MFr:Pt:Bld:Qn:Calculated
C0800962|Hgb A1c MFr Bld Calc
C0800962|Hemoglobin A1c/Hemoglobin.total:Mass Fraction:Point in time:Whole blood:Quantitative:Calculated
C0800963|Hemoglobin A1c/Hemoglobin.total in Blood by HPLC
C0800963|Hemoglobin A1c/Hemoglobin.total:MFr:Pt:Bld:Qn:HPLC
C0800963|Hemoglobin A1c/Hemoglobin.total:Mass Fraction:Point in time:Whole blood:Quantitative:HPLC
C0800963|Hgb A1c MFr Bld HPLC
C2960128|Hemoglobin A1c target value using International Federation of Clinical Chemistry and Laboratory Medicine standardized method (observable entity)
C2960128|Haemoglobin A1c target value using International Federation of Clinical Chemistry and Laboratory Medicine standardised method
C2960128|Hemoglobin A1c target value using International Federation of Clinical Chemistry and Laboratory Medicine standardized method
C2707530|Hemoglobin A1c in Blood
C2707530|Hgb A1c Bld
C2707530|Hemoglobin A1c:-:Pt:Bld:-
C2707530|Hemoglobin A1c:-:Point in time:Whole blood:-
C2923665|Hgb A1c SFr Bld IFCC
C2923665|Hemoglobin A1c/Hemoglobin.total in Blood by IFCC protocol
C2923665|Hemoglobin A1c/Hemoglobin.total:SFr:Pt:Bld:Qn:IFCC
C2923665|Hemoglobin A1c/Hemoglobin.total:Substance Fraction:Point in time:Whole blood:Quantitative:IFCC
C2973266|Hemoglobin A1c/Hemoglobin.total:Mass Fraction:Point in time:Whole blood:Quantitative:JDS/JSCC
C2973266|Hemoglobin A1c/Hemoglobin.total:MFr:Pt:Bld:Qn:JDS/JSCC
C2973266|Hemoglobin A1c/Hemoglobin.total in Blood by JDS/JSCC protocol
C2973266|Hgb A1c MFr Bld JDS/JSCC
C3484089|Hemoglobin A1c/Hemoglobin.total:Mass decimal fraction:Point in time:Whole blood:Quantitative
C3484089|Hemoglobin A1c/Hemoglobin.total:MFr.DF:Pt:Bld:Qn
C3484089|Hemoglobin A1c/Hemoglobin.total [Pure mass fraction] in Blood
C3484089|Hgb A1c MFr.DF Bld
C0438275|Hb. A1C - diabetic control NOS
C0438275|Hb. A1C - diabetic control NOS (observable entity)
C0438275|Hb. A1C - diabetic control NOS (procedure)
C0587827|HbA1 - diabetic control interpretation
C0587827|HbA1 - diabetic control interpretation (observable entity)
C0587827|HbA1 - diabetic control
C0587827|HbA1 - diabetic control (observable entity)
C2919483|High hemoglobin A1c level
C2919483|Haemoglobin A1c above reference range
C2919483|High haemoglobin A1c level
C2919483|Hemoglobin A1c above reference range
C2919483|Hemoglobin A1c above reference range (finding)
C1287394|HbA1 - diabetic control finding
C1287394|HbA1 - diabetic control finding (finding)
C1287394|Haemoglobin A1C - diabetic control finding
C1287394|Hemoglobin A1C - diabetic control finding (finding)
C1287394|Hemoglobin A1C - diabetic control finding
C0587829|HbA1 7-10% - borderline control (finding)
C0587829|HbA1 7-10% - borderline control
C0587830|HbA1 greater than 10% - bad control
C0587830|HbA1 greater than 10% - bad control (finding)
C0587828|HbA1 less than 7% - good control (finding)
C0587828|HbA1 less than 7% - good control
C0438277|HbA1C 7-10% - borderline (finding)
C0438277|Hemoglobin A1c between 7%-10% indicating borderline diabetic control (finding)
C0438277|Hb. A1C 7-10% - borderline
C0438277|Hemoglobin A1c (HbA1c) between 7%-10% indicating borderline diabetic control
C0438277|Hemoglobin A1c between 7%-10% indicating borderline diabetic control
C0438277|Haemoglobin A1c (HbA1c) between 7%-10% indicating borderline diabetic control
C0438277|Haemoglobin A1c between 7%-10% indicating borderline diabetic control
C0438277|Hb. A1C 7-10% - borderline (finding)
C0438276|Hemoglobin A1c less than 7% indicating good diabetic control
C0438276|Hb. A1C < 7% - good control
C0438276|Hemoglobin A1c less than 7% indicating good diabetic control (finding)
C0438276|Hemoglobin A1c (HbA1c) less than 7% indicating good diabetic control
C0438276|HbA1C < 7% - good control (finding)
C0438276|Haemoglobin A1c less than 7% indicating good diabetic control
C0438276|Haemoglobin A1c (HbA1c) less than 7% indicating good diabetic control
C0438276|Hb. A1C < 7% - good control (finding)
C0438278|Hemoglobin A1c greater than 10% indicating poor diabetic control (finding)
C0438278|Haemoglobin A1c (HbA1c) greater than 10% indicating poor diabetic control
C0438278|Hb. A1C > 10% - bad control
C0438278|Hemoglobin A1c greater than 10% indicating poor diabetic control
C0438278|Haemoglobin A1c greater than 10% indicating poor diabetic control
C0438278|Hemoglobin A1c (HbA1c) greater than 10% indicating poor diabetic control
C0438278|HbA1C > 10% - bad control (finding)
C0438278|Hb. A1C > 10% - bad control (finding)
C1624104|Hemoglobin A1c:MCnc:Pt:Bld:Qn
C1624104|Hemoglobin A1c [Mass/volume] in Blood
C1624104|Hgb A1c Bld-mCnc
C1624104|Hemoglobin A1c:Mass Concentration:Point in time:Whole blood:Quantitative
C1624124|HbA1c measurement device panel:-:Pt:^Patient:-
C1624124|Hemoglobin A1c measurement device panel
C1624124|Hb A1c Measurement Device Pnl
C1624124|HbA1c measurement device panel:-:Point in time:^Patient:-
C1650487|Vendor device name:ID:Pt:HbA1c measurement device:Nom
C1650487|HbA1c measurement device Vendor name
C1650487|Vendor device name:Identifier:Point in time:HbA1c measurement device:Nominal
C1650488|Vendor serial number:ID:Pt:HbA1c measurement device:Nom
C1650488|HbA1c measurement device Vendor serial number
C1650488|HbA1c Measurement Device Serial #
C1650488|Vendor serial number:Identifier:Point in time:HbA1c measurement device:Nominal
C1652140|HbA1c Measurement Device Model Cd
C1652140|Vendor device model code:ID:Pt:HbA1c measurement device:Nom
C1652140|HbA1c measurement device Vendor model code
C1652140|Vendor device model code:Identifier:Point in time:HbA1c measurement device:Nominal
C1652141|HbA1c measurement device Vendor software version
C1652141|Vendor software version:ID:Pt:HbA1c measurement device:Nom
C1652141|HbA1c Measurement Device Software vers
C1652141|Vendor software version:Identifier:Point in time:HbA1c measurement device:Nominal
C1633474|Class:Type:Pt:HbA1c measurement device:Nom
C1633474|Type of HbA1c measurement device
C1633474|HbA1c Measurement Device Class
C1633474|Class:Type:Point in time:HbA1c measurement device:Nominal
C2114374|hemoglobin A1C level > 9.0%
C2114374|hemoglobin A1C level greater 9.0%
C2114374|hemoglobin A1C level greater 9.0% (treatment)
C2114374|hemoglobin A1C results documented and reviewed - hemoglobin A1C level greater 9.0%
C2114346|hemoglobin A1C level < 7.0%
C2114346|hemoglobin A1C level less than 7.0%
C2114346|hemoglobin A1C level less than 7.0% (treatment)
C2114347|hemoglobin A1C level 7.0-9.0% (treatment)
C2114347|hemoglobin A1C level 7.0-9.0%
C1737720|Most recent hemoglobin A1c level > 9.0% (DM)
C1737720|Most recent hemoglobin A1c level greater than 9.0% (DM)
C1737720|MOST RECENT HEMOGLOBIN A1C LEVEL >9.0%
C1737720|HEMOGLOBIN A1C LEVEL >9.0%
C1964112|HG A1C LEVEL LT 7.0%
C1964112|Most recent hemoglobin A1c (HbA1c) level less than 7.0% (DM)
C1964112|MOST RECENT HEMOGLOBIN A1C LEVEL < 7.0%
C1277717|HbA1 measurement (DCCT aligned) (procedure)
C1277717|HbA1 measurement (DCCT aligned)
C1277717|Haemoglobin A1 measurement (Diabetes Control and Complications Trial aligned)
C1277717|Hemoglobin A1 measurement (Diabetes Control and Complications Trial aligned) (procedure)
C1277717|HbA1 level (DCCT aligned) (procedure)
C1277717|HbA1 level (DCCT aligned)
C1277717|Hemoglobin A1 measurement (Diabetes Control and Complications Trial aligned)
C1964113|HG A1C LEVEL 7.0-9.0%
C1964113|Most recent hemoglobin A1c (HbA1c) level 7.0-9.0% (DM)
C1964113|MOST RECENT HEMOGLOBIN A1C LEVEL GT 7.0-9.0 %
