C0019683|HIV Ab
C0019683|HIV Antibodies
C3714540|HIV Antibody Test
C3714540|HIV Antibody Measurement
C0019683|Antibodies, AIDS
C0019683|Antibodies, HIV
C0019683|Antibodies, HIV Associated
C0019683|Antibodies, HIV-Associated
C0019683|Antibodies, HTLV III
C0019683|Antibodies, HTLV-III
C0019683|Antibodies, HTLV-III-LAV
C0019683|Antibodies, LAV
C0019683|Antibodies, Lymphadenopathy Associated
C0019683|Antibodies, Lymphadenopathy-Associated
C0019683|HIV Antibodies
C0019683|HTLV WIII ANTIBODIES
C0019683|HTLV WIII LAV ANTIBODIES
C0019683|LYMPHOTROPIC VIRUS TYPE III ANTIBODIES HUMAN T
C0019683|HTLV-III Antibodies
C0019683|HIV Antibodies [Chemical/Ingredient]
C0019683|HTLV III Antibodies
C0019683|LAV Antibodies
C0019683|Lymphadenopathy Associated Antibodies
C0019683|T Lymphotropic Virus Type III Antibodies, Human
C0019683|AIDS Antibodies
C0019683|HIV Associated Antibodies
C0019683|T-Lymphotropic Virus Type III Antibodies, Human
C0019683|HIV-Associated Antibodies
C0019683|HTLV-III-LAV Antibodies
C0019683|HTLV III LAV Antibodies
C0019683|Lymphadenopathy-Associated Antibodies
C0019683|HIV antibody
C0019683|HIV - Human immunodeficiency virus antibody
C0019683|Human immunodeficiency virus antibody
C0019683|Human immunodeficiency virus antibody (substance)
C0019683|ARV Antibody
C0019683|HTLV-III Antibody
C0474652|Human immunodeficiency virus antibody titer measurement
C0474652|Human immunodeficiency virus antibody level (substance)
C0474652|Human immunodeficiency virus antibody level
C0474652|Human immunodeficiency virus antibody level (procedure)
C0474652|HIV - Human immunodeficiency virus antibody titer
C0474652|HIV - Human immunodeficiency virus antibody titre
C0474652|Human immunodeficiency virus antibody titer
C0474652|Human immunodeficiency virus antibody titre
C0474652|Human immunodeficiency virus antibody titer measurement (procedure)
C0474652|Human immunodeficiency virus antibody titre measurement
C0474652|Human immunodeficiency virus antibody assay
C3181597|4E10 MAb
C3181597|MAb 4E10
C3181597|4E10 monoclonal antibody
C4043370|3BNC117 antibody
C0369497|Human immunodeficiency virus, type I antibody
C0369497|Human immunodeficiency virus type 1 antibody
C0369497|HIV 1 Ab
C0369497|human immunodeficiency virus 1 Antibody
C0369497|Human immunodeficiency virus, type I antibody (substance)
C0369497|HIV-1 Antibody
C0369497|Human immunodeficiency virus type 1 antibody (substance)
C0369497|LAV-1 Antibody
C0369500|Human immunodeficiency virus type 2 (HIV-2) antibody
C0369500|HIV 2 Ab
C0369500|human immunodeficiency virus 2 Antibody
C0369500|Human immunodeficiency virus type 2 antibody
C0369500|Human immunodeficiency virus, type II antibody (substance)
C0369500|Human immunodeficiency virus, type II antibody
C3179325|PRO-140 monoclonal antibody
C3714540|HIV antibody
C3714540|HIV Antibody Measurement
C3714540|HIVAB
