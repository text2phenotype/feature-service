C1515945|American Indian or Alaska Native
C3261247|American indian and alaska native alone
C0078988|Asians
C0078988|Asian
C0003988|Asian Americans
C0003988|Asian American
C0438971|Other Asian ethnic group
C1524069|Asian Indian
C3261249|Asian alone
C0085756|African American
C0005680|Black race
C0027567|African race
C0085756|African American
C0085756|African
C0085756|Botswanan
C0085756|Ethiopian
C0085756|Liberian
C0085756|Namibian
C0085756|Nigerian
C0085756|Zairean
C0085756|Bahamian
C0085756|Barbadian
C0085756|Dominica Islander
C0085756|Dominican
C0085756|Haitian
C0085756|Jamaican
C0085756|Tobagoan
C0085756|Trinidadian
C0085756|West Indian
C1513907|Native Hawaiian or Other Pacific Islander
C1513907|Melanesian
C1513907|Fijian
C1513907|New Hebrides
C1513907|Papua New Guinean
C1513907|Solomon Islander
C1513907|Micronesian
C1513907|Carolinian
C1513907|Chamorro
C1513907|Chuukese
C1513907|Guamanian or Chamorro
C1513907|Guamanian
C1513907|Kiribati
C1513907|Kosraean
C1513907|Mariana Islander
C1513907|Marshallese
C1513907|Palauan
C1513907|Pohnpeian
C1513907|Saipanese
C1513907|Yapese
C1513907|Other Pacific Islander
C1513907|Polynesian
C1513907|Native Hawaiian
C1513907|Samoan
C1513907|Tahitian
C1513907|Tokelauan
C1513907|Tongan
C0043157|Caucasians
C0043157|European
C0043157|Armenian
C0043157|English
C0043157|French
C0043157|German
C0043157|Irish
C0043157|Italian
C0043157|Polish
C0043157|Scottish
C0221786|white American
C1535514|European race
C0086409|Hispanics
C0086409|Central American
C0086409|Canal Zone
C0086409|Central American Indian
C0086409|Costa Rican
C0086409|Guatemalan
C0086409|Honduran
C0086409|Nicaraguan
C0086409|Panamanian
C0086409|Salvadoran
C0086409|Cuban
C0086409|Dominican
C0086409|Latin American
C0086409|Mexican
C0086409|Chicano
C0086409|La Raza
C0086409|Mexican American Indian
C0086409|Mexican American
C0086409|Mexicano
C0086409|Puerto Rican
C0086409|South American
C0086409|Argentinean
C0086409|Bolivian
C0086409|Chilean
C0086409|Colombian
C0086409|Criollo
C0086409|Ecuadorian
C0086409|Paraguayan
C0086409|Peruvian
C0086409|South American Indian
C0086409|Uruguayan
C0086409|Venezuelan
C0086409|Spaniard
C0086409|Andalusian
C0086409|Asturian
C0086409|Belearic Islander
C0086409|Canarian
C0086409|Castillian
C0086409|Catalonian
C0086409|Gallego
C0086409|Spanish Basque
C0086409|Valencian
C3846650|Spanish,NOS; Hispanic,NOS
C0019576|Hispanic Americans
C1533017|Hispanic black finding
C1533018|Hispanic black racial group
C1533020|Hispanic white finding
C1533021|Hispanic white racial group
C1881927|Multiple Hispanic
C2741637|Hispanic or Latino:Finding:Point in time:^Patient:Ordina
C3844642|Other Hispanic
C4036190|Yes, another Hispanic, Latino-a, or Spanish origin
C3161701|cultural background alaskan native (___ %) (history)
C3161701|cultural background alaskan native (___ %)
C0002460|American Indian
C0002460|American Indians
C0002460|Indian, American
C0002460|Indians, American
C0002460|RaceAmericanIndian
C0002460|American Indian race (finding)
C0002460|American Indian race
C0002460|Amerindian race
C0002460|Amerindian
C0002460|Indians (American)
C0002460|American Indian race (racial group)
C0682125|Alaska Indian
C0682125|RaceAlaskanNative
C0682125|RaceAlaskanIndian
C0682125|Alaska Native
C0682125|Alaska Natives
C0682125|Native Alaskans
C0682125|Alaska Indians
C0152035|Chinese
C0152035|Chinese People
C0152035|Chinese (ethnic group)
C0152035|-- Chinese
C1556094|Japanese
C1556094|Race: Japanese (finding)
C1556094|Race: Japanese
C1556094|-- Japanese
C1556094|Japanese (ethnic group)
C1556094|Japanese race
C0238697|southeast Asian
C0238697|South East Asian
C0238697|South East Asian (ethnic group)
C0596476|East Indian
C1556093|Filipino
C1556093|-- Filipino
C1556093|Filipinos
C1556093|Filipinos (ethnic group)
C1556093|Filipino race
C0078988|Asian
C0078988|Asians
C0078988|oriental
C0078988|RaceAsian
C0078988|Asian race
C0078988|Race: Oriental (finding)
C0078988|Asian race (finding)
C0078988|Race: Oriental
C0078988|Oriental (ethnic group)
C0078988|Asian race (racial group)
C0438971|Other Asian ethnic group
C0438971|Other Asian (ethnic group)
C0438971|Other Asian ethnic group (ethnic group)
C0438971|Other Asian
C0438971|-- Other Asian
C0870279|Chinese Cultural Groups
C0870754|Japanese Cultural Groups
C0870776|Korean Cultural Groups
C0871579|Vietnamese Cultural Groups
C1510645|South Asian Cultural Groups
C1510577|Southeast Asian Cultural Groups
C1553332|Malagasy
C1553332|Madagascar
C1553332|Madagascar race
C1553322|Burmese
C1553322|Burmeses
C0337900|Indonesian
C0337900|Indonesians
C0337900|Indonesians (ethnic group)
C1556095|Korean
C1556095|Race: Korean
C1556095|Race: Korean (finding)
C1556095|-- Korean
C1556095|Koreans
C1556095|Koreans (ethnic group)
C1556095|Korean race
C0337910|Thai
C0337910|Thaus
C0337910|Thais (Population Group)
C0337910|Thais
C0337910|Thais (ethnic group)
C1561452|Vietnamese
C1561452|Vietnameses
C1561452|Vietnamese (ethnic group)
C1561452|-- Vietnamese
C1561452|Vietnamese race
C1553323|Cambodian
C1553323|Kampuchean
C1553323|Cambodians
C0337894|Bhutanese
C0337894|Bhutanese (ethnic group)
C1556096|Taiwanese
C1556096|Taiwanese (ethnic group)
C1556096|Race - Taiwanese
C1556107|Bangladeshi
C1556107|Bangladeshi race
C0425375|Pakistani
C0425375|Race: Pakistani
C0425375|Race: Pakistani (finding)
C0425375|Pakistani race
C0240293|Malaysian
C0240293|Malaysian race
C1524069|Indian
C1524069|Indian (East Indian)
C1524069|Indian (ethnic group)
C1524069|Indian race (finding)
C1524069|Indian sub-continent (NMO)
C1524069|Indian race
C1524069|Indian sub-continent (NMO) (ethnic group)
C1524069|Asian Indian
C1524069|-- Asian Indian
C1524069|Indian (East Indian) (ethnic group)
C1524069|Asian Indians
C1524069|Indian (racial group)
C1553324|Hmong
C1553328|Iwo Jiman
C1553328|Iwo Jiman race
C1553325|Laotian
C1553325|Laotian race
C1553329|Maldivian
C1553329|Maldivian race
C1553330|Nepalese
C1553330|Nepalese race
C1553326|Okinawan
C1553326|Okinawan race
C1553331|Singaporean
C1553331|Singaporean race
C1553327|Sri Lankan
C1553327|Sri Lankan race
C0337893|Ainu
C0337893|Ainu (ethnic group)
C0337892|Mongoloid population
C0337892|Mongol (ethnic group)
C0337892|Mongoloid
C0337892|Mongoloid (ethnic group)
C0337892|Mongol
C0337892|Mongoloid race
C0337892|Asiatic Race
C0337892|Asiatic Races
C0337892|Mongoloid Races
C0337892|Race, Asiatic
C0337892|Race, Mongoloid
C0337892|Races, Asiatic
C0337892|Races, Mongoloid
C0337892|Mongoloid, NOS
C0337920|Hawaiian
C0337920|Hawaiian population
C0337920|Native Hawaiian
C0337920|-- Native Hawaiian
C0337920|Hawaiian, Native
C0337920|Hawaiians, Native
C0337920|Native Hawaiians
C0337920|Hawaiians
C0337920|Hawaiians (ethnic group)
C0337920|Hawaii Natives
C1519427|South Asians
C1519427|South Asian
C1709065|Mongolian
C1709065|Mongolian (race)
C0008121|American, Chinese
C0008121|Americans, Chinese
C0008121|Chinese American
C0008121|Chinese Americans
C0022343|American, Japanese
C0022343|Americans, Japanese
C0022343|Japanese American
C0022343|Japanese Americans
C0597918|Filipino American
C0597919|Indochinese American
C0597920|Indonesian American
C0597921|Korean American
C0597921|Americans, Korean
C0597921|American, Korean
C0597921|Korean Americans
C0003988|American, Asian
C0003988|Americans, Asian
C0003988|Asian American
C0003988|Asian Americans
C0003988|Asian-American
C0085756|African American
C0085756|Americans, African
C0085756|Afroamerican
C0085756|black American
C0085756|United States Black
C0085756|U.S. Blacks
C0085756|RaceBlackOrAfricanAmerican
C0085756|African Americans
C0085756|Black
C0085756|BLACK OR AFRICAN AMERICAN
C0085756|Black or African-American
C0085756|African-American
C0085756|Black/African American
C0085756|African American (ethnic group)
C0085756|Black Populations
C0085756|Afro American
C0005680|Black race
C0005680|Blacks
C0005680|Negroes
C0005680|Negro
C0005680|Black
C0005680|Black - ethnic group (ethnic group)
C0005680|Black - ethnic group
C0027567|African
C0027567|African race (finding)
C0027567|African race
C0027567|Negroid
C0027567|Negroid Race
C0027567|Negroid Races
C0027567|Race, Negroid
C0027567|Races, Negroid
C0027567|Black
C0027567|African race (racial group)
C1553338|Dominican
C1553338|Dominica Islander
C1553338|Dominica Islander race
C0239806|Haitian
C0239806|Haitian race
C0240072|Jamaican
C1553339|Tobagoan
C1553339|Tobagoan race
C1553340|Trinidadian
C1553340|Trinidadian race
C0425373|West Indian
C0425373|Race: West indian
C0425373|Race: West indian (ethnic group)
C0425373|Race: West indian (finding)
C0425373|West Indian race
C1553336|Bahamian
C1553336|Bahamian race
C1553337|Barbadian
C1553337|Barbadian race
C2135340|cultural background African American (history)
C2135340|cultural background African American
C2135340|the cultural background is African American
C2135340|Social history - cultural background African American
C0422781|Black - other, mixed
C0422781|Black - other, mixed (ethnic group)
C0337824|Black African (ethnic group)
C0337824|Black African
C0337824|Black African, NOS
C0422771|African Caribbean
C0422771|black carib
C0422771|black Caribbean
C0422771|Black Caribbean (ethnic group)
C0422772|Black, other, non-mixed origin
C0422772|Black, other, non-mixed origin (ethnic group)
C1278528|Other black ethnic group
C1278528|Other black ethnic group (ethnic group)
C2135370|racial background black (history)
C2135370|racial background Black
C1531522|Black, not of hispanic origin (racial group)
C1531522|Black, not of hispanic origin
C0239304|Ethiopian
C1556088|Liberian
C1556088|Liberians
C1556088|Liberians (ethnic group)
C1556088|Liberian race
C1553334|Namibian
C1553334|Namibian race
C1556089|Nigerian
C1556089|Nigerians
C1556089|Nigerians (ethnic group)
C1556089|Nigerian race
C1553335|Zairean
C1553335|Zairean race
C1553333|Botswanan
C1553333|Motswana
C1553333|Botswanan race
C1553351|Other Pacific Islander
C1553351|-- Other Pacific Islander
C0337924|Melanesian
C0337924|RacePacificIslandMelanesian
C0337924|Melanesian, NOS
C0337924|Melanesians
C0337924|Melanesians (ethnic group)
C0337924|Melanesian-Papuan
C0337924|Melanesian (ethnic group)
C0240790|Polynesian
C0240790|RacePacificIslandPolynesian
C0240790|Polynesian race (finding)
C0240790|Polynesian race
C0240790|Polynesian, NOS
C0240790|Polynesians
C0240790|Polynesians (ethnic group)
C1556099|Micronesian
C1556099|RacePacificIslandMicronesian
C1556099|Micronesian race (finding)
C1556099|Micronesian race
C1556099|Micronesian, NOS
C1556099|Micronesians
C1556099|Micronesians (ethnic group)
C0221786|caucasian American
C0221786|white American
C0337815|Poles
C0337815|Poles (ethnic group)
C0337799|Czechs
C0337799|Czechs (ethnic group)
C1556085|German
C1556085|Germans
C1556085|Germans (ethnic group)
C1556085|german race
C0337800|Danes
C0337800|Danes (ethnic group)
C0337796|Basques
C0337796|Basques (ethnic group)
C0337806|Greek
C0337806|Greeks
C0337806|Greeks (ethnic group)
C1556083|English
C1556083|English (ethnic group)
C1556083|English race
C0337795|Austrians
C0337795|Austrians (ethnic group)
C1556087|Iraqi
C1556087|Iraqi (ethnic group)
C1556087|Iraqi race
C0337811|Irani
C0337811|Irani (ethnic group)
C0337817|Spaniards
C0337817|Spaniards (ethnic group)
C0337817|Spaniard
C0337797|Belgians
C0337797|Belgians (ethnic group)
C0337801|Egyptian
C0337801|Egyptians
C0337801|Egyptians (ethnic group)
C0032730|Portuguese population
C0032730|Portuguese
C0032730|Portuguese (ethnic group)
C0337802|Estonians
C0337802|Estonians (ethnic group)
C0013331|Dutch Population
C0013331|Dutch
C0013331|Dutch (ethnic group)
C0337809|Indians (Hindi-speaking)
C0337809|Indians (Hindi-speaking) (ethnic group)
C0337798|Bulgarians
C0337798|Bulgarians (ethnic group)
C0337821|Serbs
C0337821|Serbs (ethnic group)
C0241315|Swiss
C0241315|Swiss (ethnic group)
C0337816|Russian
C0337816|Russians
C0337816|Russians (ethnic group)
C1556084|French
C1556084|French (ethnic group)
C1556084|french race
C0337804|Georgians
C0337804|Georgians (ethnic group)
C0337820|Tristan da Cunhans
C0337820|Tristan da Cunhans (ethnic group)
C0337818|Swedes
C0337818|Swedes (ethnic group)
C0337808|Icelanders
C0337808|Icelanders (ethnic group)
C0337819|Syrian
C0337819|Syrians (ethnic group)
C0337819|Syrians
C0337822|Slovaks
C0337822|Slovaks (ethnic group)
C0337812|Norwegian
C0337812|Norwegians
C0337812|Norwegians (ethnic group)
C0043114|Welsh population
C0043114|Welsh
C0043114|Welsh (ethnic group)
C0337803|Finns
C0337803|Finns (ethnic group)
C1278525|Other white ethnic group (ethnic group)
C1278525|Other white ethnic group
C0043157|Caucasians
C0043157|caucasian
C0043157|RaceWhite
C0043157|Caucasian (living organism) (ethnic group)
C0043157|White - ethnic group (ethnic group)
C0043157|White - ethnic group
C0043157|White
C0043157|White/Caucasian
C0043157|Whites
C0043157|Caucasoid
C0043157|Caucasian (ethnic group)
C0043157|Caucasian, NOS
C0043157|Caucasian (living organism)
C1278523|White British (ethnic group)
C1278523|White British
C1278524|White Irish (ethnic group)
C1278524|White Irish
C0870136|Anglos
C0007457|Caucasoid Race
C0007457|white race
C0007457|racial background Caucasian
C0007457|racial background Caucasian (history)
C0007457|Race: Caucasian
C0007457|Caucasian race
C0007457|Race: Caucasian (racial group)
C0007457|Race: Caucasian (finding)
C0007457|Race: White
C0007457|Caucasoid
C0007457|WHITE
C0007457|Caucasian Races
C0007457|Caucasoid Races
C0007457|Race, Caucasian
C0007457|Race, Caucasoid
C0007457|Races, Caucasian
C0007457|Races, Caucasoid
C0007457|Caucasian
C0007457|Whites
C0007457|Caucasians
C0007457|Occidental
C0007457|Caucasian (racial group)
C0239307|European
C0239307|European (ethnic group)
C0239307|ethnic european
C0337794|Armenian
C0337794|Armenians
C0337794|Armenians (ethnic group)
C0087186|Irish
C0087186|Irish race
C0337810|Italian
C0337810|Italians
C0337810|Italians (ethnic group)
C0220896|Polish population
C0220896|Polish
C0240966|Scottish
C0240966|Scottish race
C1710263|Swedish
C1710525|Ukranian
C1711254|Finnish
C0019576|American, Hispanic
C0019576|Americans, Hispanic
C0019576|Americans, Spanish
C0019576|Hispanic American
C0019576|Hispanic Americans
C0019576|Spanish American
C0019576|Spanish Americans
C1553379|Cuban
C1553379|-- Cuban
C3829110|Mexican or Mexican American
C3828691|Other Hispanic or Latino(a)
C3161473|Spanish
C3161473|Spanish Person
C0086409|Hispanic
C0086409|Hispanics
C0086409|Hispanic or Latino
C0086409|EthnicityHispanic
C0086409|Hispanic origin
C0086409|Spanish
C0086409|Hispanic Populations
C0086409|Hispanics or Latinos
C0086409|Latino Population
C0086409|Spanish Origin
C0086409|Hispanic (racial group)
C0025884|American, Mexican
C0025884|Americans, Mexican
C0025884|Chicano
C0025884|Mexican American
C0025884|Mexican Americans
C0025884|Chicanos
C0025884|Chicanas
C0025884|Chicana
C0010436|Americans, Cuban
C0010436|Cuban American
C0010436|Cuban Americans
C0086528|Latino
C0086528|Latinos
C0034043|Puerto Rican
C0034043|Puertorican
C0034043|-- Puerto Rican
C0034043|Puerto Ricans
C0935556|Latinos/Latinas
C1533018|Hispanic, black (racial group)
C1533018|Hispanic, black
C1533018|Hispanic black racial group
C1533019|Hispanic, color unknown (racial group)
C1533019|Hispanic, color unknown
C1533019|Hispanic, colour unknown
C1533021|Hispanic, white (racial group)
C1533021|Hispanic, white
C1533021|Hispanic white racial group
C0425359|South American
C0425359|-- South American
C0240339|Mexican
C0240339|EthnicityHispanicMexican
C0240339|-- Mexican
C0238914|Central American
C0238914|EthnicityHispanicCentralAmerican
C0238914|-- Central American
C1328872|Dominican
C1328872|Dominican - Ethnicity
C1553378|Latin American
C1881927|Multiple Hispanic
C1880193|Cuban or Cuban American
C2135343|cultural background Hispanic (history)
C2135343|the cultural background is Hispanic
C2135343|cultural background Hispanic
C2741637|Hispanic or Latino:Finding:Point in time:^Patient:Ordinal
C2741637|Hispanic or Latino
C2741637|Hispanic or Latino:Find:Pt:^Patient:Ord
