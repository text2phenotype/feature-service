C0551008|Hepatitis C Quantitation
C0551008|Hepatitis C RNA
C0551008|HCV log10
C0551008|HCV RNA
C0551008|Hepatitis C virus RNA
C0551008|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C0551008|LOINC 11011-4
C0551008|LOINC 38180-6
C1273338|Hepatitis C viral load
C1868902|HCV viral load
C2697584|Hepatitis C Viral Load PCR Measurement
C0485398|Hepatitis C virus RNA
C0485398|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp
C0551008|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C0803231|Hepatitis C virus RNA:NCnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C0803380|Hepatitis C virus RNA:NCnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C0945037|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C1508112|Hepatitis C virus RNA:LaCnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C1623573|Hepatitis C virus RNA:LnCnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C1643191|Hepatitis C virus RNA:LaCnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C1831320|Hepatitis C virus RNA:LnCnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C1977155|Hepatitis C virus RNA:NCnc:Pt:CSF:Qn:Probe.amp.tar
C1977156|Hepatitis C virus RNA:NCnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977157|Hepatitis C virus RNA:NCnc:Pt:Tiss:Qn:Probe.amp.tar
C1977158|Hepatitis C virus RNA:LnCnc:Pt:XXX:Qn:Probe.amp.tar
C1977159|Hepatitis C virus RNA:LnCnc:Pt:CSF:Qn:Probe.amp.tar
C1977160|Hepatitis C virus RNA:LnCnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977161|Hepatitis C virus RNA:LnCnc:Pt:Tiss:Qn:Probe.amp.tar
C1977162|Hepatitis C virus RNA:ACnc:Pt:XXX:Qn:Probe.amp.tar
C1977163|Hepatitis C virus RNA:ACnc:Pt:CSF:Qn:Probe.amp.tar
C1977164|Hepatitis C virus RNA:ACnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977165|Hepatitis C virus RNA:ACnc:Pt:Tiss:Qn:Probe.amp.tar
C1977166|Hepatitis C virus RNA:NCnc:Pt:XXX:Qn:Probe.amp.tar
C1977368|Hepatitis C virus RNA:LaCnc:Pt:CSF:Qn:Probe.amp.tar
C1977369|Hepatitis C virus RNA:LaCnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977370|Hepatitis C virus RNA:LaCnc:Pt:XXX:Qn:Probe.amp.tar
C1977373|Hepatitis C virus RNA:LaCnc:Pt:Tiss:Qn:Probe.amp.tar
C1977893|Hepatitis C virus RNA panel:-:Pt:Ser/Plas:Qn:Probe.amp.tar
C4064960|hepatitis C virus RNA viral load in serum or plasma by probe and target amplification
C1369569|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar detection limit = 500 IU/mL
C1369570|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar detection limit = 50 IU/mL
C1977509|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar detection limit = 5 IU/mL
C0551008|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C0551008|HCV RNA SerPl PCR-aCnc
C0551008|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar
C0551008|Hepatitis C virus RNA [Units/volume] (viral load) in Serum or Plasma by Probe and target amplification method
C1273338|Hepatitis C viral load
C1273338|Hepatitis C viral load (procedure)
C4064960|probe & target amplif hepatitis c virus rna serum/plasma viral load
C4064960|hepatitis C virus RNA viral load in serum or plasma by probe with target amplification (lab test)
C4064960|hepatitis C virus RNA viral load in serum or plasma by probe with target amplification
C1868902|Hepatitis C Viral Load Measurement
C1868902|HCV RNA
C1868902|Hepatitis C RNA
C1868902|HCV Viral Load
C1868902|HCVVLD
C0485398|Hepatitis C virus RNA [Units/volume] (viral load) in Serum or Plasma by Probe with amplification
C0485398|HCV RNA SerPl Amp Prb-aCnc
C0485398|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp
C0485398|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp
C0803231|HCV RNA # SerPl PCR
C0803231|Hepatitis C virus RNA:NCnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C0803231|Hepatitis C virus ribonucleic acid:Number Concentration (count/vol):Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar
C0803231|Hepatitis C virus RNA [#/volume] (viral load) in Serum or Plasma by Probe and target amplification method
C0803380|HCV RNA # SerPl bDNA
C0803380|Hepatitis C virus RNA:NCnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C0803380|Hepatitis C virus ribonucleic acid:Number Concentration (count/vol):Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.sig
C0803380|Hepatitis C virus RNA [#/volume] (viral load) in Serum or Plasma by Probe and signal amplification method
C0945037|HCV RNA SerPl bDNA-aCnc
C0945037|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C0945037|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.sig
C0945037|Hepatitis C virus RNA [Units/volume] (viral load) in Serum or Plasma by Probe and signal amplification method
C1508112|Hepatitis C virus RNA:LaCnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C1508112|HCV RNA SerPl PCR-Log IU
C1508112|Hepatitis C virus ribonucleic acid:Log Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1508112|Hepatitis C virus RNA [log units/volume] (viral load) in Serum or Plasma by Probe and target amplification method
C1623573|Hepatitis C virus RNA:LnCnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C1623573|HCV RNA SerPl bDNA-Log#
C1623573|Hepatitis C virus RNA [Log #/volume] (viral load) in Serum or Plasma by Probe and signal amplification method
C1623573|Hepatitis C virus ribonucleic acid:Log Number Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.sig
C1643191|HCV RNA SerPl bDNA-Log IU
C1643191|Hepatitis C virus RNA:LaCnc:Pt:Ser/Plas:Qn:Probe.amp.sig
C1643191|Hepatitis C virus ribonucleic acid:Log Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.sig
C1643191|Hepatitis C virus RNA [log units/volume] (viral load) in Serum or Plasma by Probe and signal amplification method
C1831320|Hepatitis C virus RNA:LnCnc:Pt:Ser/Plas:Qn:Probe.amp.tar
C1831320|HCV RNA SerPl PCR-Log#
C1831320|Hepatitis C virus ribonucleic acid:Log Number Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1831320|Hepatitis C virus RNA [Log #/volume] (viral load) in Serum or Plasma by Probe and target amplification method
C1977155|HCV RNA # CSF PCR
C1977155|Hepatitis C virus RNA:NCnc:Pt:CSF:Qn:Probe.amp.tar
C1977155|Hepatitis C virus ribonucleic acid:Number Concentration (count/vol):Point in time:Cerebral spinal fluid:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977155|Hepatitis C virus RNA [#/volume] (viral load) in Cerebral spinal fluid by Probe and target amplification method
C1977156|HCV RNA # Mar PCR
C1977156|Hepatitis C virus RNA:NCnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977156|Hepatitis C virus ribonucleic acid:Number Concentration (count/vol):Point in time:Marrow (bone):Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977156|Hepatitis C virus RNA [#/volume] (viral load) in Bone marrow by Probe and target amplification method
C1977157|Hepatitis C virus RNA:NCnc:Pt:Tiss:Qn:Probe.amp.tar
C1977157|HCV RNA # Tiss PCR
C1977157|Hepatitis C virus ribonucleic acid:Number Concentration (count/vol):Point in time:Tissue, unspecified:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977157|Hepatitis C virus RNA [#/volume] (viral load) in Tissue by Probe and target amplification method
C1977158|Hepatitis C virus RNA:LnCnc:Pt:XXX:Qn:Probe.amp.tar
C1977158|HCV RNA XXX PCR-Log#
C1977158|Hepatitis C virus ribonucleic acid:Log Number Concentration:Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977158|Hepatitis C virus RNA [Log #/volume] (viral load) in Unspecified specimen by Probe and target amplification method
C1977159|Hepatitis C virus RNA:LnCnc:Pt:CSF:Qn:Probe.amp.tar
C1977159|HCV RNA CSF PCR-Log#
C1977159|Hepatitis C virus ribonucleic acid:Log Number Concentration:Point in time:Cerebral spinal fluid:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977159|Hepatitis C virus RNA [Log #/volume] (viral load) in Cerebral spinal fluid by Probe and target amplification method
C1977160|Hepatitis C virus RNA:LnCnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977160|HCV RNA Mar PCR-Log#
C1977160|Hepatitis C virus ribonucleic acid:Log Number Concentration:Point in time:Marrow (bone):Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977160|Hepatitis C virus RNA [Log #/volume] (viral load) in Bone marrow by Probe and target amplification method
C1977161|HCV RNA Tiss PCR-Log#
C1977161|Hepatitis C virus RNA:LnCnc:Pt:Tiss:Qn:Probe.amp.tar
C1977161|Hepatitis C virus ribonucleic acid:Log Number Concentration:Point in time:Tissue, unspecified:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977161|Hepatitis C virus RNA [Log #/volume] (viral load) in Tissue by Probe and target amplification method
C1977162|Hepatitis C virus RNA:ACnc:Pt:XXX:Qn:Probe.amp.tar
C1977162|HCV RNA XXX PCR-aCnc
C1977162|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977162|Hepatitis C virus RNA [Units/volume] (viral load) in Unspecified specimen by Probe and target amplification method
C1977163|HCV RNA CSF PCR-aCnc
C1977163|Hepatitis C virus RNA:ACnc:Pt:CSF:Qn:Probe.amp.tar
C1977163|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Cerebral spinal fluid:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977163|Hepatitis C virus RNA [Units/volume] (viral load) in Cerebral spinal fluid by Probe and target amplification method
C1977164|HCV RNA Mar PCR-aCnc
C1977164|Hepatitis C virus RNA:ACnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977164|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Marrow (bone):Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977164|Hepatitis C virus RNA [Units/volume] (viral load) in Bone marrow by Probe and target amplification method
C1977165|HCV RNA Tiss PCR-aCnc
C1977165|Hepatitis C virus RNA:ACnc:Pt:Tiss:Qn:Probe.amp.tar
C1977165|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Tissue, unspecified:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977165|Hepatitis C virus RNA [Units/volume] (viral load) in Tissue by Probe and target amplification method
C1977166|Hepatitis C virus RNA:NCnc:Pt:XXX:Qn:Probe.amp.tar
C1977166|HCV RNA # XXX PCR
C1977166|Hepatitis C virus ribonucleic acid:Number Concentration (count/vol):Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977166|Hepatitis C virus RNA [#/volume] (viral load) in Unspecified specimen by Probe and target amplification method
C1977368|Hepatitis C virus RNA:LaCnc:Pt:CSF:Qn:Probe.amp.tar
C1977368|HCV RNA CSF PCR-Log IU
C1977368|Hepatitis C virus ribonucleic acid:Log Arbitrary Concentration:Point in time:Cerebral spinal fluid:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977368|Hepatitis C virus RNA [log units/volume] (viral load) in Cerebral spinal fluid by Probe and target amplification method
C1977369|HCV RNA Mar PCR-Log IU
C1977369|Hepatitis C virus RNA:LaCnc:Pt:Bone mar:Qn:Probe.amp.tar
C1977369|Hepatitis C virus ribonucleic acid:Log Arbitrary Concentration:Point in time:Marrow (bone):Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977369|Hepatitis C virus RNA [log units/volume] (viral load) in Bone marrow by Probe and target amplification method
C1977370|HCV RNA XXX PCR-Log IU
C1977370|Hepatitis C virus RNA:LaCnc:Pt:XXX:Qn:Probe.amp.tar
C1977370|Hepatitis C virus ribonucleic acid:Log Arbitrary Concentration:Point in time:To be specified in another part of the message:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977370|Hepatitis C virus RNA [log units/volume] (viral load) in Unspecified specimen by Probe and target amplification method
C1977373|HCV RNA Tiss PCR-Log IU
C1977373|Hepatitis C virus RNA:LaCnc:Pt:Tiss:Qn:Probe.amp.tar
C1977373|Hepatitis C virus ribonucleic acid:Log Arbitrary Concentration:Point in time:Tissue, unspecified:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977373|Hepatitis C virus RNA [log units/volume] (viral load) in Tissue by Probe and target amplification method
C1977893|HCV RNA Pnl SerPl PCR
C1977893|Hepatitis C virus RNA panel:-:Pt:Ser/Plas:Qn:Probe.amp.tar
C1977893|Hepatitis C virus ribonucleic acid panel:-:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar
C1977893|Hepatitis C virus RNA panel (viral load) in Serum or Plasma by Probe and target amplification method
C1369569|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar detection limit = 500 IU/mL
C1369569|HCV RNA SerPl PCR DL=500-aCnc
C1369569|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar detection limit = 500 IU/mL
C1369569|Hepatitis C virus RNA [Units/volume] (viral load) in Serum or Plasma by Probe and target amplification method detection limit = 500 IU/mL
C1369570|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar detection limit = 50 IU/mL
C1369570|HCV RNA SerPl PCR DL=50-aCnc
C1369570|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar detection limit = 50 IU/mL
C1369570|Hepatitis C virus RNA [Units/volume] (viral load) in Serum or Plasma by Probe and target amplification method detection limit = 50 iU/mL
C1977509|Hepatitis C virus RNA:ACnc:Pt:Ser/Plas:Qn:Probe.amp.tar detection limit = 5 IU/mL
C1977509|HCV RNA SerPl PCR DL=5-aCnc
C1977509|Hepatitis C virus ribonucleic acid:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:DNA Nucleic Acid Probe.amp.tar detection limit = 5 IU/mL
C1977509|Hepatitis C virus RNA [Units/volume] (viral load) in Serum or Plasma by Probe and target amplification method detection limit = 5 iU/mL
