C0809969|Cancer of kidney and renal pelvis
C0809971|Cancer of brain and nervous system
C0809972|Cancer; other and unspecified primary
C0810239|Cancer of ovary and other female genital organs
C0810243|Cancer; other primary
C1140680|Malignant neoplasm of ovary
C4048328|cervical cancer
C4048331|Cancer of bronchus; lung
C0005684|Malignant neoplasm of urinary bladder
C0006142|Malignant neoplasm of breast
C0007102|Malignant tumor of colon
C0007114|Malignant neoplasm of skin
C0007115|Malignant neoplasm of thyroid
C0153448|Malignant neoplasm of liver and intrahepatic bile ducts
C0153567|Uterine Cancer
C0153594|Malignant neoplasm of testis
C0153606|malignant tumor of male genital organ
C0278996|Cancer of Head and Neck
C0346647|Malignant neoplasm of pancreas
C0346890|Malignant neoplasm of other and unspecified urinary organs
C0348371|Malignant neoplasm of urinary organ, unspecified
C0348393|Malignant tumor of lymphoid hemopoietic and related tissue
C0376358|Malignant neoplasm of prostate
C0392920|Chemotherapy Regimen
C0497581|Other male genital malignant neoplasm
C0546837|Malignant neoplasm of esophagus
C0699791|Stomach Carcinoma
C0740458|cancer of uterus and cervix
C0809960|Cancer of rectum and anus
C0809962|Cancer of other GI organs; peritoneum
C0809964|Cancer; other respiratory and intrathoracic
C0809965|Cancer of bone and connective tissue
C0809967|Cancer of other female genital organs
C0809969|Cancer of kidney and renal pelvis
C0809971|Cancer of brain and nervous system
C0809972|Cancer; other and unspecified primary
C1140680|Cancer, Ovarian
C1140680|Cancers, Ovarian
C1140680|Ovarian Cancers
C1140680|Malignant neoplasm of ovary
C1140680|ovarian cancer
C1140680|Cancer of ovary
C1140680|malignant neoplasm of ovary (diagnosis)
C1140680|ovarian cancer (diagnosis)
C1140680|Ca ovary
C1140680|Cancers, Ovary
C1140680|Ovary Cancers
C1140680|malignant tumor of ovary
C1140680|Malign neopl ovary
C1140680|Cancer, Ovary
C1140680|Malignant tumour of ovary
C1140680|Malignant tumour of ovary (disorder)
C1140680|Ovaries--Cancer
C1140680|Ovarian cancer, NOS
C1140680|-- Ovarian Cancer
C1140680|Ovarian Ca
C1140680|Ovarian cancer NOS
C1140680|Cancer of the Ovary
C1140680|Ovary Cancer
C1140680|CA - Cancer of ovary
C1140680|Malignant tumor of ovary (disorder)
C1140680|Malignant Neoplasm of the Ovary
C1140680|Malignant Ovarian Neoplasm
C1140680|Malignant Ovarian Tumor
C1140680|Malignant Tumor of the Ovary
C0809967|Cancer of other female genital organs
C0809965|Cancer of bone and connective tissue
C0278996|Malignant tumor of head and neck (disorder)
C0278996|Malignant tumor of head and/or neck (disorder)
C0278996|Head and neck cancer
C0278996|Malignant tumour of head and/or neck
C0278996|Malignant tumor of head and/or neck
C0278996|Cancer of head and neck
C0278996|malignant neoplasm of head and/or neck (diagnosis)
C0278996|malignant neoplasm of head and/or neck
C0278996|Head and neck cancer, NOS
C0278996|Cancer of the Head and Neck
C0278996|Malignant tumor of head and neck
C0278996|Malignant tumour of head and neck
C0278996|Malignant Head and Neck Neoplasm
C0278996|Malignant Head and Neck Tumor
C0278996|Malignant Neoplasm of Head and Neck
C0278996|Malignant Neoplasm of the Head and Neck
C0278996|Malignant Tumor of the Head and Neck
C0007115|Malignant neoplasm of thyroid gland
C0007115|Malignant Thyroid Gland Neoplasm
C0007115|Malignant Thyroid Neoplasm
C0007115|Thyroid cancer
C0007115|malignant neoplasm of thyroid gland (diagnosis)
C0007115|Thyroid neoplasms malignant
C0007115|malignant tumor of thyroid gland
C0007115|Malign neopl thyroid
C0007115|Cancer of thyroid
C0007115|Malignant tumour of thyroid gland
C0007115|Malignant tumour of thyroid gland (disorder)
C0007115|-- Thyroid Cancer
C0007115|Thyroid neoplasm malignant
C0007115|Thyroid gland cancer
C0007115|Thyroid Ca
C0007115|Malignant tumor of thyroid gland (disorder)
C0007115|Malignant neoplasm of thyroid
C0007115|Malignant Neoplasm of the Thyroid Gland
C0007115|Malignant Neoplasm of the Thyroid
C0007115|Malignant Thyroid Gland Tumor
C0007115|Malignant Thyroid Tumor
C0007115|Malignant Tumor of Thyroid
C0007115|Malignant Tumor of the Thyroid Gland
C0007115|Malignant Tumor of the Thyroid
C0007115|Neoplasm malig;thyroid gland
C0007115|malignant neosplasm of the thyroid gland
C0809964|Cancer; other respiratory and intrathoracic
C0948216|adenocarcinoma of ovary (diagnosis)
C0948216|adenocarcinoma of ovary
C0948216|ovarian adenocarcinoma
C0948216|Adenocarcinoma of the Ovary
C0334495|malignant Brenner tumor of ovary (diagnosis)
C0334495|malignant Brenner tumor of ovary
C0334495|Malignant Brenner Tumor
C0334495|Brenner tumor, malignant
C0334495|Malignant Brenner tumour
C0334495|Brenner tumour, malignant
C0334495|Brenner tumor, malignant (morphologic abnormality)
C0334495|Brenner; tumor, malignant
C0334495|tumor; Brenner, malignant
C0334495|Malignant Brenner Tumor of the Ovary
C0334495|Malignant Ovarian Brenner Tumor
C1297991|malignant neoplasm involving left ovary by direct extension from endometrium
C1297991|malignant neoplasm involving left ovary by direct extension from endometrium (diagnosis)
C1297991|ovarian neoplasm left by direct extension from endometrium
C1297991|Malignant tumor involving left ovary by direct extension from endometrium (disorder)
C1297991|Malignant tumor involving left ovary by direct extension from endometrium
C1297991|Malignant tumour involving left ovary by direct extension from endometrium
C1297992|Malignant tumor involving left ovary by direct extension from fallopian tube (disorder)
C1297992|Malignant tumor involving left ovary by direct extension from fallopian tube
C1297992|Malignant tumour involving left ovary by direct extension from fallopian tube
C1297993|Malignant tumor involving left ovary by direct extension from right ovary (disorder)
C1297993|Malignant tumor involving left ovary by direct extension from right ovary
C1297993|Malignant tumour involving left ovary by direct extension from right ovary
C1297994|Malignant tumor involving left ovary by direct extension from uterine cervix (disorder)
C1297994|Malignant tumor involving left ovary by direct extension from uterine cervix
C1297994|Malignant tumour involving left ovary by direct extension from uterine cervix
C1297995|malignant neoplasm involving left ovary by direct extension from uterus
C1297995|ovarian neoplasm left by direct extension from uterus
C1297995|malignant neoplasm involving left ovary by direct extension from uterus (diagnosis)
C1297995|Malignant tumor involving left ovary by direct extension from uterus (disorder)
C1297995|Malignant tumor involving left ovary by direct extension from uterus
C1297995|Malignant tumour involving left ovary by direct extension from uterus
C1297998|Malignant tumor involving right ovary by direct extension from endometrium (disorder)
C1297998|Malignant tumor involving right ovary by direct extension from endometrium
C1297998|Malignant tumour involving right ovary by direct extension from endometrium
C1297999|ovarian neoplasm right by direct extension from fallopian tube
C1297999|malignant neoplasm involving right ovary by direct extension from fallopian tube (diagnosis)
C1297999|malignant neoplasm involving right ovary by direct extension from fallopian tube
C1297999|Malignant tumor involving right ovary by direct extension from fallopian tube (disorder)
C1297999|Malignant tumor involving right ovary by direct extension from fallopian tube
C1297999|Malignant tumour involving right ovary by direct extension from fallopian tube
C1298000|Malignant tumor involving right ovary by direct extension from left ovary (disorder)
C1298000|Malignant tumor involving right ovary by direct extension from left ovary
C1298000|Malignant tumour involving right ovary by direct extension from left ovary
C1298001|ovarian neoplasm right by direct extension from uterine cervix
C1298001|malignant neoplasm involving right ovary by direct extension from uterine cervix (diagnosis)
C1298001|malignant neoplasm involving right ovary by direct extension from uterine cervix
C1298001|Malignant tumor involving right ovary by direct extension from uterine cervix (disorder)
C1298001|Malignant tumor involving right ovary by direct extension from uterine cervix
C1298001|Malignant tumour involving right ovary by direct extension from uterine cervix
C1298026|malignant neoplasm involving left ovary by direct extension from vagina (diagnosis)
C1298026|malignant neoplasm involving left ovary by direct extension from vagina
C1298026|ovarian neoplasm left by direct extension from vagina
C1298026|Malignant tumor involving left ovary by direct extension from vagina (disorder)
C1298026|Malignant tumor involving left ovary by direct extension from vagina
C1298026|Malignant tumour involving left ovary by direct extension from vagina
C1298033|Malignant tumor involving right ovary by direct extension from uterus (disorder)
C1298033|Malignant tumor involving right ovary by direct extension from uterus
C1298033|Malignant tumour involving right ovary by direct extension from uterus
C1298034|Malignant tumor involving right ovary by direct extension from vagina (disorder)
C1298034|Malignant tumor involving right ovary by direct extension from vagina
C1298034|Malignant tumour involving right ovary by direct extension from vagina
C0346182|malignant teratoma of ovary (diagnosis)
C0346182|malignant teratoma of ovary
C0346182|Immature teratoma of ovary
C0346182|Immature teratoma of ovary (diagnosis)
C0346182|ovarian neoplasm malignant immature teratoma
C0346182|Immature teratoma of ovary (disorder)
C0346182|ovarian germ cell immature teratoma
C0346182|immature teratoma, ovarian germ cell
C0346182|teratoma, immature, ovarian germ cell
C0346182|Immature Germ Cell Teratoma of Ovary
C0346182|Immature Germ Cell Teratoma of the Ovary
C0346182|Immature Ovarian Teratoma
C0346182|Immature Teratoma of the Ovary
C0346182|Malignant Germ Cell Teratoma of Ovary
C0346182|Malignant Germ Cell Teratoma of the Ovary
C0346182|Malignant Ovarian Germ Cell Teratoma
C0346182|Malignant Ovarian Teratoma
C0346182|Malignant Teratoma of the Ovary
C0346182|Ovarian Immature Germ Cell Teratoma
C0346182|Ovarian Immature Teratoma
C2842146|Malignant neoplasm of right ovary
C2842147|Malignant neoplasm of unspecified ovary
C2016058|carcinoma simplex of ovary (diagnosis)
C2016058|carcinoma simplex of ovary
C2212041|adenocarcinoid tumor of ovary
C2212041|adenocarcinoid tumor of ovary (diagnosis)
C0392998|carcinosarcoma of ovary
C0392998|carcinosarcoma of ovary (diagnosis)
C0392998|Carcinosarcoma of ovary (disorder)
C0392998|Ovarian carcinosarcoma
C0392998|Malignant Mixed Mesodermal Müllerian Neoplasm of Ovary
C0392998|Ovarian Malignant Mixed Müllerian Tumor
C0392998|Malignant Mixed Mesodermal Müllerian Tumor of the Ovary
C0392998|Ovarian Malignant Mixed Müllerian Neoplasm
C0392998|Malignant Mixed Mesodermal Müllerian Neoplasm of the Ovary
C0392998|Ovarian Malignant Mixed Mesodermal Müllerian Tumor
C0392998|Malignant Mixed Mesodermal Müllerian Tumor of Ovary
C0392998|Ovarian Malignant Mixed Mesodermal Müllerian Neoplasm
C0392998|Ovarian Malignant Mixed Mesodermal (Müllerian) Tumor
C0392998|Ovarian Malignant Mesodermal (Müllerian) Mixed Tumor
C0392998|Mullerian sarcoma, ovarian malignant mixed mesodermal
C0392998|Mullerian tumor, ovarian malignant mixed mesodermal
C0392998|carcinosarcoma, ovarian
C0392998|malignant mixed mesodermal Mullerian tumor, ovarian
C0392998|Ovarian MMMT
C0392998|Carcinosarcoma of the Ovary
C2212004|malignant small cell neoplasm of ovary (diagnosis)
C2212004|ovarian neoplasm malignant small cell type
C2212004|malignant small cell neoplasm of ovary
C2011392|giant cell type neoplasm of ovary (diagnosis)
C2011392|ovarian neoplasm malignant giant cell type
C2011392|giant cell type neoplasm of ovary
C2018675|spindle cell type neoplasm of ovary (diagnosis)
C2018675|spindle cell type neoplasm of ovary
C2018675|ovarian neoplasm malignant spindle cell type
C2075635|ovarian neoplasm malignant clear cell type
C2075635|malignant clear cell type neoplasm of the ovary (diagnosis)
C2075635|malignant clear cell type neoplasm of the ovary
C2075635|clear cell type neoplasm of ovary
C0029925|Ovarian carcinoma
C0029925|carcinoma of ovary (diagnosis)
C0029925|carcinoma of ovary
C2212016|malignant epithelioid trophoblastic tumor of ovary
C2212016|malignant epithelioid trophoblastic tumor of ovary (diagnosis)
C0334525|malignant struma ovarii
C0334525|malignant struma ovarii (diagnosis)
C0334525|Struma ovarii, malignant
C0334525|Struma ovarii, malignant (morphologic abnormality)
C0334525|struma; ovarii, malignant
C0280746|Sarcoma of ovary
C0280746|Sarcoma of ovary (disorder)
C0280746|sarcoma of ovary (diagnosis)
C0280746|ovarian sarcoma
C0280746|sarcoma of the ovary
C0280746|sarcoma, ovarian
C1335161|fibrosarcoma of ovary (diagnosis)
C1335161|fibrosarcoma of ovary
C1335161|Fibrosarcoma of the Ovary
C1335161|Ovarian Fibrosarcoma
C2212040|myosarcoma of ovary (diagnosis)
C2212040|myosarcoma of ovary
C2212048|malignant gonadal neoplasm of ovary (diagnosis)
C2212048|malignant gonadal neoplasm of ovary
C2212049|malignant mesonephroma of ovary (diagnosis)
C2212049|malignant mesonephroma of ovary
C2212050|malignant lymphoma of ovary
C2212050|malignant lymphoma of ovary (diagnosis)
C2212053|malignant plasmacytoma of ovary
C2212053|malignant plasmacytoma of ovary (diagnosis)
C2212055|malignant mastocytosis of ovary (diagnosis)
C2212055|malignant mastocytosis of ovary
C2212056|Mullerian mixed tumor of ovary (diagnosis)
C2212056|Mullerian mixed tumor of ovary
C2212057|malignant mesodermal mixed tumor of ovary (diagnosis)
C2212057|malignant mesodermal mixed tumor of ovary
C2212058|adenocarcinofibroma of ovary
C2212058|adenocarcinofibroma of ovary (diagnosis)
C2217304|malignant neoplasm of ovary staging
C2217304|malignant neoplasm of ovary staging (diagnosis)
C2217304|malignant ovarian neoplasm staging
C2217304|malignant tumor of ovary staging
C2217304|ovarian cancer staging
C0346181|choriocarcinoma of ovary (diagnosis)
C0346181|choriocarcinoma of ovary
C0346181|Ovarian germ cell choriocarcinoma
C0346181|Choriocarcinoma of ovary (disorder)
C0346181|choriocarcinoma, ovarian germ cell
C0346181|Choriocarcinoma of the Ovary
C0346181|Germ Cell Choriocarcinoma of Ovary
C0346181|Germ Cell Choriocarcinoma of the Ovary
C0346181|Ovarian Choriocarcinoma
C2062541|malignant carcinoid tumor of ovary (diagnosis)
C2062541|malignant carcinoid tumor of ovary
C2011182|germinoma of ovary
C2011182|germinoma of ovary (diagnosis)
C2212020|ovarian adenocarcinoma scirrhous
C2212020|scirrhous adenocarcinoma of ovary (diagnosis)
C2212020|scirrhous adenocarcinoma of ovary
C2037342|ovarian adenocarcinoma superficial spreading
C2037342|superficial spreading adenocarcinoma of ovary (diagnosis)
C2037342|superficial spreading adenocarcinoma of ovary
C2212021|basal cell adenocarcinoma of ovary
C2212021|basal cell adenocarcinoma of ovary (diagnosis)
C2033126|papillary adenocarcinoma of ovary (diagnosis)
C2033126|papillary adenocarcinoma of ovary
C2189642|villous adenocarcinoma of ovary (diagnosis)
C2189642|villous adenocarcinoma of ovary
C2016016|adenocarcinoma in villous adenoma of ovary (diagnosis)
C2016016|adenocarcinoma in villous adenoma of ovary
C2016015|adenocarcinoma in tubulovillous adenoma of ovary
C2016015|adenocarcinoma in tubulovillous adenoma of ovary (diagnosis)
C2212022|mixed cell adenocarcinoma of ovary
C2212022|mixed cell adenocarcinoma of ovary (diagnosis)
C2212026|endocervical type mucinous adenocarcinoma of ovary (diagnosis)
C2212026|endocervical type mucinous adenocarcinoma of ovary
C2212027|mucin-producing adenocarcinoma of ovary (diagnosis)
C2212027|mucin-producing adenocarcinoma of ovary
C2212028|adenocarcinoma of ovary with metaplasia
C2212028|adenocarcinoma of ovary with metaplasia (diagnosis)
C2212028|ovarian adenocarcinoma with metaplasia
C2212029|adenocarcinoma of ovary with squamous metaplasia
C2212029|ovarian adenocarcinoma with squamous metaplasia
C2212029|adenocarcinoma of ovary with squamous metaplasia (diagnosis)
C2016017|adenocarcinoma with cartilaginous or osseous metaplasia of ovary
C2016017|adenocarcinoma of ovary with cartilaginous and osseous metaplasia (diagnosis)
C2016017|adenocarcinoma of ovary with cartilaginous and osseous metaplasia
C2016017|ovarian adenocarcinoma with cartilaginous or osseous metaplasia
C2016017|ovarian adenocarcinoma with cartilaginous and osseous metaplasia
C2212030|ovarian adenocarcinoma with spindle cell metaplasia
C2212030|adenocarcinoma of ovary with spindle cell metaplasia
C2212030|adenocarcinoma of ovary with spindle cell metaplasia (diagnosis)
C2212031|adenocarcinoma of ovary with apocrine metaplasia
C2212031|ovarian adenocarcinoma with apocrine metaplasia
C2212031|adenocarcinoma of ovary with apocrine metaplasia (diagnosis)
C2016018|adenocarcinoma of ovary with neuroendocrine differentiation
C2016018|adenocarcinoma of ovary with neuroendocrine differentiation (diagnosis)
C2016018|ovarian adenocarcinoma with neuroendocrine differentiation
C1335167|mucinous adenocarcinoma of ovary (diagnosis)
C1335167|mucinous adenocarcinoma of ovary
C1335167|Mucinous Adenocarcinoma of the Ovary
C1335167|Mucinous Carcinoma of Ovary
C1335167|Mucinous Carcinoma of the Ovary
C1335167|Ovarian Mucinous Adenocarcinoma
C1335167|Ovarian Mucinous Carcinoma
C0346163|Ovarian Endometrioid Adenocarcinoma NOS
C0346163|endometrioid adenocarcinoma of ovary (diagnosis)
C0346163|endometrioid adenocarcinoma of ovary
C0346163|Ovarian endometrioid carcinoma
C0346163|ovarian malignant carcinoma endometrioid
C0346163|endometrioid carcinoma of ovary
C0346163|endometrioid carcinoma of ovary (diagnosis)
C0346163|Ovarian Endometrioid Adenocarcinoma Not Otherwise Specified
C0346163|Endometrioid carcinoma ovary
C0346163|Endometrioid carcinoma ovary (disorder)
C0346163|ovarian endometrioid adenocarcinoma
C0346163|adenocarcinoma of the ovary, endometrioid
C0346163|endometrioid adenocarcinoma of the ovary
C0346163|ovarian cancer, endometrioid adenocarcinoma
C0346163|ovary cancer, endometrioid adenocarcinoma
C0346163|Endometrioid Cancer of Ovary
C0346163|Endometrioid Cancer of the Ovary
C0346163|Endometrioid Carcinoma of the Ovary
C0346163|Ovarian Endometrioid Cancer
C1518693|clear cell adenocarcinoma of ovary (diagnosis)
C1518693|clear cell adenocarcinoma of ovary
C1518693|Ovarian Clear Cell Adenocarcinoma
C2977928|Malignant neoplasm of left ovary
C2212005|malignant epithelioma of ovary
C2212005|malignant epithelioma of ovary (diagnosis)
C2111648|large cell carcinoma of ovary (diagnosis)
C2111648|large cell carcinoma of ovary
C1335174|large cell neuroendocrine carcinoma of ovary (diagnosis)
C1335174|large cell neuroendocrine carcinoma of ovary
C1335174|Ovarian Large Cell NEC
C1335174|Large Cell Neuroendocrine Carcinoma of the Ovary
C1335174|Large-Cell Neuroendocrine Carcinoma of Ovary
C1335174|Large-Cell Neuroendocrine Carcinoma of the Ovary
C1335174|Non-Small-Cell Type Neuroendocrine Carcinoma of Ovary
C1335174|Non-Small-Cell Type Neuroendocrine Carcinoma of the Ovary
C1335174|Ovarian Non-Small-Cell Type Neuroendocrine Carcinoma
C1335174|Ovarian Large Cell Neuroendocrine Carcinoma
C2111649|ovarian malignant carcinoma large cell with rhabdoid phenotype
C2111649|large cell carcinoma of ovary with rhabdoid phenotype
C2111649|large cell carcinoma of ovary with rhabdoid phenotype (diagnosis)
C2012100|glassy cell carcinoma of ovary (diagnosis)
C2012100|glassy cell carcinoma of ovary
C0334398|malignant thecoma of ovary (diagnosis)
C0334398|malignant thecoma of ovary
C0334398|THECOMA, OVARIAN, MALIGNANT
C0334398|Malignant Ovarian Thecal Cell Neoplasm
C0334398|Thecoma, Malignant
C0334398|Malignant Thecal Cell Tumor of the Ovary
C0334398|Malignant Thecal Cell Neoplasm of Ovary
C0334398|Malignant Thecal Cell Tumor of Ovary
C0334398|Malignant Thecoma of the Ovary
C0334398|Malignant Ovarian Thecal Cell Tumor
C0334398|Malignant Thecal Cell Neoplasm of the Ovary
C0334398|Malignant thecoma
C0334398|Thecoma, malignant (morphologic abnormality)
C0334398|malignant; thecoma
C0334398|thecoma; malignant
C0334398|Malignant Ovarian Thecoma
C0346167|undifferentiated carcinoma of ovary
C0346167|anaplastic carcinoma of ovary
C0346167|anaplastic carcinoma of ovary (diagnosis)
C0346167|undifferentiated carcinoma of ovary (diagnosis)
C0346167|Undifferentiated ovarian cancer
C0346167|Undifferentiated carcinoma of ovary (disorder)
C0346167|Anaplastic Carcinoma of the Ovary
C0346167|Anaplastic Ovarian Carcinoma
C0346167|Undifferentiated Carcinoma of the Ovary
C0346167|Undifferentiated Ovarian Carcinoma
C2082449|pleomorphic carcinoma of ovary
C2082449|pleomorphic carcinoma of ovary (diagnosis)
C2011259|giant cell carcinoma of ovary (diagnosis)
C2011259|giant cell carcinoma of ovary
C2018399|spindle cell carcinoma of ovary
C2018399|spindle cell carcinoma of ovary (diagnosis)
C2011224|giant cell and spindle cell carcinoma of ovary
C2011224|giant cell and spindle cell carcinoma of ovary (diagnosis)
C2142929|pseudosarcomatous carcinoma of ovary (diagnosis)
C2142929|pseudosarcomatous carcinoma of ovary
C2111811|polygonal cell carcinoma of ovary (diagnosis)
C2111811|polygonal cell carcinoma of ovary
C2016059|carcinoma of ovary with osteoclast-like giant cells (diagnosis)
C2016059|carcinoma of ovary with osteoclast-like giant cells
C2212006|small cell carcinoma of ovary (diagnosis)
C2212006|small cell carcinoma of ovary
C2212006|Ovarian Small Cell Neuroendocrine Carcinoma
C2212006|Ovarian Small Cell NEC
C2212006|Ovarian Small Cell Carcinoma
C2033226|papillary carcinoma of ovary
C2033226|papillary carcinoma of ovary (diagnosis)
C2033303|papillary squamous cell carcinoma of ovary (diagnosis)
C2033303|papillary squamous cell carcinoma of ovary
C2189355|verrucous carcinoma of ovary (diagnosis)
C2189355|verrucous carcinoma of ovary
C2019443|squamous cell carcinoma of ovary (diagnosis)
C2019443|squamous cell carcinoma of ovary
C2019443|Ovarian Squamous Cell Carcinoma
C2109313|keratinizing squamous cell carcinoma of ovary
C2109313|keratinizing squamous cell carcinoma of ovary (diagnosis)
C2212007|nonkeratinizing large cell squamous carcinoma cell of ovary (diagnosis)
C2212007|nonkeratinizing large cell squamous carcinoma cell of ovary
C2212007|ovarian malignant carcinoma squamous cell large cell nonkeratinizing
C2212008|ovarian malignant carcinoma squamous cell small cell nonkeratinizing
C2212008|nonkeratinizing small cell squamous cell carcinoma of ovary (diagnosis)
C2212008|nonkeratinizing small cell squamous cell carcinoma of ovary
C2018560|spindle cell squamous cell carcinoma of ovary (diagnosis)
C2018560|spindle cell squamous cell carcinoma of ovary
C2212009|adenoid squamous cell carcinoma of ovary
C2212009|adenoid squamous cell carcinoma of ovary (diagnosis)
C2212010|microinvasive squamous cell carcinoma of ovary (diagnosis)
C2212010|microinvasive squamous cell carcinoma of ovary
C2019488|ovarian malignant carcinoma squamous cell with horn formation
C2019488|squamous cell carcinoma with horn formation of ovary
C2019488|squamous cell carcinoma of ovary with horn formation (diagnosis)
C2019488|squamous cell carcinoma of ovary with horn formation
C2212012|myxosarcoma of ovary
C2212012|myxosarcoma of ovary (diagnosis)
C2212013|Ovarian Serous Adenocarcinofibroma
C2212013|serous adenocarcinofibroma of ovary
C2212013|serous adenocarcinofibroma of ovary (diagnosis)
C2212014|mucinous adenocarcinofibroma of ovary
C2212014|mucinous adenocarcinofibroma of ovary (diagnosis)
C2212014|Ovarian Mucinous Adenocarcinofibroma
C2212014|Ovarian Mucinous Malignant Adenofibroma
C2212017|adenosquamous carcinoma of ovary (diagnosis)
C2212017|adenosquamous carcinoma of ovary
C2212017|Ovarian Adenoacanthoma
C2212017|Ovarian Adenosquamous Carcinoma
C2212017|Ovarian Endometrioid Adenocarcinoma with Squamous Differentiation
C2212018|epithelial-myoepithelial carcinoma of ovary
C2212018|epithelial-myoepithelial carcinoma of ovary (diagnosis)
C2017451|solid carcinoma of ovary (diagnosis)
C2017451|solid carcinoma of ovary
C2012542|granular cell carcinoma of ovary (diagnosis)
C2012542|granular cell carcinoma of ovary
C2212019|medullary carcinoma of ovary
C2212019|medullary carcinoma of ovary (diagnosis)
C2212023|secretory variant endometrioid adenocarcinoma of ovary (diagnosis)
C2212023|secretory variant endometrioid adenocarcinoma of ovary
C2075006|ciliated cell variant endometrioid adenocarcinoma of ovary (diagnosis)
C2075006|ciliated cell variant endometrioid adenocarcinoma of ovary
C2212024|endometrioid adenofibroma of ovary (diagnosis)
C2212024|endometrioid adenofibroma of ovary
C2212024|Ovarian Endometrioid Adenofibroma
C2018502|spindle cell sarcoma of ovary (diagnosis)
C2018502|spindle cell sarcoma of ovary
C2011316|giant cell sarcoma of ovary (diagnosis)
C2011316|giant cell sarcoma of ovary
C2212032|small cell sarcoma of ovary (diagnosis)
C2212032|small cell sarcoma of ovary
C2212033|epithelioid sarcoma of ovary
C2212033|epithelioid sarcoma of ovary (diagnosis)
C2188139|undifferentiated sarcoma of ovary (diagnosis)
C2188139|undifferentiated sarcoma of ovary
C2188139|High Grade Ovarian Endometrioid Stromal Sarcoma
C2188139|Undifferentiated Ovarian Sarcoma
C2016060|desmoplastic small round cell tumor of ovary
C2016060|desmoplastic small round cell tumor of ovary (diagnosis)
C2212034|malignant enterochromaffin cell carcinoid tumor of ovary (diagnosis)
C2212034|malignant enterochromaffin cell carcinoid tumor of ovary
C2046334|histiocytic sarcoma of ovary
C2046334|histiocytic sarcoma of ovary (diagnosis)
C2111171|Langerhans cell sarcoma of ovary (diagnosis)
C2111171|Langerhans cell sarcoma of ovary
C2077757|interdigitating dendritic cell sarcoma of ovary
C2077757|interdigitating dendritic cell sarcoma of ovary (diagnosis)
C2212036|follicular dendritic cell sarcoma of ovary
C2212036|follicular dendritic cell sarcoma of ovary (diagnosis)
C2212037|malignant enterochromaffin-like cell carcinoid tumor of ovary
C2212037|malignant enterochromaffin-like cell carcinoid tumor of ovary (diagnosis)
C2212038|fibromyxosarcoma of ovary (diagnosis)
C2212038|fibromyxosarcoma of ovary
C2212039|fascial fibrosarcoma of ovary (diagnosis)
C2212039|fascial fibrosarcoma of ovary
C2016039|infantile fibrosarcoma of ovary (diagnosis)
C2016039|infantile fibrosarcoma of ovary
C2016081|malignant solitary fibrous tumor of ovary
C2016081|malignant solitary fibrous tumor of ovary (diagnosis)
C2016056|goblet cell carcinoid of ovary
C2016056|goblet cell carcinoid of ovary (diagnosis)
C2106919|composite carcinoid tumor of ovary (diagnosis)
C2106919|composite carcinoid tumor of ovary
C2016057|neuroendocrine carcinoma of ovary
C2016057|neuroendocrine carcinoma of ovary (diagnosis)
C2212042|atypical carcinoid tumor of ovary (diagnosis)
C2212042|atypical carcinoid tumor of ovary
C2212043|angiomyosarcoma of ovary
C2212043|angiomyosarcoma of ovary (diagnosis)
C2075522|clear cell adenocarcinofibroma of ovary (diagnosis)
C2075522|clear cell adenocarcinofibroma of ovary
C2075522|Ovarian Clear Cell Adenocarcinofibroma
C2075522|Ovarian Clear Cell Malignant Adenofibroma
C2212044|embryonal carcinosarcoma of ovary (diagnosis)
C2212044|embryonal carcinosarcoma of ovary
C2212045|malignant myoepithelioma of ovary
C2212045|malignant myoepithelioma of ovary (diagnosis)
C2033248|papillary cystadenocarcinoma of ovary
C2033248|papillary cystadenocarcinoma of ovary (diagnosis)
C2212047|signet ring cell carcinoma of ovary (diagnosis)
C2212047|signet ring cell carcinoma of ovary
C1335178|serous surface papillary carcinoma of ovary (diagnosis)
C1335178|serous surface papillary carcinoma of ovary
C1335178|Serous Surface Papillary Carcinoma of the Ovary
C1335178|Ovarian Serous Surface Papillary Adenocarcinoma
C2016082|teratoma of ovary with malignant transformation
C2016082|teratoma of ovary with malignant transformation (diagnosis)
C2217294|malignant neoplasm of ovary stage Ia
C2217294|malignant neoplasm of ovary stage Ia (diagnosis)
C2217294|malignant ovarian neoplasm stage Ia
C2217294|malignant tumor of ovary stage Ia
C2217294|ovarian cancer stage Ia
C2217295|malignant ovarian neoplasm stage Ib
C2217295|malignant neoplasm of ovary stage Ib
C2217295|malignant neoplasm of ovary stage Ib (diagnosis)
C2217295|malignant tumor of ovary stage Ib
C2217295|ovarian cancer stage Ib
C2217296|malignant neoplasm of ovary stage Ic
C2217296|malignant neoplasm of ovary stage Ic (diagnosis)
C2217296|malignant ovarian neoplasm stage Ic
C2217296|ovarian cancer stage Ic
C2217296|malignant tumor of ovary stage Ic
C2217297|malignant neoplasm of ovary stage IIa (diagnosis)
C2217297|malignant ovarian neoplasm stage IIa
C2217297|malignant neoplasm of ovary stage IIa
C2217297|ovarian cancer stage IIa
C2217297|malignant tumor of ovary stage IIa
C2217298|malignant neoplasm of ovary stage IIb (diagnosis)
C2217298|malignant ovarian neoplasm stage IIb
C2217298|malignant neoplasm of ovary stage IIb
C2217298|malignant tumor of ovary stage IIb
C2217298|ovarian cancer stage IIb
C2217299|malignant neoplasm of ovary stage IIc
C2217299|malignant neoplasm of ovary stage IIc (diagnosis)
C2217299|malignant ovarian neoplasm stage IIc
C2217299|malignant tumor of ovary stage IIc
C2217299|ovarian cancer stage IIc
C2217300|malignant neoplasm of ovary stage IIIa (diagnosis)
C2217300|malignant ovarian neoplasm stage IIIa
C2217300|malignant neoplasm of ovary stage IIIa
C2217300|malignant tumor of ovary stage IIIa
C2217300|ovarian cancer stage IIIa
C2217301|malignant ovarian neoplasm stage IIIb
C2217301|malignant neoplasm of ovary stage IIIb
C2217301|malignant neoplasm of ovary stage IIIb (diagnosis)
C2217301|malignant tumor of ovary stage IIIb
C2217301|ovarian cancer stage IIIb
C2217302|malignant neoplasm of ovary stage IIIc (diagnosis)
C2217302|malignant ovarian neoplasm stage IIIc
C2217302|malignant neoplasm of ovary stage IIIc
C2217302|ovarian cancer stage IIIc
C2217302|malignant tumor of ovary stage IIIc
C2217303|malignant neoplasm of ovary stage IV
C2217303|malignant ovarian neoplasm stage IV
C2217303|malignant neoplasm of ovary stage IV (diagnosis)
C2217303|malignant tumor of ovary stage IV
C2217303|ovarian cancer stage IV
C0346188|yolk sac tumor of ovary (diagnosis)
C0346188|yolk sac tumor of ovary
C0346188|Ovarian germ cell endodermal sinus tumour
C0346188|Endodermal sinus tumor of ovary
C0346188|Endodermal sinus tumor of ovary (diagnosis)
C0346188|ovarian neoplasm malignant germ cell tumor endodermal sinus
C0346188|Ovarian germ cell yolk sac tumor
C0346188|Ovarian germ cell endodermal sinus tumor
C0346188|Ovarian germ cell yolk sac tumour
C0346188|Endodermal sinus tumour of ovary
C0346188|Yolk sac tumour of ovary
C0346188|Endodermal sinus tumor of ovary (disorder)
C0346188|endodermal sinus tumor, ovarian germ cell
C0346188|ovarian germ cell yolk sac carcinoma
C0346188|yolk sac carcinoma, ovarian germ cell
C0346188|Endodermal Sinus Neoplasm of Ovary
C0346188|Endodermal Sinus Neoplasm of the Ovary
C0346188|Endodermal Sinus Tumor of the Ovary
C0346188|Germ Cell Endodermal Sinus Neoplasm of Ovary
C0346188|Germ Cell Endodermal Sinus Neoplasm of the Ovary
C0346188|Germ Cell Endodermal Sinus Tumor of Ovary
C0346188|Germ Cell Endodermal Sinus Tumor of the Ovary
C0346188|Ovarian Endodermal Sinus Neoplasm
C0346188|Ovarian Endodermal Sinus Tumor
C0346188|Ovarian Germ Cell Endodermal Sinus Neoplasm
C0346188|Ovarian Yolk Sac Neoplasm
C0346188|Ovarian Yolk Sac Tumor
C0346188|Yolk Sac Neoplasm of Ovary
C0346188|Yolk Sac Neoplasm of the Ovary
C0346188|Yolk Sac Tumor of the Ovary
C0346161|Carcinoma of ovary
C0346161|Malignant epithelial tumor of ovary
C0346161|Malignant epithelial tumour of ovary
C0346161|Malignant epithelial tumor of ovary (disorder)
C3469523|ovarian cancer susceptibility (diagnosis)
C3469523|ovarian cancer susceptibility
C3469523|OVARIAN CANCER, SUSCEPTIBILITY TO
C0153577|Malignant neoplasm of ovary and other uterine adnexa
C0153577|Ca ovary/other uterine adnexa
C0153577|Ca ovary/other uterine adnexa (disorder)
C0153577|Malignant neoplasm of ovary and other uterine adnexa (disorder)
C1299247|Primary malignant neoplasm of ovary and other uterine adnexa (disorder)
C1299247|Primary malignant neoplasm of ovary and other uterine adnexa
C1306468|Primary malignant neoplasm of ovary
C1306468|ovarian malignant neoplasm primary
C1306468|Primary malignant neoplasm of ovary (diagnosis)
C1306468|Primary malignant neoplasm of ovary (disorder)
C1299248|Carcinoma of ovary and other uterine adnexa (disorder)
C1299248|Carcinoma of ovary and other uterine adnexa
C3693886|malignant neoplasm involving left ovary by direct extension from fallopian tube (diagnosis)
C3693886|malignant neoplasm involving left ovary by direct extension from fallopian tube
C3693886|ovarian neoplasm left by direct extension from fallopian tube
C0346180|OVARIAN GERM CELL CANCER
C0346180|Ovarian germ cell neoplasms malignant
C0346180|malignant germ cell tumor of ovary (diagnosis)
C0346180|malignant germ cell tumor of ovary
C0346180|ovarian neoplasm malignant germ cell tumor
C0346180|Ovarian germ cell cancer NOS
C0346180|Malignant germ cell tumour of ovary
C0346180|Malignant germ cell tumor of ovary (disorder)
C0346180|Malignant Ovarian Germ Cell Neoplasm
C0346180|Malignant Germ Cell Neoplasm of Ovary
C0346180|Malignant Germ Cell Neoplasm of the Ovary
C0346180|Malignant Germ Cell Tumor of the Ovary
C0346180|Malignant Ovarian Germ Cell Tumor
C3693885|malignant neoplasm involving left ovary by direct extension from right ovary
C3693885|malignant neoplasm involving left ovary by direct extension from right ovary (diagnosis)
C3693885|ovarian neoplasm left by direct extension from right ovary
C3647143|Secondary malignant neoplasm of ovary
C3647143|metastasis of malignant neoplasm to ovary (diagnosis)
C3647143|metastasis of malignant neoplasm to ovary
C3647143|Metastases to ovary
C3647143|Second malig neo ovary
C3647143|secondary malignant neoplasm of ovary (diagnosis)
C3647143|secondary malignant neoplasm genital organs ovary
C3647143|Metastasis to ovary (disorder)
C3647143|Metastasis to ovary
C3647143|Metastatic Malignant Neoplasm to the Ovary
C3647143|Metastatic Malignant Neoplasm in the Ovary
C3647143|Ovarian metastases
C3647143|Metastasis to ovary [Ambiguous]
C3647143|Metastatic Malignant Tumor to the Ovary
C3647143|Ovarian Metastasis
C3693879|ovarian neoplasm right by direct extension from vagina
C3693879|malignant neoplasm involving right ovary by direct extension from vagina (diagnosis)
C3693879|malignant neoplasm involving right ovary by direct extension from vagina
C3693881|ovarian neoplasm right by direct extension from left ovary
C3693881|malignant neoplasm involving right ovary by direct extension from left ovary (diagnosis)
C3693881|malignant neoplasm involving right ovary by direct extension from left ovary
C0346175|malignant granulosa cell tumor of ovary
C0346175|malignant granulosa cell tumor of ovary (diagnosis)
C0346175|ovarian neoplasm malignant granulosa cell
C0346175|malignant granulosa cell neoplasm of ovary
C0346175|malignant granulosa cell neoplasm of ovary (diagnosis)
C0346175|Malignant granulosa cell tumour of ovary
C0346175|Malignant granulosa cell tumor of ovary (disorder)
C0346175|Malignant Granulosa Cell Neoplasm of the Ovary
C0346175|Malignant Granulosa Cell Tumor of the Ovary
C0346175|Malignant Ovarian Granulosa Cell Neoplasm
C0346175|Malignant Ovarian Granulosa Cell Tumor
C3693882|malignant neoplasm involving right ovary by direct extension from endometrium (diagnosis)
C3693882|ovarian neoplasm right by direct extension from endometrium
C3693882|malignant neoplasm involving right ovary by direct extension from endometrium
C3693884|malignant neoplasm involving left ovary by direct extension from uterine cervix (diagnosis)
C3693884|malignant neoplasm involving left ovary by direct extension from uterine cervix
C3693884|ovarian neoplasm left by direct extension from uterine cervix
C3693880|ovarian neoplasm right by direct extension from uterus
C3693880|malignant neoplasm involving right ovary by direct extension from uterus (diagnosis)
C3693880|malignant neoplasm involving right ovary by direct extension from uterus
C3250633|malig ovarian neoplasm tnm staging distant metastasis (m) m0 (diagnosis)
C3250633|malig ovarian neoplasm tnm staging distant metastasis (m) m0
C3250634|malig ovarian neoplasm tnm staging distant metastasis (m) m1
C3250634|malig ovarian neoplasm tnm staging distant metastasis (m) m1 (diagnosis)
C3250632|malig ovarian neoplasm tnm staging distant metastasis (m) (diagnosis)
C3250632|malig ovarian neoplasm tnm staging distant metastasis (m)
C4030088|biopsy ovary malignant neoplasm fibrosarcoma solitary fibrous tumor
C4030088|biopsy ovary malignant neoplasm fibrosarcoma solitary fibrous tumor (procedure)
C4030115|biopsy ovary malignant lymphoma precursor cell lymphoblastic (procedure)
C4030115|biopsy ovary malignant lymphoma precursor cell lymphoblastic
C4030090|biopsy ovary malignant neoplasm fibrosarcoma fibromyxosarcoma (procedure)
C4030090|biopsy ovary malignant neoplasm fibrosarcoma fibromyxosarcoma
C4030122|biopsy ovary malignant lymphoma mantle cell
C4030122|biopsy ovary malignant lymphoma mantle cell (procedure)
C4030071|biopsy ovary malignant neoplasm immature teratoma
C4030071|biopsy ovary malignant neoplasm immature teratoma (procedure)
C4030060|biopsy ovary malignant neoplasm plasmacytoma
C4030060|biopsy ovary malignant neoplasm plasmacytoma (procedure)
C4030059|biopsy ovary malignant neoplasm plasmacytoma extramedullary
C4030059|biopsy ovary malignant neoplasm plasmacytoma extramedullary (procedure)
C4030166|biopsy ovary malignant carcinoma medullary (procedure)
C4030166|biopsy ovary malignant carcinoma medullary
C4030051|biopsy ovary malignant neoplasm teratoma teratocarcinoma
C4030051|biopsy ovary malignant neoplasm teratoma teratocarcinoma (procedure)
C4030045|biopsy ovary malignant sarcoma histiocytic
C4030045|biopsy ovary malignant sarcoma histiocytic (procedure)
C4030186|biopsy ovary malig lymphoma precursor cell lymphoblastic t-cell
C4030186|biopsy ovary malig lymphoma precursor cell lymphoblastic t-cell (procedure)
C4030114|biopsy ovary malignant lymphoma small b-cell lymphocytic
C4030114|biopsy ovary malignant lymphoma small b-cell lymphocytic (procedure)
C4030201|biopsy ovary malig adenocarcinoma metaplastic cartilaginous & osseous (procedure)
C4030201|biopsy ovary malig adenocarcinoma metaplastic cartilaginous & osseous
C4030104|biopsy ovary malignant neoplasm carcinoid tumor composite (procedure)
C4030104|biopsy ovary malignant neoplasm carcinoid tumor composite
C4030191|biopsy ovary malig lymphoma hodgkin's lymphocyt deplet reticular
C4030191|biopsy ovary malig lymphoma hodgkin's lymphocyt deplet reticular (procedure)
C4030058|biopsy ovary malignant neoplasm sarcoma (procedure)
C4030058|biopsy ovary malignant neoplasm sarcoma
C4030044|biopsy ovary malignant sarcoma interdigitating dendritic cell (procedure)
C4030044|biopsy ovary malignant sarcoma interdigitating dendritic cell
C4030040|biopsy ovary malignant sarcoma small cell
C4030040|biopsy ovary malignant sarcoma small cell (procedure)
C4030168|biopsy ovary malignant carcinoma large cell neuroendocrine (procedure)
C4030168|biopsy ovary malignant carcinoma large cell neuroendocrine
C4030160|biopsy ovary malignant carcinoma serous surface papillary (procedure)
C4030160|biopsy ovary malignant carcinoma serous surface papillary
C4030054|biopsy ovary malignant neoplasm teratoma (procedure)
C4030054|biopsy ovary malignant neoplasm teratoma
C4030102|biopsy ovary malignant neoplasm carcinoid tumor goblet cell (procedure)
C4030102|biopsy ovary malignant neoplasm carcinoid tumor goblet cell
C4030065|biopsy ovary malignant neoplasm myosarcoma
C4030065|biopsy ovary malignant neoplasm myosarcoma (procedure)
C4030134|biopsy ovary malignant lymphoma follicular grade 3 (procedure)
C4030134|biopsy ovary malignant lymphoma follicular grade 3
C4030129|biopsy ovary malignant lymphoma hodgkin's lymphocytic depletion
C4030129|biopsy ovary malignant lymphoma hodgkin's lymphocytic depletion (procedure)
C4030083|biopsy ovary malignant neoplasm germinoma nonseminomatous (procedure)
C4030083|biopsy ovary malignant neoplasm germinoma nonseminomatous
C4030112|biopsy ovary malignant neoplasm adenocarcinofibroma clear cell (procedure)
C4030112|biopsy ovary malignant neoplasm adenocarcinofibroma clear cell
C4030049|biopsy ovary malignant sarcoma desmoplastic small round cell
C4030049|biopsy ovary malignant sarcoma desmoplastic small round cell (procedure)
C4030135|biopsy ovary malignant lymphoma follicular grade 2 (procedure)
C4030135|biopsy ovary malignant lymphoma follicular grade 2
C4030177|biopsy ovary malignant carcinoma embryonal yolk sac tumor (procedure)
C4030177|biopsy ovary malignant carcinoma embryonal yolk sac tumor
C4030097|biopsy ovary malignant neoplasm carcinosarcoma myoepithelioma
C4030097|biopsy ovary malignant neoplasm carcinosarcoma myoepithelioma (procedure)
C4030111|biopsy ovary malignant neoplasm adenocarcinofibroma mucinous
C4030111|biopsy ovary malignant neoplasm adenocarcinofibroma mucinous (procedure)
C4030039|biopsy ovary malignant sarcoma spindle cell
C4030039|biopsy ovary malignant sarcoma spindle cell (procedure)
C4030064|biopsy ovary malignant neoplasm myosarcoma angiomyosarcoma
C4030064|biopsy ovary malignant neoplasm myosarcoma angiomyosarcoma (procedure)
C4030139|biopsy ovary malignant lymphoma burkitt's (procedure)
C4030139|biopsy ovary malignant lymphoma burkitt's
C4030120|biopsy ovary malignant lymphoma mature t-cell (procedure)
C4030120|biopsy ovary malignant lymphoma mature t-cell
C4030179|biopsy ovary malignant carcinoma embryonal
C4030179|biopsy ovary malignant carcinoma embryonal (procedure)
C4030178|biopsy ovary malignant carcinoma embryonal polyembryoma
C4030178|biopsy ovary malignant carcinoma embryonal polyembryoma (procedure)
C4030184|biopsy ovary malig neoplasm teratoma with malignant transformation (procedure)
C4030184|biopsy ovary malig neoplasm teratoma with malignant transformation
C4030062|biopsy ovary malignant neoplasm myosarcoma leiomyosarcoma epithelioid
C4030062|biopsy ovary malignant neoplasm myosarcoma leiomyosarcoma epithelioid (procedure)
C4030095|biopsy ovary malignant neoplasm clear cell type (procedure)
C4030095|biopsy ovary malignant neoplasm clear cell type
C4030069|biopsy ovary malignant neoplasm mastocytosis
C4030069|biopsy ovary malignant neoplasm mastocytosis (procedure)
C4030043|biopsy ovary malignant sarcoma langerhans cell
C4030043|biopsy ovary malignant sarcoma langerhans cell (procedure)
C4030038|biopsy ovary malignant sarcoma undifferentiated (procedure)
C4030038|biopsy ovary malignant sarcoma undifferentiated
C4030189|biopsy ovary malig lymphoma hodgkin's nodular sclerosis grade 2
C4030189|biopsy ovary malig lymphoma hodgkin's nodular sclerosis grade 2 (procedure)
C4030132|biopsy ovary malignant lymphoma hodgkin's (procedure)
C4030132|biopsy ovary malignant lymphoma hodgkin's
C4030586|biopsy ovary malig lymphoma hodgkin's nodular sclerosis grade 1
C4030586|biopsy of ovary showed Hodgkin's lymphoma with grade 1 nodular sclerosis (procedure)
C4030586|biopsy of ovary showed Hodgkin's lymphoma with grade 1 nodular sclerosis
C4030066|biopsy ovary malignant neoplasm mullerian mixed tumor (procedure)
C4030066|biopsy ovary malignant neoplasm mullerian mixed tumor
C4030068|biopsy ovary malignant neoplasm mesodermal mixed tumor (procedure)
C4030068|biopsy ovary malignant neoplasm mesodermal mixed tumor
C4030101|biopsy ovary malignant neoplasm carcinoid tumor neuroendocrine
C4030101|biopsy ovary malignant neoplasm carcinoid tumor neuroendocrine (procedure)
C4030182|biopsy ovary malignant adenocarcinoma villous (procedure)
C4030182|biopsy ovary malignant adenocarcinoma villous
C4030061|biopsy ovary malignant neoplasm myosarcoma leiomyosarcoma myxoid
C4030061|biopsy ovary malignant neoplasm myosarcoma leiomyosarcoma myxoid (procedure)
C4030056|biopsy ovary malignant neoplasm spindle cell type
C4030056|biopsy ovary malignant neoplasm spindle cell type (procedure)
C4030192|biopsy ovary malig lymphoma hodgkin's lymphocyt deplet diffuse fibrosis
C4030192|biopsy ovary malig lymphoma hodgkin's lymphocyt deplet diffuse fibrosis (procedure)
C4030190|biopsy ovary malig lymphoma hodgkin's nodular lymphocyte predominance (procedure)
C4030190|biopsy ovary malig lymphoma hodgkin's nodular lymphocyte predominance
C4030048|biopsy ovary malignant sarcoma epithelioid
C4030048|biopsy ovary malignant sarcoma epithelioid (procedure)
C4030123|biopsy ovary malignant lymphoma lymphoplasmacytic (procedure)
C4030123|biopsy ovary malignant lymphoma lymphoplasmacytic
C4030583|biopsy of ovary showed malignant neoplasm
C4030583|biopsy of ovary showed malignant neoplasm (procedure)
C4030204|biopsy ovary malig adenocarc metaplastic neuroendocrine differentiation (procedure)
C4030204|biopsy ovary malig adenocarc metaplastic neuroendocrine differentiation
C4030047|biopsy ovary malignant sarcoma follicular dendritic cell (procedure)
C4030047|biopsy ovary malignant sarcoma follicular dendritic cell
C4030092|biopsy ovary malignant neoplasm fibrosarcoma
C4030092|biopsy ovary malignant neoplasm fibrosarcoma (procedure)
C4030187|biopsy ovary malig lymphoma precursor cell lymphoblastic b-cell
C4030187|biopsy ovary malig lymphoma precursor cell lymphoblastic b-cell (procedure)
C4030105|biopsy ovary malignant neoplasm carcinoid tumor atypical
C4030105|biopsy ovary malignant neoplasm carcinoid tumor atypical (procedure)
C4030202|biopsy ovary malig adenocarcinoma endometrioid secretory variant (procedure)
C4030202|biopsy ovary malig adenocarcinoma endometrioid secretory variant
C4030042|biopsy ovary malignant sarcoma mast cell (procedure)
C4030042|biopsy ovary malignant sarcoma mast cell
C4030138|biopsy ovary malignant lymphoma composite hodgkin's and non-hodgkin's
C4030138|biopsy ovary malignant lymphoma composite hodgkin's and non-hodgkin's (procedure)
C4030108|biopsy ovary malignant neoplasm brenner tumor (procedure)
C4030108|biopsy ovary malignant neoplasm brenner tumor
C4030110|biopsy ovary malignant neoplasm adenocarcinofibroma serous
C4030110|biopsy ovary malignant neoplasm adenocarcinofibroma serous (procedure)
C4030106|biopsy ovary malignant neoplasm carcinoid tumor adenocarcinoid (procedure)
C4030106|biopsy ovary malignant neoplasm carcinoid tumor adenocarcinoid
C4030103|biopsy ovary malignant neoplasm carcinoid tumor enterochromaffin cell (procedure)
C4030103|biopsy ovary malignant neoplasm carcinoid tumor enterochromaffin cell
C4030057|biopsy ovary malignant neoplasm small cell type
C4030057|biopsy ovary malignant neoplasm small cell type (procedure)
C4030137|biopsy ovary malignant lymphoma follicular
C4030137|biopsy ovary malignant lymphoma follicular (procedure)
C4030128|biopsy ovary malignant lymphoma hodgkin's mixed cellularity
C4030128|biopsy ovary malignant lymphoma hodgkin's mixed cellularity (procedure)
C4030127|biopsy ovary malignant lymphoma hodgkin's nodular sclerosis
C4030127|biopsy ovary malignant lymphoma hodgkin's nodular sclerosis (procedure)
C4030125|biopsy ovary malignant lymphoma large b-cell diffuse (procedure)
C4030125|biopsy ovary malignant lymphoma large b-cell diffuse
C4030119|biopsy ovary malignant lymphoma mature t-cell angioimmunoblastic (procedure)
C4030119|biopsy ovary malignant lymphoma mature t-cell angioimmunoblastic
C4030203|biopsy ovary malig adenocarcinoma endometrioid ciliated cell variant
C4030203|biopsy ovary malig adenocarcinoma endometrioid ciliated cell variant (procedure)
C4030113|biopsy ovary malignant neoplasm adenocarcinofibroma
C4030113|biopsy ovary malignant neoplasm adenocarcinofibroma (procedure)
C4030063|biopsy ovary malignant neoplasm myosarcoma leiomyosarcoma (procedure)
C4030063|biopsy ovary malignant neoplasm myosarcoma leiomyosarcoma
C4030126|biopsy ovary malignant lymphoma hodgkin's sarcoma
C4030126|biopsy ovary malignant lymphoma hodgkin's sarcoma (procedure)
C4030089|biopsy ovary malignant neoplasm fibrosarcoma infantile
C4030089|biopsy ovary malignant neoplasm fibrosarcoma infantile (procedure)
C4030133|biopsy ovary malignant lymphoma histiocytosis
C4030133|biopsy ovary malignant lymphoma histiocytosis (procedure)
C4030131|biopsy ovary malignant lymphoma hodgkin's granuloma
C4030131|biopsy ovary malignant lymphoma hodgkin's granuloma (procedure)
C4030093|biopsy ovary malignant neoplasm epithelioid trophoblastic tumor (procedure)
C4030093|biopsy ovary malignant neoplasm epithelioid trophoblastic tumor
C4030584|biopsy of ovary showed malignant endometrioid adenofibroma (procedure)
C4030584|biopsy of ovary showed malignant endometrioid adenofibroma
C4030584|biopsy ovary malignant adenocarcinoma endometrioid adenofibroma
C4030050|biopsy ovary malignant neoplasm teratoma undifferentiated (procedure)
C4030050|biopsy ovary malignant neoplasm teratoma undifferentiated
C4030052|biopsy ovary malignant neoplasm teratoma mixed germ cell tumor (procedure)
C4030052|biopsy ovary malignant neoplasm teratoma mixed germ cell tumor
C4030596|biopsy of ovary showed adenocarcinoma with metaplasia
C4030596|biopsy of ovary showed adenocarcinoma with metaplasia (procedure)
C4030596|biopsy ovary malignant adenocarcinoma metaplastic
C4030181|biopsy ovary malignant carcinoma adenosquamous (procedure)
C4030181|biopsy ovary malignant carcinoma adenosquamous
C4030121|biopsy ovary malignant lymphoma marginal zone b-cell (procedure)
C4030121|biopsy ovary malignant lymphoma marginal zone b-cell
C4030585|biopsy of ovary showed Hodgkin's lymphoma with nodular sclerosis, cellular phase (procedure)
C4030585|biopsy of ovary showed Hodgkin's lymphoma with nodular sclerosis, cellular phase
C4030585|biopsy ovary malig lymphoma hodgkin's nodular sclerosis cellular phase
C4030053|biopsy ovary malignant neoplasm teratoma intermediate
C4030053|biopsy ovary malignant neoplasm teratoma intermediate (procedure)
C4030153|biopsy ovary malignant carcinoma squamous cell adenoid
C4030153|biopsy ovary malignant carcinoma squamous cell adenoid (procedure)
C4030107|biopsy ovary malignant neoplasm carcinoid tumor (procedure)
C4030107|biopsy ovary malignant neoplasm carcinoid tumor
C4030046|biopsy ovary malignant sarcoma giant cell (procedure)
C4030046|biopsy ovary malignant sarcoma giant cell
C4030041|biopsy ovary malignant sarcoma myxosarcoma (procedure)
C4030041|biopsy ovary malignant sarcoma myxosarcoma
C4030091|biopsy ovary malignant neoplasm fibrosarcoma fascial
C4030091|biopsy ovary malignant neoplasm fibrosarcoma fascial (procedure)
C4030188|biopsy ovary malig lymphoma mixed small and large cell, diffuse
C4030188|biopsy ovary malig lymphoma mixed small and large cell, diffuse (procedure)
C4030130|biopsy ovary malignant lymphoma hodgkin's lymphocyte-rich
C4030130|biopsy ovary malignant lymphoma hodgkin's lymphocyte-rich (procedure)
C4030124|biopsy ovary malignant lymphoma large b-cell diffuse immunoblastic
C4030124|biopsy ovary malignant lymphoma large b-cell diffuse immunoblastic (procedure)
C4030070|biopsy ovary malignant neoplasm lymphoma
C4030070|biopsy ovary malignant neoplasm lymphoma (procedure)
C4030067|biopsy ovary malignant neoplasm mesonephroma (procedure)
C4030067|biopsy ovary malignant neoplasm mesonephroma
C4030098|biopsy ovary malignant neoplasm carcinosarcoma embryonal (procedure)
C4030098|biopsy ovary malignant neoplasm carcinosarcoma embryonal
C4030159|biopsy ovary malignant carcinoma signet ring cell (procedure)
C4030159|biopsy ovary malignant carcinoma signet ring cell
C4030200|biopsy ovary malig carcinoid tumor enterochromaffin-like cell
C4030200|biopsy ovary malig carcinoid tumor enterochromaffin-like cell (procedure)
C4030082|biopsy ovary malignant neoplasm giant cell type
C4030082|biopsy ovary malignant neoplasm giant cell type (procedure)
C4030136|biopsy ovary malignant lymphoma follicular grade 1
C4030136|biopsy ovary malignant lymphoma follicular grade 1 (procedure)
C4030055|biopsy ovary malignant neoplasm struma ovarii (procedure)
C4030055|biopsy ovary malignant neoplasm struma ovarii
C4030196|biopsy ovary malig choriocarcinoma combined w/ other germ cell elements
C4030196|biopsy ovary malig choriocarcinoma combined w/ other germ cell elements (procedure)
C0022790|Krukenberg Tumor
C0022790|Krukenbergs Tumor
C0022790|Tumor, Krukenberg's
C0022790|Tumor, Krukenberg
C0022790|Krukenberg tumour
C0022790|Krukenburg tumour
C0022790|Krukenburg tumor
C0022790|Krukenberg tumor (disorder)
C0022790|Krukenburg tumor (disorder)
C0022790|signet ring cell adenocarcinoma metastatic to ovary (diagnosis)
C0022790|signet ring cell adenocarcinoma metastatic to ovary
C0022790|metastatic carcinoma to the ovary (Krukenberg tumor)
C0022790|Carcinoma, Krukenberg
C0022790|Krukenberg Tumor [Disease/Finding]
C0022790|Krukenberg's Tumor
C0022790|Krukenberg Carcinoma
C0022790|Cancer metastatic to ovary
C0022790|Secondary malignant neoplasm of ovary
C0022790|Metastasis to ovary
C0022790|Ovarian metastasis
C0022790|Secondary tumor to ovary
C0022790|Secondary tumour to ovary
C0022790|Secondary cancer of ovary
C0022790|Metastatic malignant neoplasm to ovary
C0022790|Secondary malignant neoplasm of ovary (disorder)
C0022790|Krukenberg; tumor
C0022790|tumor; Krukenberg
C0022790|Krukenberg Neoplasm
C1386260|endometrioid; adenocarcinoma, unspecified site, female
C1386260|adenocarcinoma; endometrioid, unspecified site, female
C1386284|adenocarcinoma; papillary, serous, unspecified site
C1386284|adenocarcinoma; serous papillary, unspecified site
C1386284|papillary; adenocarcinoma, serous, unspecified site
C1386284|serous; adenocarcinoma, papillary, unspecified site
C1386285|adenocarcinoma; papillocystic, unspecified site
C1386285|papillocystic; adenocarcinoma, unspecified site
C1386286|adenocarcinoma; pseudomucinous, unspecified site
C1386286|pseudomucinous; adenocarcinoma, unspecified site
C0334341|Endometrioid adenofibroma, malignant
C0334341|Endometrioid cystadenofibroma, malignant
C0334341|Malignant endometrioid adenofibroma
C0334341|Malignant endometrioid cystadenofibroma
C0334341|Endometrioid adenofibroma, malignant (morphologic abnormality)
C0334341|cystadenofibroma; endometrioid, malignant
C0334341|endometrioid; adenofibroma, malignant
C0334341|endometrioid; cystadenofibroma, malignant
C0334341|adenofibroma; endometrioid, malignant
C1388418|malignant; androblastoma, unspecified site, female
C1388418|malignant; arrhenoblastoma, unspecified site, female
C1388418|androblastoma; malignant, unspecified site, female
C1388418|arrhenoblastoma; malignant, unspecified site, female
C1390413|borderline malignancy; mucinous cystadenoma, unspecified site
C1390413|cystadenoma; mucinous, borderline malignancy, unspecified site
C1390413|mucinous; cystadenoma, borderline malignancy, unspecified site
C0851188|borderline malignancy; mucinous cystadenoma, ovary
C0851188|cystadenoma; mucinous, borderline malignancy, ovary
C0851188|mucinous; cystadenoma, borderline malignancy, ovary
C0851188|ovary; cystadenoma, mucinous, borderline malignancy
C0851188|ovary; mucinous cystadenoma, borderline malignancy
C1390414|borderline malignancy; mucinous papillary cystadenoma, unspecified site
C1390414|borderline malignancy; papillary mucinous cystadenoma, unspecified site
C1390414|cystadenoma; mucinous, papillary, borderline malignancy, unspecified site
C1390414|cystadenoma; papillary, mucinous, borderline malignancy, unspecified site
C1390414|mucinous; cystadenoma, papillary, borderline malignancy, unspecified site
C1390414|papillary; cystadenoma, mucinous, borderline malignancy, unspecified site
C0851177|papillary mucinous cystadenoma of ovary of borderline malignancy (diagnosis)
C0851177|papillary mucinous cystadenoma of ovary of borderline malignancy
C0851177|papillary mucinous ovarian cystadenoma of borderline malignancy
C0851177|borderline malignancy; mucinous papillary cystadenoma, ovary
C0851177|borderline malignancy; papillary mucinous cystadenoma, ovary
C0851177|cystadenoma; mucinous, papillary, borderline malignancy, ovary
C0851177|cystadenoma; papillary, mucinous, borderline malignancy, ovary
C0851177|mucinous; cystadenoma, papillary, borderline malignancy, ovary
C0851177|ovary; cystadenoma, mucinous papillary, borderline malignancy
C0851177|ovary; cystadenoma, papillary mucinous, borderline malignancy
C0851177|ovary; mucinous papillary cystadenoma, borderline malignancy
C0851177|ovary; papillary mucinous cystadenoma, borderline malignancy
C0851177|papillary; cystadenoma, mucinous, borderline malignancy, ovary
C0334356|Papillary cystadenoma, borderline malignancy -RETIRED-
C0334356|Papillary cystadenoma - borderline malignancy
C0334356|Papillary cystadenoma - borderline malignancy (disorder)
C0334356|Papillary cystadenoma, borderline malignancy
C0334356|Papillary cystadenoma, borderline malignancy (morphologic abnormality)
C0334356|[M] Papillary cystadenoma, borderline malignancy
C0334356|[M]Papillary cystadenoma, borderline malignancy
C0334356|borderline malignancy; papillary cystadenoma, unspecified site
C0334356|cystadenoma; papillary, borderline malignancy, unspecified site
C0334356|papillary; cystadenoma, borderline malignancy, unspecified site
C0334356|Low Malignancy Potential Papillary Cystadenoma
C0334356|Borderline Malignancy Papillary Cystadenoma
C0334356|Borderline Papillary Cystadenoma
C0851186|papillary cystadenoma of ovary of borderline malignancy (diagnosis)
C0851186|papillary cystadenoma of ovary of borderline malignancy
C0851186|papillary ovarian cystadenoma of borderline malignancy
C0851186|borderline malignancy; papillary cystadenoma, ovary
C0851186|cystadenoma; papillary, borderline malignancy, ovary
C0851186|ovary; cystadenoma, papillary, borderline malignancy
C0851186|ovary; papillary cystadenoma, borderline malignancy
C0851186|papillary; cystadenoma, borderline malignancy, ovary
C1390415|borderline malignancy; papillary pseudomucinous cystadenoma, unspecified site
C1390415|borderline malignancy; pseudomucinous papillary cystadenoma, unspecified site
C1390415|cystadenoma; papillary, pseudomucinous, borderline malignancy, unspecified site
C1390415|cystadenoma; pseudomucinous, papillary, borderline malignancy, unspecified site
C1390415|papillary; cystadenoma, pseudomucinous, borderline malignancy, unspecified site
C1390415|pseudomucinous; cystadenoma, papillary, borderline malignancy, unspecified site
C1390416|borderline malignancy; papillary pseudomucinous cystadenoma, ovary
C1390416|borderline malignancy; pseudomucinous papillary cystadenoma, ovary
C1390416|cystadenoma; papillary, pseudomucinous, borderline malignancy, ovary
C1390416|cystadenoma; pseudomucinous, papillary, borderline malignancy, ovary
C1390416|ovary; cystadenoma, papillary pseudomucinous, borderline malignancy
C1390416|ovary; cystadenoma, pseudomucinous papillary, borderline malignancy
C1390416|ovary; papillary pseudomucinous cystadenoma, borderline malignancy
C1390416|ovary; pseudomucinous papillary cystadenoma, borderline malignancy
C1390416|papillary; cystadenoma, pseudomucinous, borderline malignancy, ovary
C1390416|pseudomucinous; cystadenoma, papillary, borderline malignancy, ovary
C1390417|borderline malignancy; papillary serous cystadenoma, unspecified site
C1390417|borderline malignancy; serous papillary cystadenoma, unspecified site
C1390417|cystadenoma; papillary, serous, borderline malignancy, unspecified site
C1390417|cystadenoma; serous, papillary, borderline malignancy, unspecified site
C1390417|papillary; cystadenoma, serous, borderline malignancy, unspecified site
C1390417|serous; cystadenoma, papillary, borderline malignancy, unspecified site
C0851187|borderline malignancy; papillary serous cystadenoma, ovary
C0851187|borderline malignancy; serous papillary cystadenoma, ovary
C0851187|cystadenoma; papillary, serous, borderline malignancy, ovary
C0851187|cystadenoma; serous, papillary, borderline malignancy, ovary
C0851187|ovary; cystadenoma, papillary serous, borderline malignancy
C0851187|ovary; cystadenoma, serous papillary, borderline malignancy
C0851187|ovary; papillary serous cystadenoma, borderline malignancy
C0851187|ovary; serous papillary cystadenoma, borderline malignancy
C0851187|papillary; cystadenoma, serous, borderline malignancy, ovary
C0851187|serous; cystadenoma, papillary, borderline malignancy, ovary
C1390418|borderline malignancy; pseudomucinous cystadenoma, unspecified site
C1390418|cystadenoma; pseudomucinous, borderline malignancy, unspecified site
C1390418|pseudomucinous; cystadenoma, borderline malignancy, unspecified site
C1390419|borderline malignancy; pseudomucinous cystadenoma, ovary
C1390419|cystadenoma; pseudomucinous, borderline malignancy, ovary
C1390419|ovary; cystadenoma, pseudomucinous, borderline malignancy
C1390419|ovary; pseudomucinous cystadenoma, borderline malignancy
C1390419|pseudomucinous; cystadenoma, borderline malignancy, ovary
C1390420|borderline malignancy; serous cystadenoma, unspecified site
C1390420|cystadenoma; serous, borderline malignancy, unspecified site
C1390420|serous; cystadenoma, borderline malignancy, unspecified site
C0851185|serous cystadenoma of borderline malignancy of ovary
C0851185|serous cystadenoma of borderline malignancy of ovary (diagnosis)
C0851185|serous ovarian cystadenoma of borderline malignancy
C0851185|borderline malignancy; serous cystadenoma, ovary
C0851185|cystadenoma; serous, borderline malignancy, ovary
C0851185|ovary; cystadenoma, serous, borderline malignancy
C0851185|ovary; serous cystadenoma, borderline malignancy
C0851185|serous; cystadenoma, borderline malignancy, ovary
C0206687|Carcinoma, Endometrioid
C0206687|Carcinomas, Endometrioid
C0206687|Endometrioid Carcinomas
C0206687|Endometrioid Carcinoma
C0206687|endometrioid carcinoma (diagnosis)
C0206687|Carcinoma, Endometrioid [Disease/Finding]
C0206687|Endometrioid Adenocarcinoma
C0206687|Endometrioid carcinoma (morphologic abnormality)
C0206687|carcinoma; endometrioid, unspecified site, female
C0206687|endometrioid; carcinoma, unspecified site, female
C0206687|Endometrioid Carcinoma of Female Reproductive System
C0206687|Endometrioid Carcinoma of the Female Reproductive System
C0206687|Female Reproductive Endometrioid Carcinoma
C0334401|Malignant Granulosa Cell Tumor
C0334401|GRANULOSA CELL TUMOR, MALIGNANT
C0334401|Granulosa cell carcinoma
C0334401|Malignant granulosa cell tumour
C0334401|Granulosa cell tumour, malignant
C0334401|Granulosa cell tumor, malignant (morphologic abnormality)
C0334401|Granulosa cell tumor, sarcomatoid
C0334401|Granulosa cell tumour, sarcomatoid
C0334401|carcinoma; granulosa cell
C0334401|granulosa cell; carcinoma
C0334401|granulosa cell; tumor, malignant
C0334401|tumor; granulosa cell, malignant
C0334401|Malignant Granulosa Cell Neoplasm
C1391921|carcinoma; Leydig cell, unspecified site, female
C1391921|Leydig cell; carcinoma, unspecified site, female
C1391935|carcinoma; papillary, serous, unspecified site
C1391935|carcinoma; serous, papillary, unspecified site
C1391935|papillary; carcinoma, serous, unspecified site
C1391935|serous; carcinoma, papillary, unspecified site
C1391936|carcinoma; papillary, serous, superficial, unspecified site
C1391936|carcinoma; serous, superficial, papillary, unspecified site
C1391936|papillary; carcinoma, serous, superficial, unspecified site
C1391936|serous; carcinoma, superficial, papillary, unspecified site
C1391937|carcinoma; papillocystic, unspecified site
C1391937|papillocystic; carcinoma, unspecified site
C1391941|carcinoma; pseudomucinous, unspecified site
C1391941|pseudomucinous; carcinoma, unspecified site
C1391945|carcinoma; Sertoli cell, unspecified site, female
C1391945|Sertoli cell; carcinoma, unspecified site, female
C0728814|[M]Theca cell carcinoma (morphologic abnormality)
C0728814|[M]Theca cell carcinoma
C0728814|carcinoma; theca cell
C0728814|theca cell; carcinoma
C1394299|cystadenocarcinoma; endometrioid, unspecified site, female
C1394299|endometrioid; cystadenocarcinoma, unspecified site, female
C0206699|Cystadenocarcinoma, Mucinous
C0206699|Cystadenocarcinomas, Mucinous
C0206699|Mucinous Cystadenocarcinomas
C0206699|Mucinous Cystadenocarcinoma
C0206699|Cystadenocarcinoma, Mucinous [Disease/Finding]
C0206699|[M]Mucinous cystadenocarcinoma NOS
C0206699|[M]Mucinous cystadenocarcinoma NOS (morphologic abnormality)
C0206699|Pseudomucinous adenocarcinoma
C0206699|Pseudomucinous cystadenocarcinoma
C0206699|Mucinous cystadenocarcinoma (morphologic abnormality)
C0206699|cystadenocarcinoma; mucinous, unspecified site
C0206699|cystadenocarcinoma; pseudomucinous, unspecified site
C0206699|mucinous; cystadenocarcinoma, unspecified site
C0206699|pseudomucinous; cystadenocarcinoma, unspecified site
C0206699|Mucinous cystadenocarcinoma, NOS
C0206699|Pseudomucinous cystadenocarcinoma, NOS
C0334364|Papillary Mucinous Cystadenocarcinoma
C0334364|Papillary pseudomucinous adenocarcinoma
C0334364|Papillary pseudomucinous cystadenocarcinoma
C0334364|Papillary mucinous cystadenocarcinoma (morphologic abnormality)
C0334364|cystadenocarcinoma; mucinous, papillary, unspecified site
C0334364|cystadenocarcinoma; papillary, mucinous, unspecified site
C0334364|mucinous; cystadenocarcinoma, papillary, unspecified site
C0334364|papillary; cystadenocarcinoma, mucinous, unspecified site
C0206700|Cystadenocarcinoma, Papillary
C0206700|Cystadenocarcinomas, Papillary
C0206700|Papillary Cystadenocarcinomas
C0206700|Papillary Cystadenocarcinoma
C0206700|Cystadenocarcinoma, Papillary [Disease/Finding]
C0206700|[M]Papillary cystadenocarcinoma, NOS (morphologic abnormality)
C0206700|[M]Papillary cystadenocarcinoma, NOS
C0206700|CYSTADENOCARCINOMA, PAPILLARY, MALIGNANT
C0206700|Papillocystic adenocarcinoma
C0206700|Papillary cystadenocarcinoma (morphologic abnormality)
C0206700|cystadenocarcinoma; papillary, unspecified site
C0206700|papillary; cystadenocarcinoma, unspecified site
C0206700|Papillary cystadenocarcinoma, NOS
C1394300|cystadenocarcinoma; papillary, pseudomucinous, unspecified site
C1394300|cystadenocarcinoma; pseudomucinous, papillary, unspecified site
C1394300|papillary; cystadenocarcinoma, pseudomucinous, unspecified site
C1394300|pseudomucinous; cystadenocarcinoma, papillary, unspecified site
C1394301|cystadenocarcinoma; papillary, serous, unspecified site
C1394301|cystadenocarcinoma; serous, papillary, unspecified site
C1394301|papillary; cystadenocarcinoma, serous, unspecified site
C1394301|serous; cystadenocarcinoma, papillary, unspecified site
C1394302|cystadenocarcinoma; serous, unspecified site
C1394302|serous; cystadenocarcinoma, unspecified site
C0334523|teratoma with malignant transformation (diagnosis)
C0334523|teratoma with malignant transformation
C0334523|Teratoma with malignant transformation (morphologic abnormality)
C0334523|Dermoid cyst with malignant transformation
C0334523|Dermoid cyst with malignant transformation (morphologic abnormality)
C0334523|Dermoid cyst with secondary tumor
C0334523|Dermoid cyst with secondary tumour
C0334523|dermoid; cyst, with malignant transformation
C0334523|malignant; transformation dermoid cyst
C0334523|Teratoma with malignant transformation [dup] (morphologic abnormality)
C0334523|:: Dermoid cyst with malignant transformation
C1395294|dermoid; tumor, with malignant transformation
C1395294|malignant; transformation dermoid tumor
C1395294|tumor; dermoid, with malignant transformation
C1395294|transformation; malignant, in dermoid tumor
C1395771|tumor; yolk sac, unspecified site, female
C1395771|yolk sac; tumor, unspecified site, female
C1395937|dysgerminoma; unspecified site, female
C1396616|endodermal; sinus, tumor, unspecified site, female
C1396616|tumor; endodermal sinus, unspecified site, female
C1402882|Leydig cell; tumor, malignant, unspecified site, female
C1402882|tumor; Leydig cell, malignant, unspecified site, female
C1403527|malignant; transformation dermoid
C1334811|mucinous; tumor, unspecified site
C1334811|tumor; mucinous, unspecified site
C1334811|Mucinous Neoplasm
C1334811|Mucinous Tumor
C1408999|ovarii; goiter, malignant
C1406886|ovary; teratoma, embryonal, immature or malignant
C1406886|teratoma; ovary, embryonal, immature or malignant
C1407806|papillary; tumor, mucinous, unspecified site
C1407806|tumor; papillary mucinous, unspecified site
C0334366|Papillary mucinous cystadenoma, borderline malignancy -RETIRED-
C0334366|Papillary mucinous cystadenoma, borderline malignancy
C0334366|Papillary mucinous cystadenoma, borderline malignancy (morphologic abnormality)
C0334366|Papillary mucinous cystadenoma - borderline malignancy
C0334366|Papillary mucinous tumor of low malignant potential
C0334366|Papillary mucinous tumour of low malignant potential
C0334366|Papillary pseudomucinous cystadenoma, borderline malignancy
C0334366|papillary; tumor, mucinous, of low malignant potential
C0334366|tumor; papillary, mucinous, of low malignant potential
C0334366|Low Malignancy Potential Papillary Mucinous Cystadenoma
C0334366|Low Malignancy Potential Papillary Pseudomucinous Cystadenoma
C0334366|Papillary Mucinous Neoplasm of Low Malignant Potential
C0334366|Borderline Malignancy Papillary Mucinous Cystadenoma
C0334366|Borderline Malignancy Papillary Pseudomucinous Cystadenoma
C0334366|Borderline Papillary Mucinous Cystadenoma
C0334366|Borderline Papillary Pseudomucinous Cystadenoma
C1407807|papillary; tumor, serous, low malignant potential, unspecified site
C1407807|tumor; papillary serous, low malignant potential, unspecified site
C1405367|polyvesicular; tumor, unspecified site, female
C1405367|tumor; polyvesicular, unspecified site, female
C1407812|serous; tumor, unspecified site
C1407812|tumor; serous, unspecified site
C1518236|Malignant Ovarian Surface Epithelial-Stromal Tumor
C1518236|Ovarian stromal cancer
C1518236|Malignant Ovarian Epithelial Tumor
C1518236|cancer, ovarian stromal
C1518236|stromal cancer, ovarian
C1518236|Malignant Ovarian Surface Epithelial-Stromal Neoplasm
C1518721|Ovarian Malignant Mesothelioma
C1335169|Ovarian Müllerian Adenosarcoma
C1335169|Ovarian Mesodermal Adenosarcoma
C1335169|Ovarian Adenosarcoma
C1518720|Primary Ovarian Lymphoma
C1518720|Ovarian Lymphoma
C0235770|Malignant ovarian cyst
C0235770|Ovarian cyst malignant
C1334609|Malignant Ovarian Sex Cord-Stromal Neoplasm
C1334609|Malignant Ovarian Sex Cord-Stromal Tumor
C1334609|Malignant Sex Cord-Stromal Tumor of Ovary
C1334609|Malignant Sex Cord-Stromal Tumor of the Ovary
C1518746|Ovarian Wilms' Tumor
C1518746|Ovarian Wilms Tumor
C1827462|Carcinoma of ovary, stage 2 (finding)
C1827462|Carcinoma of ovary, stage 2
C1827462|Ovarian cancer stage 2
C1827462|Cancer of ovary, stage 2
C0346162|serous papillary cystadenocarcinoma of ovary
C0346162|serous papillary cystadenocarcinoma of ovary (diagnosis)
C0346162|Serous papillary cystadenocarcinoma ovary
C0346162|Serous papillary cystadenocarcinoma ovary (disorder)
C0279665|mucinous cystadenocarcinoma of ovary
C0279665|mucinous cystadenocarcinoma of ovary (diagnosis)
C0279665|Mucinous cystadenocarcinoma ovary
C0279665|Mucinous cystadenocarcinoma of ovary (disorder)
C0279665|ovarian mucinous cystadenocarcinoma
C0279665|cystadenocarcinoma of the ovary, mucinous
C0279665|cystadenocarcinoma, mucinous, ovarian
C0279665|cystadenocarcinoma, ovarian mucinous
C0279665|mucinous cystadenocarcinoma of the ovary
C0279665|ovarian cancer, mucinous cystadenocarcinoma
C0279665|ovary cancer, mucinous cystadenocarcinoma
C0521156|Epithelial ovarian tumor, International Federation of Gynecology and Obstetrics stage IV (finding)
C0521156|Epithelial ovarian tumor, FIGO stage IV (finding)
C0521156|Epithelial ovarian tumor, International Federation of Gynecology and Obstetrics stage IV
C0521156|Epithelial ovarian tumour, International Federation of Gynecology and Obstetrics stage IV
C0521156|Epithelial ovarian tumor, FIGO stage IV
C0521156|Epithelial ovarian tumour, FIGO stage IV
C0521156|Epithelial ovarian tumor, FIGO stage IV (tumor staging)
C1096638|cystadenocarcinoma of ovary (diagnosis)
C1096638|cystadenocarcinoma of ovary
C1096638|Cystadenocarcinoma ovary
C1096638|Cystadenocarcinoma of ovary (disorder)
C1096638|Cystadenocarcinoma of the Ovary
C1096638|Ovarian Cystadenocarcinoma
C0346174|ovarian neoplasm malignant gonadal stromal tumor sex cord
C0346174|malignant sex cord tumor of ovary
C0346174|malignant sex cord tumor of ovary (diagnosis)
C0346174|Malignant sex cord tumour of ovary
C0346174|Malignant sex cord tumor of ovary (disorder)
C1827620|Carcinoma of ovary, stage 4
C1827620|Carcinoma of ovary, stage 4 (finding)
C1827620|Ovarian cancer stage 4
C1827620|Cancer of ovary, stage 4
C0346183|embryonal carcinoma of ovary
C0346183|embryonal carcinoma of ovary (diagnosis)
C0346183|Ovarian embryonal carcinoma
C0346183|Embryonal carcinoma of ovary (disorder)
C0346183|Embryonal Carcinoma of the Ovary
C0521152|Epithelial ovarian tumor, International Federation of Gynecology and Obstetrics stage IIA (finding)
C0521152|Epithelial ovarian tumor, FIGO stage IIA (finding)
C0521152|Epithelial ovarian tumor, International Federation of Gynecology and Obstetrics stage IIA
C0521152|Epithelial ovarian tumour, International Federation of Gynaecology and Obstetrics stage IIA
C0521152|Epithelial ovarian tumor, FIGO stage IIA
C0521152|Epithelial ovarian tumour, FIGO stage IIA
C0521152|Epithelial ovarian tumor, FIGO stage IIA (tumor staging)
C1562619|Malignant mesonephroid tumor of ovary
C1562619|Malignant mesonephroid tumour of ovary
C1562619|Primary malignant clear cell tumor of ovary (disorder)
C1562619|Primary malignant clear cell tumor of ovary
C1562619|Primary malignant clear cell tumour of ovary
C0521154|Epithelial ovarian tumor, International Federation of Gynecology and Obstetrics stage IIC
C0521154|Epithelial ovarian tumor, International Federation of Gynecology and Obstetrics stage IIC (finding)
C0521154|Epithelial ovarian tumor, FIGO stage IIC (finding)
C0521154|Epithelial ovarian tumour, International Federation of Gynecology and Obstetrics stage IIC
C0521154|Epithelial ovarian tumor, FIGO stage IIC
C0521154|Epithelial ovarian tumour, FIGO stage IIC
C0521154|Epithelial ovarian tumor, FIGO stage IIC (tumor staging)
C0346166|ovarian neoplasm epithelial mixed
C0346166|mixed epithelial neoplasm of ovary
C0346166|mixed epithelial neoplasm of ovary (diagnosis)
C0346166|Mixed epithelial tumor of ovary
C0346166|Mixed epithelial tumour of ovary
C0346166|Mixed epithelial tumor of ovary (disorder)
C0346166|Mixed Epithelial Neoplasm of the Ovary
C0346166|Mixed Epithelial Tumor of the Ovary
C0346166|Ovarian Mixed Epithelial Neoplasm
C0346166|Ovarian Mixed Epithelial Tumor
C1297996|Primary malignant neoplasm of right ovary (diagnosis)
C1297996|Primary malignant neoplasm of right ovary
C1297996|ovarian malignant neoplasm primary right
C1297996|Primary malignant neoplasm of right ovary (disorder)
C2016048|mixed cellularity Hodgkin's lymphoma of ovary (diagnosis)
C2016048|mixed cellularity Hodgkin's lymphoma of ovary
C2046511|ovarian malignant lymphoma Hodgkin's and non-Hodgkin's
C2046511|composite Hodgkin's and non-Hodgkin's lymphoma of ovary (diagnosis)
C2046511|composite Hodgkin's and non-Hodgkin's lymphoma of ovary
C2016073|mantle cell lymphoma of ovary (diagnosis)
C2016073|mantle cell lymphoma of ovary
C2016078|NK/T-cell lymphoma of ovary (diagnosis)
C2016078|NK/T-cell lymphoma of ovary
C2212025|Sezary syndrome of ovary (diagnosis)
C2212025|Sezary syndrome of ovary
C2016046|ovarian Hodgkin lymphoma lymphocytic depletion diffuse fibrosis
C2016046|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of ovary
C2016046|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of ovary (diagnosis)
C2016049|lymphocyte-rich nodular Hodgkin's lymphoma of ovary (diagnosis)
C2016049|lymphocyte-rich nodular Hodgkin's lymphoma of ovary
C2016077|mixed small and large cell diffuse lymphoma of ovary (diagnosis)
C2016077|mixed small and large cell diffuse lymphoma of ovary
C2016071|immunoblastic large B-cell diffuse lymphoma of ovary (diagnosis)
C2016071|immunoblastic large B-cell diffuse lymphoma of ovary
C2016068|grade 3 follicular lymphoma of ovary (diagnosis)
C2016068|grade 3 follicular lymphoma of ovary
C2016070|large B-cell diffuse lymphoma of ovary (diagnosis)
C2016070|large B-cell diffuse lymphoma of ovary
C2016076|angioimmunoblastic T-cell lymphoma of ovary (diagnosis)
C2016076|angioimmunoblastic T-cell lymphoma of ovary
C2016076|angioimmunoblastic lymphadenopathy with dysproteinemia (AILD) of ovary
C2016044|lymphocyte-rich Hodgkin's lymphoma of ovary
C2016044|lymphocyte-rich Hodgkin's lymphoma of ovary (diagnosis)
C2016047|Hodgkin's disease, lymphocytic depletion, reticular of ovary
C2016047|Hodgkin's disease, lymphocytic depletion, reticular of ovary (diagnosis)
C2113645|precursor B-cell lymphoblastic lymphoma of ovary (diagnosis)
C2113645|precursor B-cell lymphoblastic lymphoma of ovary
C2212035|mast cell sarcoma of ovary (diagnosis)
C2212035|mast cell sarcoma of ovary
C2016067|grade 2 follicular lymphoma of ovary (diagnosis)
C2016067|grade 2 follicular lymphoma of ovary
C2016050|nodular sclerosing Hodgkin's lymphoma of ovary (diagnosis)
C2016050|nodular sclerosing Hodgkin's lymphoma of ovary
C2046584|Hodgkin's granuloma of ovary
C2046584|Hodgkin's granuloma of ovary (diagnosis)
C2016066|grade 1 follicular lymphoma of ovary
C2016066|grade 1 follicular lymphoma of ovary (diagnosis)
C2016075|mature T-cell lymphoma of ovary
C2016075|mature T-cell lymphoma of ovary (diagnosis)
C2113785|precursor T-cell lymphoblastic lymphoma of ovary
C2113785|precursor T-cell lymphoblastic lymphoma of ovary (diagnosis)
C2016045|Hodgkin's disease, lymphocytic depletion of ovary (diagnosis)
C2016045|Hodgkin's disease, lymphocytic depletion of ovary
C2016052|grade 1 nodular sclerosing Hodgkin's lymphoma of ovary
C2016052|grade 1 nodular sclerosing Hodgkin's lymphoma of ovary (diagnosis)
C2016053|grade 2 nodular sclerosing Hodgkin's lymphoma of ovary
C2016053|grade 2 nodular sclerosing Hodgkin's lymphoma of ovary (diagnosis)
C2016079|small B-cell lymphocytic lymphoma of ovary (diagnosis)
C2016079|small B-cell lymphocytic lymphoma of ovary
C2016074|marginal zone B-cell lymphoma of ovary (diagnosis)
C2016074|marginal zone B-cell lymphoma of ovary
C2113716|precursor cell lymphoblastic lymphoma of ovary (diagnosis)
C2113716|precursor cell lymphoblastic lymphoma of ovary
C2016051|nodular sclerosing Hodgkin's lymphoma in cellular phase of ovary (diagnosis)
C2016051|nodular sclerosing Hodgkin's lymphoma in cellular phase of ovary
C2046724|Hodgkin's sarcoma of ovary (diagnosis)
C2046724|Hodgkin's sarcoma of ovary
C2016072|lymphoplasmacytic lymphoma of ovary (diagnosis)
C2016072|lymphoplasmacytic lymphoma of ovary
C2016069|malignant histiocytosis of ovary
C2016069|malignant histiocytosis of ovary (diagnosis)
C0302592|CARCINOMA OF CERVIX
C0302592|Ca cervix
C0302592|Cervical carcinoma
C0302592|carcinoma of cervix (diagnosis)
C0302592|Carcinoma uterine cerix
C0302592|Carcinoma;cervix
C0302592|Ca cervix uteri NOS (disorder)
C0302592|Cancer of cervix
C0302592|Cervical carcinoma (uterus)
C0302592|Carcinoma cervix uteri
C0302592|Ca cervix uteri NOS
C0302592|cervical cancer
C0302592|Cervical cancer, NOS
C0302592|Cervix uteri cancer
C0302592|Cervical carcinoma NOS
C0302592|Cervix carcinoma
C0302592|Carcinoma cervix
C0302592|Carcinoma uterine cervix
C0302592|Carcinoma of cervix (disorder)
C0302592|Cancer of the Cervix
C0302592|Cervix Cancer
C0302592|Uterine Cervix Cancer
C0302592|Uterine Cervix Carcinoma
C0302592|Cancer of Uterine Cervix
C0302592|Cancer of the Uterine Cervix
C0302592|Carcinoma of Cervix Uteri
C0302592|Carcinoma of Uterine Cervix
C0302592|Carcinoma of the Cervix Uteri
C0302592|Carcinoma of the Cervix
C0302592|Carcinoma of the Uterine Cervix
C0302592|Cervix Uteri Carcinoma
C4048328|cervix cancer
C4048328|cervical cancer
C4048328|Cancer of cervix
C4048328|cervical cancer (diagnosis)
C4048328|Cancers, Cervix
C4048328|Cancer, Cervix
C4048328|Cervix uteri--Cancer
C4048328|Ca cervix
C4048328|Cancer of the Uterine Cervix
C4048328|Cancer of the Cervix
C4048328|Uterine Cervical Cancer
C4048328|uterine cervix cancer
C4048328|Cancer, Uterine Cervical
C4048328|Cancers, Uterine Cervical
C4048328|Cervical Cancer, Uterine
C4048328|Cervical Cancers, Uterine
C4048328|Uterine Cervical Cancers
C0279888|cellular diagnosis, cervical cancer
C0279888|cervical cancer cellular diagnosis
C0280232|stage, cervical cancer
C0280232|cervical cancer stage
C1280511|Primary malignant neoplasm of uterine cervix
C1280511|Primary malignant neoplasm of uterine cervix (disorder)
C4048331|Cancer of bronchus; lung
C0153615|Urachus
C0153615|Malignant neoplasm of urachus
C0153615|malignant neoplasm of urachus (diagnosis)
C0153615|malignant tumor of urachus
C0153615|Malig neo urachus
C0153615|Malignant tumour of urachus
C0153615|Malignant tumor of urachus (disorder)
C0153611|Malignant neoplasm of anterior wall of urinary bladder
C0153611|Anterior wall of bladder
C0153611|Malignant neoplasm of anterior wall of bladder
C0153611|malignant neoplasm of anterior wall of bladder (diagnosis)
C0153611|malignant tumor of anterior wall of bladder
C0153611|Mal neo bladder-anterior
C0153611|Malignant neoplasm of anterior wall of urinary bladder (disorder)
C0153613|Malignant neoplasm of bladder neck
C0153613|Bladder neck
C0153613|Malignant neoplasm of urinary bladder neck
C0153613|malignant neoplasm of neck of bladder
C0153613|malignant neoplasm of neck of bladder (diagnosis)
C0153613|malignant tumor of neck of bladder
C0153613|Mal neo bladder neck
C0153613|Malignant tumor of bladder neck
C0153613|Malignant tumour of bladder neck
C0153613|Malignant tumor of bladder neck (disorder)
C0005684|Malignant neoplasm of bladder
C0005684|Bladder, unspecified
C0005684|Malignant neoplasm of bladder, unspecified
C0005684|Cancer, Urinary Bladder
C0005684|BLADDER CANCER
C0005684|malignant neoplasm of bladder (diagnosis)
C0005684|bladder cancer (diagnosis)
C0005684|Ca bladder
C0005684|Bladder Cancers
C0005684|malignant tumor of bladder
C0005684|Malig neo bladder NOS
C0005684|Cancer of bladder
C0005684|Cancer, Bladder
C0005684|Bladder neoplasms malignant
C0005684|Urinary Bladder Cancer
C0005684|Malignant tumour of urinary bladder
C0005684|Malignant tumor of urinary bladder (disorder)
C0005684|Bladder Ca
C0005684|CA - Bladder cancer
C0005684|Malignant tumor of urinary bladder
C0005684|Malignant neoplasm of urinary bladder NOS
C0005684|Malignant neoplasm of urinary bladder NOS (disorder)
C0005684|Malignant neoplasm of urinary bladder
C0005684|Bladder--Cancer
C0005684|Bladder cancer NOS
C0005684|Malignant neoplasm of bladder, part unspecified
C0005684|Cancer of the Bladder
C0005684|Malignant neoplasm of bladder, NOS
C0005684|Malignant Bladder Neoplasm
C0005684|Malignant Bladder Tumor
C0005684|Malignant Neoplasm of the Bladder
C0005684|Malignant Neoplasm of the Urinary Bladder
C0005684|Malignant Neoplasm, Bladder
C0005684|Malignant Neoplasm, Urinary Bladder
C0005684|Malignant Tumor of the Bladder
C0005684|Malignant Tumor of the Urinary Bladder
C0005684|Malignant Tumor, Urinary Bladder
C0005684|Malignant Urinary Bladder Neoplasm
C0005684|Malignant Urinary Bladder Tumor
C0005684|Urinary Bladder Malignant Neoplasm
C0005684|Urinary Bladder Malignant Tumor
C0005684|Neoplasm malig;bladder
C0005684|malignant neosplasm of the bladder
C0496827|Dome of bladder
C0496827|Malignant neoplasm of dome of bladder
C0496827|Malignant neoplasm of apex of urinary bladder
C0496827|malignant neoplasm of dome of bladder (diagnosis)
C0496827|malignant tumor of dome of bladder
C0496827|Mal neo bladder-dome
C0496827|Malignant neoplasm of dome of urinary bladder
C0496827|BLADDER, DOME
C0496827|Dome of the Bladder
C0496827|Malignant tumor of bladder dome
C0496827|Malignant tumor of vault of bladder
C0496827|Malignant tumour of bladder dome
C0496827|Malignant tumour of vault of bladder
C0496827|Malignant neoplasm of vault of bladder
C0496827|Malignant tumor of vault of bladder (disorder)
C0496827|Superior Surface of Bladder
C0496827|Superior Surface of the Bladder
C0496828|Lateral wall of bladder
C0496828|Malignant neoplasm of lateral wall of bladder
C0496828|Malignant neoplasm of lateral wall of urinary bladder
C0496828|malignant neoplasm of lateral wall of bladder (diagnosis)
C0496828|malignant tumor of lateral wall of bladder
C0496828|Mal neo bladder-lateral
C0496828|Malignant neoplasm of lateral wall of urinary bladder (disorder)
C0496828|Lateral Wall of the Bladder
C0349054|Malignant neoplasm overlapping bladder site
C0349054|Overlapping lesion of bladder
C0349054|Malignant neoplasm of overlapping sites of bladder
C0349054|malignant neoplasm bladder overlapping sites
C0349054|malignant neoplasm of overlapping sites of bladder (diagnosis)
C0349054|Overlapping malignant neoplasm of bladder
C0349054|Overlapping malignant neoplasm of urinary bladder (disorder)
C0349054|Overlapping malignant neoplasm of urinary bladder
C0349054|Malignant neoplasm, overlapping lesion of bladder
C0349054|Malignant neoplasm, overlapping lesion of bladder (disorder)
C0153612|Malignant neoplasm of posterior wall of urinary bladder
C0153612|Malignant neoplasm of posterior wall of bladder
C0153612|Posterior wall of bladder
C0153612|malignant neoplasm of posterior wall of bladder (diagnosis)
C0153612|malignant tumor of posterior wall of bladder
C0153612|Mal neo bladder-post
C0153612|Malignant neoplasm of posterior wall of urinary bladder (disorder)
C0496826|Malignant neoplasm of trigone of bladder
C0496826|Trigone of bladder
C0496826|Malignant neoplasm of trigone of urinary bladder
C0496826|malignant neoplasm of trigone of bladder (diagnosis)
C0496826|malignant tumor of trigone of bladder
C0496826|Mal neo bladder-trigone
C0496826|Malignant tumour of trigone of bladder
C0496826|Malignant tumor of trigone of bladder (disorder)
C0496826|Malignant tumor of trigone of urinary bladder
C0496826|Malignant tumour of trigone of urinary bladder
C0496826|Malignant tumor of trigone of urinary bladder (disorder)
C0153614|Malignant neoplasm of ureteric orifice
C0153614|Ureteric orifice
C0153614|Malignant neoplasm of ureteric orifice of urinary bladder
C0153614|malignant neoplasm of ureteric orifice (diagnosis)
C0153614|malignant tumor of ureteric orifice
C0153614|Mal neo ureteric orifice
C0153614|cancer of ureteral orifice
C0153614|cancer of ureteric orifice
C0153614|Ureteral Opening
C0153614|Uteric Orifice
C0153614|Malignant tumour of ureteric orifice
C0153614|Malignant tumor of ureteric orifice (disorder)
C0153614|Orifice of the Ureter
C0855174|Bladder adenocarcinoma recurrent
C0855174|Recurrent Adenocarcinoma of Bladder
C0855174|Recurrent Adenocarcinoma of Urinary Bladder
C0855174|Recurrent Adenocarcinoma of the Bladder
C0855174|Recurrent Adenocarcinoma of the Urinary Bladder
C0855174|Recurrent Bladder Adenocarcinoma
C0855174|Recurrent Urinary Bladder Adenocarcinoma
C0855174|Relapsed Adenocarcinoma of Bladder
C0855174|Relapsed Adenocarcinoma of Urinary Bladder
C0855174|Relapsed Adenocarcinoma of the Bladder
C0855174|Relapsed Adenocarcinoma of the Urinary Bladder
C0855174|Relapsed Bladder Adenocarcinoma
C0855174|Relapsed Urinary Bladder Adenocarcinoma
C0855174|Bladder Adenocarcinoma, Recurrent
C0855175|Bladder adenocarcinoma stage 0
C0855175|Stage 0 Bladder Adenocarcinoma AJCC v7
C0855175|Stage 0 Bladder Adenocarcinoma AJCC v6
C0855175|Stage 0 Bladder Adenocarcinoma
C0855176|Bladder adenocarcinoma stage I
C0855176|Stage I Bladder Adenocarcinoma AJCC v7
C0855176|Stage I Bladder Adenocarcinoma AJCC v6
C0855176|Stage I Bladder Adenocarcinoma
C0855177|Bladder adenocarcinoma stage II
C0855177|Stage II Bladder Adenocarcinoma AJCC v6
C0855177|Stage II Bladder Adenocarcinoma AJCC v7
C0855177|Stage II Bladder Adenocarcinoma
C0855178|Bladder adenocarcinoma stage III
C0855178|Stage III Bladder Adenocarcinoma AJCC v7
C0855178|Stage III Bladder Adenocarcinoma AJCC v6
C0855178|Stage III Bladder Adenocarcinoma
C0855179|Bladder adenocarcinoma stage IV
C0855179|Stage IV Bladder Adenocarcinoma AJCC v7
C0855179|Stage IV Bladder Adenocarcinoma
C0855180|Bladder adenocarcinoma stage unspecified
C0278827|Ca bladder recurrent
C0278827|Bladder cancer recurrent
C0278827|Recurrent Bladder Cancer
C0278827|Recurrent Bladder Carcinoma
C0278827|Carcinoma urinary bladder recurrent
C0278827|Urinary bladder carcinoma recurrent
C0278827|Carcinoma bladder recurrent
C0278827|Bladder carcinoma recurrent
C0278827|bladder cancer, recurrent
C0278827|cancer of the bladder, recurrent
C0278827|carcinoma of the bladder, recurrent
C0278827|recurrent cancer of the bladder
C0278827|recurrent carcinoma of the bladder
C0278827|Recurrent Cancer of Bladder
C0278827|Recurrent Cancer of Urinary Bladder
C0278827|Recurrent Cancer of the Urinary Bladder
C0278827|Recurrent Urinary Bladder Cancer
C0278827|Relapsed Bladder Cancer
C0278827|Relapsed Cancer of Bladder
C0278827|Relapsed Cancer of Urinary Bladder
C0278827|Relapsed Cancer of the Bladder
C0278827|Relapsed Cancer of the Urinary Bladder
C0278827|Relapsed Urinary Bladder Cancer
C0855181|Ca bladder stage 0, with cancer in situ
C0855181|Bladder cancer stage 0, with cancer in situ
C0855181|Malignant neoplasm of bladder stage 0, with cancer in situ
C0855182|Ca bladder stage 0, without cancer in situ
C0855182|Bladder cancer stage 0, without cancer in situ
C0855182|Malignant neoplasm of bladder stage 0, without cancer in situ
C0855183|Ca bladder stage I, with cancer in situ
C0855183|Bladder cancer stage I, with cancer in situ
C0855183|Malignant neoplasm of bladder stage I, with cancer in situ
C0855185|Ca bladder stage I, without cancer in situ
C0855185|Bladder cancer stage I, without cancer in situ
C0855185|Malignant neoplasm of bladder stage I, without cancer in situ
C0278823|Ca bladder stage II
C0278823|Bladder cancer stage II
C0278823|Stage II Bladder Carcinoma AJCC v7
C0278823|Stage II Bladder Cancer AJCC v7
C0278823|Stage II Bladder Cancer AJCC v6
C0278823|Stage II Bladder Carcinoma AJCC v6
C0278823|stage II bladder cancer
C0278823|Carcinoma urinary bladder stage II
C0278823|Carcinoma bladder stage II
C0278823|Bladder carcinoma stage II
C0278823|Urinary bladder carcinoma stage II
C0278823|bladder cancer, stage B1
C0278823|bladder cancer, stage II
C0278823|cancer of the bladder, stage B1
C0278823|cancer of the bladder, stage II
C0278823|carcinoma of the bladder, stage B1
C0278823|carcinoma of the bladder, stage II
C0278823|stage B1 cancer of the bladder
C0278823|stage B1 carcinoma of the bladder
C0278823|stage II cancer of the bladder
C0278823|stage II carcinoma of the bladder
C0278823|Jewett-Marshall Stage B Bladder Cancer
C0278823|Jewett-Marshall Stage B Bladder Carcinoma
C0278823|Jewett-Marshall Stage B Urinary Bladder Cancer
C0278823|Jewett-Marshall Stage B Urinary Bladder Carcinoma
C0278823|Stage II Bladder Carcinoma
C0278823|Stage II Carcinoma of Bladder
C0278823|Stage II Carcinoma of Urinary Bladder
C0278823|Stage II Carcinoma of the Urinary Bladder
C0278823|Stage II Urinary Bladder Carcinoma
C0278823|Cancer of Bladder Stage II
C0278823|Cancer of the Bladder Stage II
C0278824|Ca bladder stage III
C0278824|Bladder cancer stage III
C0278824|Stage III Bladder Cancer AJCC v6
C0278824|Stage III Bladder Carcinoma AJCC v7
C0278824|Stage III Bladder Cancer AJCC v7
C0278824|Stage III Bladder Carcinoma AJCC v6
C0278824|stage III bladder cancer
C0278824|Carcinoma bladder stage III
C0278824|Carcinoma urinary bladder stage III
C0278824|Bladder carcinoma stage III
C0278824|Urinary bladder carcinoma stage III
C0278824|bladder cancer, stage III
C0278824|cancer of the bladder, stage III
C0278824|carcinoma of the bladder, stage III
C0278824|stage III cancer of the bladder
C0278824|stage III carcinoma of the bladder
C0278824|Jewett-Marshall Stage C Bladder Cancer
C0278824|Jewett-Marshall Stage C Urinary Bladder Cancer
C0278824|Jewett-Marshall Stage C Urinary Bladder Carcinoma
C0278824|Stage III Bladder Carcinoma
C0278824|Stage III Carcinoma of Bladder
C0278824|Stage III Carcinoma of Urinary Bladder
C0278824|Stage III Carcinoma of the Urinary Bladder
C0278824|Stage III Urinary Bladder Carcinoma
C0278824|Cancer of Bladder Stage III
C0278824|Cancer of the Bladder Stage III
C0278828|Ca bladder stage IV
C0278828|Bladder cancer stage IV
C0278828|Cancer of Bladder Stage IV AJCC v6
C0278828|Stage IV Carcinoma of the Bladder AJCC v6
C0278828|Cancer of the Bladder Stage IV AJCC v6
C0278828|Stage IV Carcinoma of Urinary Bladder AJCC v6
C0278828|Stage IV Carcinoma of the Urinary Bladder AJCC v6
C0278828|Stage IV Urinary Bladder Carcinoma AJCC v6
C0278828|Stage IV Carcinoma of Bladder AJCC v6
C0278828|Stage IV Bladder Cancer AJCC v6
C0278828|Stage IV Bladder Carcinoma AJCC v6
C0278828|Metastatic carcinoma of the bladder
C0278828|stage IV bladder cancer
C0278828|Urinary bladder carcinoma stage IV
C0278828|Carcinoma bladder stage IV
C0278828|Carcinoma urinary bladder stage IV
C0278828|Bladder carcinoma stage IV
C0278828|bladder cancer, metastatic
C0278828|bladder cancer, stage IV
C0278828|cancer of the bladder, metastatic
C0278828|cancer of the bladder, stage IV
C0278828|carcinoma of the bladder, metastatic
C0278828|carcinoma of the bladder, stage IV
C0278828|metastatic bladder cancer
C0278828|metastatic cancer of the bladder
C0278828|stage IV cancer of the bladder
C0278828|stage IV carcinoma of the bladder
C0278828|Jewett-Marshall Stage D Bladder Cancer
C0278828|Jewett-Marshall Stage D Bladder Carcinoma
C0278828|Jewett-Marshall Stage D Urinary Bladder Cancer
C0278828|Jewett-Marshall Stage D Urinary Bladder Carcinoma
C0855186|Bladder squamous cell carcinoma recurrent
C0855186|Squamous cell carcinoma of the bladder recurrent
C0855186|Squamous cell bladder carcinoma recurrent
C0855186|Recurrent Bladder Epidermoid Carcinoma
C0855186|Recurrent Bladder Squamous Cell Carcinoma
C0855186|Recurrent Epidermoid Carcinoma of Bladder
C0855186|Recurrent Epidermoid Carcinoma of Urinary Bladder
C0855186|Recurrent Epidermoid Carcinoma of the Bladder
C0855186|Recurrent Epidermoid Carcinoma of the Urinary Bladder
C0855186|Recurrent Squamous Cell Carcinoma of Bladder
C0855186|Recurrent Squamous Cell Carcinoma of Urinary Bladder
C0855186|Recurrent Squamous Cell Carcinoma of the Bladder
C0855186|Recurrent Squamous Cell Carcinoma of the Urinary Bladder
C0855186|Recurrent Urinary Bladder Epidermoid Carcinoma
C0855186|Recurrent Urinary Bladder Squamous Cell Carcinoma
C0855186|Relapsed Bladder Epidermoid Carcinoma
C0855186|Relapsed Bladder Squamous Cell Carcinoma
C0855186|Relapsed Epidermoid Carcinoma of Bladder
C0855186|Relapsed Epidermoid Carcinoma of Urinary Bladder
C0855186|Relapsed Epidermoid Carcinoma of the Bladder
C0855186|Relapsed Epidermoid Carcinoma of the Urinary Bladder
C0855186|Relapsed Squamous Cell Carcinoma of Bladder
C0855186|Relapsed Squamous Cell Carcinoma of Urinary Bladder
C0855186|Relapsed Squamous Cell Carcinoma of the Bladder
C0855186|Relapsed Squamous Cell Carcinoma of the Urinary Bladder
C0855186|Relapsed Urinary Bladder Epidermoid Carcinoma
C0855186|Relapsed Urinary Bladder Squamous Cell Carcinoma
C0855186|Squamous Cell Carcinoma of Bladder, Recurrent
C0855186|Squamous Cell Carcinoma of the Bladder, Recurrent
C0855187|Bladder squamous cell carcinoma stage 0
C0855187|Stage 0 Bladder Squamous Cell Carcinoma AJCC v6
C0855187|Stage 0 Bladder Squamous Cell Carcinoma AJCC v7
C0855187|Squamous cell carcinoma of the bladder stage 0
C0855187|Squamous cell bladder carcinoma stage 0
C0855187|Stage 0 Bladder Squamous Cell Carcinoma
C0855187|Stage 0 Squamous Cell Carcinoma of Bladder
C0855187|Stage 0 Squamous Cell Carcinoma of the Bladder
C0855188|Bladder squamous cell carcinoma stage I
C0855188|Stage I Squamous Cell Carcinoma of the Bladder AJCC v7
C0855188|Stage I Squamous Cell Carcinoma of the Bladder AJCC v6
C0855188|Squamous cell carcinoma of the bladder stage I
C0855188|Squamous cell bladder carcinoma stage I
C0855188|Stage I Squamous Cell Carcinoma of Bladder
C0855188|Stage I Squamous Cell Carcinoma of the Bladder
C0855189|Bladder squamous cell carcinoma stage II
C0855189|Stage II Bladder Squamous Cell Carcinoma AJCC v6
C0855189|Stage II Bladder Squamous Cell Carcinoma AJCC v7
C0855189|Squamous cell bladder carcinoma stage II
C0855189|Squamous cell carcinoma of the bladder stage II
C0855189|Stage II Bladder Squamous Cell Carcinoma
C0855190|Bladder squamous cell carcinoma stage III
C0855190|Stage III Bladder Squamous Cell Carcinoma AJCC v6
C0855190|Stage III Bladder Squamous Cell Carcinoma AJCC v7
C0855190|Squamous cell bladder carcinoma stage III
C0855190|Squamous cell carcinoma of the bladder stage III
C0855190|Stage III Bladder Squamous Cell Carcinoma
C0855191|Bladder squamous cell carcinoma stage IV
C0855191|Stage IV Bladder Squamous Cell Carcinoma AJCC v7
C0855191|Squamous cell bladder carcinoma stage IV
C0855191|Squamous cell carcinoma of the bladder stage IV
C0855191|Stage IV Bladder Squamous Cell Carcinoma
C0855192|Bladder squamous cell carcinoma stage unspecified
C0855192|Squamous cell carcinoma of the bladder stage unspecified
C0279680|Bladder transitional cell carcinoma
C0279680|Transitional cell carcinoma of the bladder
C0279680|transitional cell carcinoma of bladder
C0279680|transitional cell carcinoma of bladder (diagnosis)
C0279680|Transitional cell carcinoma of bladder (disorder)
C0279680|Bladder Urothelial Carcinoma
C0279680|Transitional cell bladder carcinoma
C0279680|Urothelial carcinoma bladder
C0279680|TCC - Transitional cell carcinoma of bladder
C0279680|bladder cancer, transitional cell carcinoma
C0279680|carcinoma, transitional cell, bladder
C0279680|Transitional Cell Carcinoma of the Urinary Bladder
C0279680|Urinary Bladder Transitional Cell Carcinoma
C0279680|Urinary Bladder Urothelial Carcinoma
C0279680|Urothelial Carcinoma of the Urinary Bladder
C1336089|Non-Invasive Bladder Urothelial Carcinoma
C1336089|Bladder transitional cell carcinoma stage 0
C1336089|Stage 0 Bladder Urothelial Carcinoma AJCC v7
C1336089|Stage 0 Bladder Urothelial Carcinoma AJCC v6
C1336089|Stage 0 Transitional Cell Carcinoma of Bladder
C1336089|Stage 0 Transitional Cell Carcinoma of Urinary Bladder
C1336089|Stage 0 Transitional Cell Carcinoma of the Bladder
C1336089|Stage 0 Transitional Cell Carcinoma of the Urinary Bladder
C1336089|Stage 0 Urinary Bladder Transitional Cell Carcinoma
C1336089|Stage 0 Bladder Urothelial Carcinoma
C1739113|Bladder transitional cell carcinoma recurrent
C1336450|Bladder transitional cell carcinoma stage I
C1336450|Stage I Bladder Urothelial Carcinoma AJCC v6
C1336450|Stage I Bladder Urothelial Carcinoma AJCC v7
C1336450|Stage I Transitional Cell Carcinoma of Bladder
C1336450|Stage I Transitional Cell Carcinoma of Urinary Bladder
C1336450|Stage I Transitional Cell Carcinoma of the Bladder
C1336450|Stage I Transitional Cell Carcinoma of the Urinary Bladder
C1336450|Stage I Urinary Bladder Transitional Cell Carcinoma
C1336450|Stage I Bladder Urothelial Carcinoma
C0862432|Bladder transitional cell carcinoma stage IV
C0862432|Stage IV Bladder Urothelial Carcinoma AJCC v7
C0862432|Transitional cell carcinoma of the bladder stage IV
C0862432|Urothelial carcinoma bladder stage IV
C0862432|Stage IV Transitional Cell Carcinoma of Bladder
C0862432|Stage IV Transitional Cell Carcinoma of Urinary Bladder
C0862432|Stage IV Transitional Cell Carcinoma of the Bladder
C0862432|Stage IV Transitional Cell Carcinoma of the Urinary Bladder
C0862432|Stage IV Urinary Bladder Transitional Cell Carcinoma
C0862432|Stage IV Bladder Urothelial Carcinoma
C0862402|Bladder transitional cell carcinoma stage II
C0862402|Stage II Bladder Urothelial Carcinoma AJCC v6
C0862402|Stage II Bladder Urothelial Carcinoma AJCC v7
C0862402|Urothelial carcinoma bladder stage II
C0862402|Transitional cell carcinoma of the bladder stage II
C0862402|Stage II Transitional Cell Carcinoma of Bladder
C0862402|Stage II Transitional Cell Carcinoma of Urinary Bladder
C0862402|Stage II Transitional Cell Carcinoma of the Bladder
C0862402|Stage II Transitional Cell Carcinoma of the Urinary Bladder
C0862402|Stage II Urinary Bladder Transitional Cell Carcinoma
C0862402|Stage II Bladder Urothelial Carcinoma
C0862417|Bladder transitional cell carcinoma stage III
C0862417|Stage III Bladder Urothelial Carcinoma AJCC v7
C0862417|Stage III Bladder Urothelial Carcinoma AJCC v6
C0862417|Transitional cell carcinoma of the bladder stage III
C0862417|Urothelial carcinoma bladder stage III
C0862417|Stage III Transitional Cell Carcinoma of Bladder
C0862417|Stage III Transitional Cell Carcinoma of Urinary Bladder
C0862417|Stage III Transitional Cell Carcinoma of the Bladder
C0862417|Stage III Transitional Cell Carcinoma of the Urinary Bladder
C0862417|Stage III Urinary Bladder Transitional Cell Carcinoma
C0862417|Stage III Bladder Urothelial Carcinoma
C1297936|malignant neoplasm bladder by direct extension from endometrium
C1297936|malignant neoplasm involving bladder by direct extension from endometrium (diagnosis)
C1297936|malignant neoplasm involving bladder by direct extension from endometrium
C1297936|Malignant tumor involving bladder by direct extension from endometrium (disorder)
C1297936|Malignant tumor involving bladder by direct extension from endometrium
C1297936|Malignant tumour involving bladder by direct extension from endometrium
C1297937|malignant neoplasm involving bladder by direct extension from fallopian tube
C1297937|malignant neoplasm bladder by direct extension from fallopian tube
C1297937|malignant neoplasm involving bladder by direct extension from fallopian tube (diagnosis)
C1297937|Malignant tumor involving bladder by direct extension from fallopian tube (disorder)
C1297937|Malignant tumor involving bladder by direct extension from fallopian tube
C1297937|Malignant tumour involving bladder by direct extension from fallopian tube
C1297938|malignant neoplasm involving bladder by direct extension from ovary (diagnosis)
C1297938|malignant neoplasm involving bladder by direct extension from ovary
C1297938|malignant neoplasm bladder by direct extension from ovary
C1297938|Malignant tumor involving bladder by direct extension from ovary (disorder)
C1297938|Malignant tumor involving bladder by direct extension from ovary
C1297938|Malignant tumour involving bladder by direct extension from ovary
C1297939|malignant neoplasm involving bladder by direct extension from prostate
C1297939|malignant neoplasm bladder by direct extension from prostate
C1297939|malignant neoplasm involving bladder by direct extension from prostate (diagnosis)
C1297939|Malignant tumor involving bladder by direct extension from prostate (disorder)
C1297939|Malignant tumor involving bladder by direct extension from prostate
C1297939|Malignant tumour involving bladder by direct extension from prostate
C1297940|malignant neoplasm involving bladder by direct extension from uterine cervix
C1297940|malignant neoplasm bladder by direct extension from uterine cervix
C1297940|malignant neoplasm involving bladder by direct extension from uterine cervix (diagnosis)
C1297940|Malignant tumor involving bladder by direct extension from uterine cervix (disorder)
C1297940|Malignant tumor involving bladder by direct extension from uterine cervix
C1297940|Malignant tumour involving bladder by direct extension from uterine cervix
C1297941|malignant neoplasm involving bladder by direct extension from uterus
C1297941|malignant neoplasm involving bladder by direct extension from uterus (diagnosis)
C1297941|malignant neoplasm bladder by direct extension from uterus
C1297941|Malignant tumor involving bladder by direct extension from uterus (disorder)
C1297941|Malignant tumor involving bladder by direct extension from uterus
C1297941|Malignant tumour involving bladder by direct extension from uterus
C1297942|malignant neoplasm involving bladder by direct extension from vagina
C1297942|malignant neoplasm involving bladder by direct extension from vagina (diagnosis)
C1297942|malignant neoplasm bladder by direct extension from vagina
C1297942|Malignant tumor involving bladder by direct extension from vagina (disorder)
C1297942|Malignant tumor involving bladder by direct extension from vagina
C1297942|Malignant tumour involving bladder by direct extension from vagina
C2033201|papillary carcinoma of bladder (diagnosis)
C2033201|papillary carcinoma of bladder
C2212520|Mullerian mixed tumor of bladder
C2212520|Mullerian mixed tumor of bladder (diagnosis)
C2212529|malignant mesodermal mixed tumor of bladder
C2212529|malignant mesodermal mixed tumor of bladder (diagnosis)
C2212590|malignant small cell neoplasm of bladder (diagnosis)
C2212590|malignant small cell neoplasm of bladder
C2011424|giant cell type neoplasm of bladder
C2011424|giant cell type neoplasm of bladder (diagnosis)
C2018634|spindle cell type neoplasm of bladder (diagnosis)
C2018634|spindle cell type neoplasm of bladder
C2075593|clear cell type neoplasm of bladder (diagnosis)
C2075593|clear cell type neoplasm of bladder
C1334563|malignant paraganglioma of bladder (diagnosis)
C1334563|malignant paraganglioma of bladder
C1334563|Malignant Bladder Paraganglioma
C1334563|Malignant Paraganglioma of Urinary Bladder
C1334563|Malignant Paraganglioma of the Bladder
C1334563|Malignant Paraganglioma of the Urinary Bladder
C1334563|Malignant Urinary Bladder Paraganglioma
C2212603|myosarcoma of bladder
C2212603|myosarcoma of bladder (diagnosis)
C2212605|fibrous histiocytoma of bladder (diagnosis)
C2212605|fibrous histiocytoma of bladder
C0279682|adenocarcinoma of bladder
C0279682|adenocarcinoma of bladder (diagnosis)
C0279682|bladder adenocarcinoma
C0279682|Adenocarcinoma of bladder (disorder)
C0279682|adenocarcinoma of the bladder
C0279682|adenocarcinoma, bladder
C0279682|bladder cancer, adenocarcinoma
C0279682|Adenocarcinoma of Urinary Bladder
C0279682|Adenocarcinoma of the Urinary Bladder
C0279682|Urinary Bladder Adenocarcinoma
C0279682|Bladder Adenocarcinoma NOS
C0279682|Bladder Adenocarcinoma, NOS
C0279682|Bladder Adenocarcinoma, Not Otherwise Specified
C2007062|carcinosarcoma of bladder (diagnosis)
C2007062|carcinosarcoma of bladder
C0349666|sarcoma of bladder
C0349666|sarcoma of bladder (diagnosis)
C0349666|Urinary bladder sarcoma
C0349666|Sarcoma of bladder (disorder)
C0349666|Sarcoma of Urinary Bladder
C0349666|Sarcoma of the Bladder
C0349666|Sarcoma of the Urinary Bladder
C0349666|Bladder Sarcoma
C2212616|fibrosarcoma of bladder (diagnosis)
C2212616|fibrosarcoma of bladder
C2212627|malignant mesenchymoma of bladder (diagnosis)
C2212627|malignant mesenchymoma of bladder
C2212628|malignant lymphoma of bladder (diagnosis)
C2212628|malignant lymphoma of bladder
C2212659|malignant plasmacytoma of bladder
C2212659|malignant plasmacytoma of bladder (diagnosis)
C2212661|malignant mastocytosis of bladder
C2212661|malignant mastocytosis of bladder (diagnosis)
C2216667|staging of bladder cancer
C2216667|staging of malignant neoplasm of bladder (diagnosis)
C2216667|staging of malignant neoplasm of bladder
C2216667|malignant neoplasm of bladder staging
C0699885|CARCINOMA OF BLADDER
C0699885|Bladder carcinoma
C0699885|carcinoma of bladder (diagnosis)
C0699885|Carcinoma;bladder
C0699885|Carcinoma bladder
C0699885|bladder cancer
C0699885|Bladder carcinoma NOS
C0699885|Carcinoma urinary bladder
C0699885|Urinary bladder carcinoma
C0699885|Carcinoma of bladder (disorder)
C0699885|carcinoma of the bladder
C0699885|Cancer of Bladder
C0699885|Cancer of the Bladder
C0699885|Urinary Bladder Cancer
C0699885|Cancer of the Urinary Bladder
C0699885|Carcinoma of Urinary Bladder
C0699885|Carcinoma of the Urinary Bladder
C0699885|Cancer of Urinary Bladder
C2212587|noninvasive papillary transitional cell carcinoma in situ of bladder
C2212587|noninvasive papillary transitional cell carcinoma in situ of bladder (diagnosis)
C2212587|bladder carcinoma in situ papillary transitional cell noninvasive
C2212591|signet ring cell carcinoma of bladder (diagnosis)
C2212591|signet ring cell carcinoma of bladder
C2212592|malignant epithelioma of bladder (diagnosis)
C2212592|malignant epithelioma of bladder
C2111591|large cell carcinoma of bladder
C2111591|large cell carcinoma of bladder (diagnosis)
C2111710|large cell neuroendocrine carcinoma of bladder (diagnosis)
C2111710|large cell neuroendocrine carcinoma of bladder
C2111592|large cell carcinoma of bladder with rhabdoid phenotype
C2111592|bladder malignant carcinoma large cell with rhabdoid phenotype
C2111592|large cell carcinoma of bladder with rhabdoid phenotype (diagnosis)
C2012070|glassy cell carcinoma of bladder
C2012070|glassy cell carcinoma of bladder (diagnosis)
C2188054|undifferentiated carcinoma of bladder (diagnosis)
C2188054|undifferentiated carcinoma of bladder
C2212593|anaplastic carcinoma of bladder (diagnosis)
C2212593|anaplastic carcinoma of bladder
C2082422|pleomorphic carcinoma of bladder (diagnosis)
C2082422|pleomorphic carcinoma of bladder
C2011242|giant cell carcinoma of bladder (diagnosis)
C2011242|giant cell carcinoma of bladder
C2018384|spindle cell carcinoma of bladder (diagnosis)
C2018384|spindle cell carcinoma of bladder
C2011207|giant cell and spindle cell carcinoma of bladder (diagnosis)
C2011207|giant cell and spindle cell carcinoma of bladder
C2142912|pseudosarcomatous carcinoma of bladder
C2142912|pseudosarcomatous carcinoma of bladder (diagnosis)
C2111794|polygonal cell carcinoma of bladder
C2111794|polygonal cell carcinoma of bladder (diagnosis)
C2007057|carcinoma of bladder with osteoclast-like giant cells (diagnosis)
C2007057|carcinoma of bladder with osteoclast-like giant cells
C2007057|bladder carcinoma with osteoclast-like giant cells
C2212594|small cell carcinoma of bladder (diagnosis)
C2212594|small cell carcinoma of bladder
C2009873|fusiform type small cell carcinoma of bladder (diagnosis)
C2009873|fusiform type small cell carcinoma of bladder
C2212595|medullary carcinoma of bladder (diagnosis)
C2212595|medullary carcinoma of bladder
C2033276|papillary squamous cell carcinoma of bladder
C2033276|papillary squamous cell carcinoma of bladder (diagnosis)
C1511208|verrucous carcinoma of bladder (diagnosis)
C1511208|verrucous carcinoma of bladder
C1511208|Bladder Verrucous Carcinoma
C1511208|Bladder Verrucous Squamous Cell Carcinoma
C2018592|spindle cell transitional cell carcinoma of bladder
C2018592|spindle cell transitional cell carcinoma of bladder (diagnosis)
C1735888|papillary transitional cell carcinoma of bladder (diagnosis)
C1735888|papillary transitional cell carcinoma of bladder
C2212600|micropapillary transitional cell carcinoma of bladder
C2212600|micropapillary transitional cell carcinoma of bladder (diagnosis)
C2212601|Schneiderian carcinoma of bladder
C2212601|Schneiderian carcinoma of bladder (diagnosis)
C2212602|basaloid carcinoma of bladder
C2212602|basaloid carcinoma of bladder (diagnosis)
C2075828|cloacogenic carcinoma of bladder (diagnosis)
C2075828|cloacogenic carcinoma of bladder
C2007045|carcinoma simplex of bladder (diagnosis)
C2007045|carcinoma simplex of bladder
C2012537|granular cell carcinoma of bladder (diagnosis)
C2012537|granular cell carcinoma of bladder
C2017446|solid carcinoma of bladder (diagnosis)
C2017446|solid carcinoma of bladder
C3203710|Bladder transitional cell carcinoma metastatic
C2033152|papillary carcinoma in situ of bladder (diagnosis)
C2033152|papillary carcinoma in situ of bladder
C2212585|bladder carcinoma in situ papillary squamous cell noninvasive
C2212585|noninvasive papillary squamous cell carcinoma in situ of bladder
C2212585|noninvasive papillary squamous cell carcinoma in situ of bladder (diagnosis)
C2019360|squamous cell carcinoma in situ of bladder (diagnosis)
C2019360|squamous cell carcinoma in situ of bladder
C2212586|bladder CIS squamous cell with questionable stromal invasion
C2212586|bladder carcinoma in situ squamous cell with questionable stromal invasion
C2212586|squamous cell carcinoma in situ of bladder with questionable stromal invasion (diagnosis)
C2212586|squamous cell carcinoma in situ of bladder with questionable stromal invasion
C2145423|transitional cell carcinoma in situ of bladder
C2145423|transitional cell carcinoma in situ of bladder (diagnosis)
C2212589|bladder adenocarcinoma in situ in villous adenoma
C2212589|adenocarcinoma in situ in villous adenoma of bladder
C2212589|adenocarcinoma in situ in villous adenoma of bladder (diagnosis)
C2199211|ductal carcinoma in situ of bladder
C2199211|ductal carcinoma in situ of bladder (diagnosis)
C0346893|Malignant neoplasm of other site of urinary bladder (disorder)
C0346893|Malignant neoplasm of other site of urinary bladder
C1314699|bladder malignant neoplasm primary
C1314699|Primary malignant neoplasm of bladder (diagnosis)
C1314699|Primary malignant neoplasm of bladder
C1314699|Primary malignant neoplasm of bladder (disorder)
C1282481|malignant neoplasm bladder, local recurrence
C1282481|local recurrence of malignant neoplasm of bladder
C1282481|local recurrence of malignant neoplasm of bladder (diagnosis)
C1282481|Local recurrence of malignant tumor of urinary bladder (disorder)
C1282481|Local recurrence of malignant tumor of urinary bladder
C1282481|Local recurrence of malignant tumour of urinary bladder
C0347011|Metastatic Neoplasm to the Bladder
C0347011|metastasis to bladder (diagnosis)
C0347011|metastasis to bladder
C0347011|metastasis to the bladder
C0347011|Secondary malignant neoplasm of bladder
C0347011|Metastases to bladder
C0347011|secondary malignant neoplasm urinary bladder
C0347011|secondary malignant neoplasm of bladder (diagnosis)
C0347011|Metastatic Malignant Neoplasm to the Bladder
C0347011|Metastatic Malignant Neoplasm in the Bladder
C0347011|Cancer metastatic to urinary bladder
C0347011|Metastatic tumor to bladder
C0347011|Metastatic tumour to bladder
C0347011|Metastatic malignant neoplasm to bladder
C0347011|Secondary malignant neoplasm of bladder (disorder)
C0347011|Metastatic malignant neoplasm to bladder, NOS
C0347011|Secondary malignant neoplasm of bladder, NOS
C0347011|Metastatic Neoplasm to the Urinary Bladder
C0347011|Metastatic Tumor to the Bladder
C0347011|Metastatic Tumor to the Urinary Bladder
C3694329|malignant neoplasm of apex of bladder (diagnosis)
C3694329|malignant neoplasm of apex of bladder
C3694329|malignant neoplasm bladder apex
C1282497|metastasis from malignant neoplasm of bladder
C1282497|metastasis from malignant neoplasm of bladder (diagnosis)
C1282497|Metastasis from malignant tumor of bladder (disorder)
C1282497|Metastasis from malignant tumor of bladder
C1282497|Metastasis from malignant tumour of bladder
C3839273|Malignant neoplasm of augmented bladder (disorder)
C3839273|Malignant neoplasm of augmented bladder
C3839273|Malignant tumor of augmented bladder
C3839273|Malignant tumour of augmented bladder
C4031688|biopsy of bladder showed hodgkin's lymphoma nodular lymphocytic predominance
C4031688|biopsy of bladder showed hodgkin's lymphoma nodular lymphocytic predominance (procedure)
C4031667|biopsy of bladder showed lymphoma mantle cell
C4031667|biopsy of bladder showed lymphoma mantle cell (procedure)
C4031656|biopsy of bladder showed mastocytosis
C4031656|biopsy of bladder showed mastocytosis (procedure)
C4031722|biopsy of bladder showed carcinoma squamous cell keratinizing (procedure)
C4031722|biopsy of bladder showed carcinoma squamous cell keratinizing
C4031707|biopsy of bladder showed carcinosarcoma embryonal type
C4031707|biopsy of bladder showed carcinosarcoma embryonal type (procedure)
C4031671|biopsy of bladder showed lymphoma histiocytosis
C4031671|biopsy of bladder showed lymphoma histiocytosis (procedure)
C4031670|biopsy of bladder showed lymphoma large b-cell diffuse
C4031670|biopsy of bladder showed lymphoma large b-cell diffuse (procedure)
C4031648|biopsy of bladder showed myosarcoma leiomyosarcoma epithelioid
C4031648|biopsy of bladder showed myosarcoma leiomyosarcoma epithelioid (procedure)
C4031736|biopsy of bladder showed carcinoma papillary
C4031736|biopsy of bladder showed carcinoma papillary (procedure)
C4031735|biopsy of bladder showed carcinoma papillary squamous cell
C4031735|biopsy of bladder showed carcinoma papillary squamous cell (procedure)
C4031714|biopsy of bladder showed carcinoma transitional cell micropapillary (procedure)
C4031714|biopsy of bladder showed carcinoma transitional cell micropapillary
C4031661|biopsy of bladder showed lymphoma precursor cell lymphoblastic
C4031661|biopsy of bladder showed lymphoma precursor cell lymphoblastic (procedure)
C4031655|biopsy of bladder showed mesenchymoma (procedure)
C4031655|biopsy of bladder showed mesenchymoma
C4031641|biopsy of bladder showed myosarcoma rhabdomyosarcoma spindle cell (procedure)
C4031641|biopsy of bladder showed myosarcoma rhabdomyosarcoma spindle cell
C4031628|biopsy of bladder showed sarcoma follicular dendritic cell (procedure)
C4031628|biopsy of bladder showed sarcoma follicular dendritic cell
C4031749|biopsy of bladder showed carcinoma basaloid (procedure)
C4031749|biopsy of bladder showed carcinoma basaloid
C4031717|biopsy of bladder showed carcinoma squamous cell with horn formation
C4031717|biopsy of bladder showed carcinoma squamous cell with horn formation (procedure)
C4031706|biopsy of bladder showed carcinosarcoma myoepithelioma
C4031706|biopsy of bladder showed carcinosarcoma myoepithelioma (procedure)
C4031703|biopsy of bladder showed clear cell type
C4031703|biopsy of bladder showed clear cell type (procedure)
C4031702|biopsy of bladder showed fibrosarcoma
C4031702|biopsy of bladder showed fibrosarcoma (procedure)
C4031691|biopsy of bladder showed hodgkin's lymphoma lymphocytic depletion
C4031691|biopsy of bladder showed hodgkin's lymphoma lymphocytic depletion (procedure)
C4031672|biopsy of bladder showed lymphoma follicular grade 3 (procedure)
C4031672|biopsy of bladder showed lymphoma follicular grade 3
C4031652|biopsy of bladder showed mullerian mixed tumor
C4031652|biopsy of bladder showed mullerian mixed tumor (procedure)
C4031644|biopsy of bladder showed myosarcoma rhabdomyosarcoma embryonal
C4031644|biopsy of bladder showed myosarcoma rhabdomyosarcoma embryonal (procedure)
C4031640|biopsy of bladder showed myosarcoma rhabdomyosarcoma with ganglionic differentiation
C4031640|biopsy of bladder showed myosarcoma rhabdomyosarcoma with ganglionic differentiation (procedure)
C4031746|biopsy of bladder showed carcinoma giant cell (procedure)
C4031746|biopsy of bladder showed carcinoma giant cell
C4031745|biopsy of bladder showed carcinoma giant sell and spindle cell
C4031745|biopsy of bladder showed carcinoma giant sell and spindle cell (procedure)
C4031726|biopsy of bladder showed carcinoma solid (procedure)
C4031726|biopsy of bladder showed carcinoma solid
C4031695|biopsy of bladder showed hepatoid adenocarcinoma (procedure)
C4031695|biopsy of bladder showed adenocarcinoma hepatoid
C4031695|biopsy of bladder showed hepatoid adenocarcinoma
C4031687|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis
C4031687|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis (procedure)
C4031677|biopsy of bladder showed lymphoma burkitt's
C4031677|biopsy of bladder showed lymphoma burkitt's (procedure)
C4031659|biopsy of bladder showed lymphoma precursor cell lymphoblastic t-cell
C4031659|biopsy of bladder showed lymphoma precursor cell lymphoblastic t-cell (procedure)
C4031647|biopsy of bladder showed myosarcoma leiomyosarcoma myxoid (procedure)
C4031647|biopsy of bladder showed myosarcoma leiomyosarcoma myxoid
C4031645|biopsy of bladder showed myosarcoma rhabdomyosarcoma alveolar (procedure)
C4031645|biopsy of bladder showed myosarcoma rhabdomyosarcoma alveolar
C4031627|biopsy of bladder showed sarcoma giant cell (procedure)
C4031627|biopsy of bladder showed sarcoma giant cell
C4031623|biopsy of bladder showed sarcoma mast cell (procedure)
C4031623|biopsy of bladder showed sarcoma mast cell
C4031728|biopsy of bladder showed carcinoma small cell (procedure)
C4031728|biopsy of bladder showed carcinoma small cell
C4031690|biopsy of bladder showed hodgkin's lymphoma lymphocytic depletion reticular
C4031690|biopsy of bladder showed hodgkin's lymphoma lymphocytic depletion reticular (procedure)
C4031686|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis cellular phase
C4031686|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis cellular phase (procedure)
C4031683|biopsy of bladder showed hodgkin's lymphoma sarcoma
C4031683|biopsy of bladder showed hodgkin's lymphoma sarcoma (procedure)
C4031674|biopsy of bladder showed lymphoma follicular grade 1 (procedure)
C4031674|biopsy of bladder showed lymphoma follicular grade 1
C4031669|biopsy of bladder showed lymphoma large b-cell diffuse immunoblastic (procedure)
C4031669|biopsy of bladder showed lymphoma large b-cell diffuse immunoblastic
C4031651|biopsy of bladder showed myosarcoma
C4031651|biopsy of bladder showed myosarcoma (procedure)
C4031634|biopsy of bladder showed plasmacytoma
C4031634|biopsy of bladder showed plasmacytoma (procedure)
C4031632|biopsy of bladder showed sarcoma (procedure)
C4031632|biopsy of bladder showed sarcoma
C4031625|biopsy of bladder showed sarcoma interdigitating dendritic cell (procedure)
C4031625|biopsy of bladder showed sarcoma interdigitating dendritic cell
C4031620|biopsy of bladder showed sarcoma undifferentiated
C4031620|biopsy of bladder showed sarcoma undifferentiated (procedure)
C4031730|biopsy of bladder showed carcinoma signet ring cell
C4031730|biopsy of bladder showed carcinoma signet ring cell (procedure)
C4031729|biopsy of bladder showed carcinoma simplex
C4031729|biopsy of bladder showed carcinoma simplex (procedure)
C4031701|biopsy of bladder showed fibrosarcoma fascial
C4031701|biopsy of bladder showed fibrosarcoma fascial (procedure)
C4031697|biopsy of bladder showed fibrous histiocytoma (procedure)
C4031697|biopsy of bladder showed fibrous histiocytoma
C4031668|biopsy of bladder showed lymphoma lymphoplasmacytic (procedure)
C4031668|biopsy of bladder showed lymphoma lymphoplasmacytic
C4031630|biopsy of bladder showed sarcoma embryonal (procedure)
C4031630|biopsy of bladder showed sarcoma embryonal
C4031626|biopsy of bladder showed sarcoma histiocytic
C4031626|biopsy of bladder showed sarcoma histiocytic (procedure)
C4031621|biopsy of bladder showed sarcoma spindle cell (procedure)
C4031621|biopsy of bladder showed sarcoma spindle cell
C4031750|biopsy of bladder showed carcinoma anaplastic
C4031750|biopsy of bladder showed carcinoma anaplastic (procedure)
C4031743|biopsy of bladder showed carcinoma granular cell (procedure)
C4031743|biopsy of bladder showed carcinoma granular cell
C4031739|biopsy of bladder showed carcinoma large cell neuroendocrine
C4031739|biopsy of bladder showed carcinoma large cell neuroendocrine (procedure)
C4031737|biopsy of bladder showed carcinoma medullary
C4031737|biopsy of bladder showed carcinoma medullary (procedure)
C4031732|biopsy of bladder showed carcinoma pseudosarcomatous
C4031732|biopsy of bladder showed carcinoma pseudosarcomatous (procedure)
C4031719|biopsy of bladder showed carcinoma squamous cell small cell, nonkeratinizing (procedure)
C4031719|biopsy of bladder showed carcinoma squamous cell small cell, nonkeratinizing
C4031698|biopsy of bladder showed fibrosarcoma solitary fibrous tumor
C4031698|biopsy of bladder showed fibrosarcoma solitary fibrous tumor (procedure)
C4031684|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis grade 2 (procedure)
C4031684|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis grade 2
C4031675|biopsy of bladder showed lymphoma follicular
C4031675|biopsy of bladder showed lymphoma follicular (procedure)
C4031633|biopsy of bladder showed plasmacytoma extramedullary
C4031633|biopsy of bladder showed plasmacytoma extramedullary (procedure)
C4031624|biopsy of bladder showed sarcoma langerhans cell (procedure)
C4031624|biopsy of bladder showed sarcoma langerhans cell
C4031725|biopsy of bladder showed carcinoma spindle cell (procedure)
C4031725|biopsy of bladder showed carcinoma spindle cell
C4031700|biopsy of bladder showed fibrosarcoma fibromyxosarcoma (procedure)
C4031700|biopsy of bladder showed fibrosarcoma fibromyxosarcoma
C4031681|biopsy of bladder showed lymphoma (procedure)
C4031681|biopsy of bladder showed lymphoma
C4031666|biopsy of bladder showed lymphoma marginal zone b-cell (procedure)
C4031666|biopsy of bladder showed lymphoma marginal zone b-cell
C4031664|biopsy of bladder showed lymphoma mature t-cell angioimmunoblastic (procedure)
C4031664|biopsy of bladder showed lymphoma mature t-cell angioimmunoblastic
C4031657|biopsy of bladder showed malignant neoplasm
C4031657|biopsy of bladder showed malignant neoplasm (procedure)
C4031654|biopsy of bladder showed mesodermal mixed tumor
C4031654|biopsy of bladder showed mesodermal mixed tumor (procedure)
C4031619|biopsy of bladder showed small cell type (procedure)
C4031619|biopsy of bladder showed small cell type
C4031616|biopsy of bladder showed spindle cell type
C4031616|biopsy of bladder showed spindle cell type (procedure)
C4031738|biopsy of bladder showed carcinoma large cell with rhabdoid phenotype
C4031738|biopsy of bladder showed carcinoma large cell with rhabdoid phenotype (procedure)
C4031694|biopsy of bladder showed hodgkin's lymphoma
C4031694|biopsy of bladder showed hodgkin's lymphoma (procedure)
C4031660|biopsy of bladder showed lymphoma precursor cell lymphoblastic b-cell (procedure)
C4031660|biopsy of bladder showed lymphoma precursor cell lymphoblastic b-cell
C4031635|biopsy of bladder showed paraganglioma (procedure)
C4031635|biopsy of bladder showed paraganglioma
C4031631|biopsy of bladder showed sarcoma desmoplastic small round cell tumor (procedure)
C4031631|biopsy of bladder showed sarcoma desmoplastic small round cell tumor
C4031744|biopsy of bladder showed carcinoma glassy cell
C4031744|biopsy of bladder showed carcinoma glassy cell (procedure)
C4031740|biopsy of bladder showed carcinoma large cell (procedure)
C4031740|biopsy of bladder showed carcinoma large cell
C4031721|biopsy of bladder showed carcinoma squamous cell large cell, nonkeratinizing (procedure)
C4031721|biopsy of bladder showed carcinoma squamous cell large cell, nonkeratinizing
C4031720|biopsy of bladder showed carcinoma squamous cell microinvasive
C4031720|biopsy of bladder showed carcinoma squamous cell microinvasive (procedure)
C4031712|biopsy of bladder showed carcinoma transitional cell spindle cell
C4031712|biopsy of bladder showed carcinoma transitional cell spindle cell (procedure)
C4031710|biopsy of bladder showed carcinoma verrucous
C4031710|biopsy of bladder showed carcinoma verrucous (procedure)
C4031693|biopsy of bladder showed hodgkin's lymphoma granuloma (procedure)
C4031693|biopsy of bladder showed hodgkin's lymphoma granuloma
C4031692|biopsy of bladder showed hodgkin's lymphoma lymphocyte-rich (procedure)
C4031692|biopsy of bladder showed hodgkin's lymphoma lymphocyte-rich
C4031642|biopsy of bladder showed myosarcoma rhabdomyosarcoma pleomorphic, adult type (procedure)
C4031642|biopsy of bladder showed myosarcoma rhabdomyosarcoma pleomorphic, adult type
C4031639|biopsy of bladder showed non-hodgkin's lymphoma (procedure)
C4031639|biopsy of bladder showed non-hodgkin's lymphoma
C4031731|biopsy of bladder showed carcinoma schneiderian (procedure)
C4031731|biopsy of bladder showed carcinoma schneiderian
C4031727|biopsy of bladder showed carcinoma small cell fusiform cell (procedure)
C4031727|biopsy of bladder showed carcinoma small cell fusiform cell
C4031713|biopsy of bladder showed carcinoma transitional cell papillary
C4031713|biopsy of bladder showed carcinoma transitional cell papillary (procedure)
C4031699|biopsy of bladder showed fibrosarcoma infantile
C4031699|biopsy of bladder showed fibrosarcoma infantile (procedure)
C4031673|biopsy of bladder showed lymphoma follicular grade 2 (procedure)
C4031673|biopsy of bladder showed lymphoma follicular grade 2
C4031665|biopsy of bladder showed lymphoma mature t-cell
C4031665|biopsy of bladder showed lymphoma mature t-cell (procedure)
C4031646|biopsy of bladder showed myosarcoma rhabdomyosarcoma
C4031646|biopsy of bladder showed myosarcoma rhabdomyosarcoma (procedure)
C4031748|biopsy of bladder showed carcinoma cloacogenic
C4031748|biopsy of bladder showed carcinoma cloacogenic (procedure)
C4031747|biopsy of bladder showed carcinoma epithelioma
C4031747|biopsy of bladder showed carcinoma epithelioma (procedure)
C4031724|biopsy of bladder showed carcinoma squamous cell (procedure)
C4031724|biopsy of bladder showed carcinoma squamous cell
C4031711|biopsy of bladder showed carcinoma undifferentiated (procedure)
C4031711|biopsy of bladder showed carcinoma undifferentiated
C4031709|biopsy of bladder showed carcinoma with osteoclast-like giant cells
C4031709|biopsy of bladder showed carcinoma with osteoclast-like giant cells (procedure)
C4031696|biopsy of bladder showed giant cell type (procedure)
C4031696|biopsy of bladder showed giant cell type
C4031663|biopsy of bladder showed lymphoma mixed small and large cell, diffuse
C4031663|biopsy of bladder showed lymphoma mixed small and large cell, diffuse (procedure)
C4031649|biopsy of bladder showed myosarcoma leiomyosarcoma
C4031649|biopsy of bladder showed myosarcoma leiomyosarcoma (procedure)
C4031658|biopsy of bladder showed lymphoma small b-cell lymphocytic
C4031658|biopsy of bladder showed lymphoma small b-cell lymphocytic (procedure)
C4031643|biopsy of bladder showed myosarcoma rhabdomyosarcoma mixed type (procedure)
C4031643|biopsy of bladder showed myosarcoma rhabdomyosarcoma mixed type
C4031734|biopsy of bladder showed carcinoma pleomorphic
C4031734|biopsy of bladder showed carcinoma pleomorphic (procedure)
C4031723|biopsy of bladder showed carcinoma squamous cell adenoid (procedure)
C4031723|biopsy of bladder showed carcinoma squamous cell adenoid
C4031685|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis grade 1
C4031685|biopsy of bladder showed hodgkin's lymphoma nodular sclerosis grade 1 (procedure)
C4031629|biopsy of bladder showed sarcoma epithelioid
C4031629|biopsy of bladder showed sarcoma epithelioid (procedure)
C4031733|biopsy of bladder showed carcinoma polygonal cell
C4031733|biopsy of bladder showed carcinoma polygonal cell (procedure)
C4031718|biopsy of bladder showed carcinoma squamous cell spindle cell
C4031718|biopsy of bladder showed carcinoma squamous cell spindle cell (procedure)
C4031715|biopsy of bladder showed carcinoma transitional cell (procedure)
C4031715|biopsy of bladder showed carcinoma transitional cell
C4031708|biopsy of bladder showed carcinosarcoma
C4031708|biopsy of bladder showed carcinosarcoma (procedure)
C4031682|biopsy of bladder showed Hodgkin's lymphoma with lymphocytic depletion with diffuse fibrosis (procedure)
C4031682|biopsy of bladder showed Hodgkin's lymphoma with lymphocytic depletion with diffuse fibrosis
C4031689|biopsy of bladder showed hodgkin's lymphoma mixed cellularity (procedure)
C4031689|biopsy of bladder showed hodgkin's lymphoma mixed cellularity
C4031676|biopsy of bladder showed lymphoma composite hodgkin's and non-hodgkin's (procedure)
C4031676|biopsy of bladder showed lymphoma composite hodgkin's and non-hodgkin's
C4031650|biopsy of bladder showed myosarcoma angiomyosarcoma (procedure)
C4031650|biopsy of bladder showed myosarcoma angiomyosarcoma
C4031622|biopsy of bladder showed sarcoma small cell
C4031622|biopsy of bladder showed sarcoma small cell (procedure)
C0279681|squamous cell carcinoma of bladder (diagnosis)
C0279681|squamous cell carcinoma of bladder
C0279681|Bladder squamous cell carcinoma
C0279681|Squamous cell carcinoma of bladder (disorder)
C0279681|squamous cell carcinoma of the bladder
C0279681|bladder cancer, squamous cell carcinoma
C0279681|carcinoma, squamous cell, bladder
C0279681|Epidermoid Carcinoma of Bladder
C0279681|Epidermoid Carcinoma of Urinary Bladder
C0279681|Epidermoid Carcinoma of the Bladder
C0279681|Epidermoid Carcinoma of the Urinary Bladder
C0279681|Squamous Cell Carcinoma of Urinary Bladder
C0279681|Squamous Cell Carcinoma of the Urinary Bladder
C0279681|Urinary Bladder Epidermoid Carcinoma
C0279681|Urinary Bladder Squamous Cell Carcinoma
C0279681|Bladder Epidermoid Carcinoma
C1827293|Carcinoma of urinary bladder, invasive (disorder)
C1827293|Carcinoma of urinary bladder, invasive
C1827293|carcinoma of bladder, invasive
C1827293|carcinoma of bladder, invasive (diagnosis)
C1827293|bladder malignant carcinoma invasive
C1827293|Invasive bladder cancer
C0153616|Malignant neoplasm of other specified sites of bladder
C0153616|Malig neo bladder NEC
C0864967|Malignant neoplasm of bladder wall NOS
C1336527|Carcinoma of urinary bladder, superficial (disorder)
C1336527|Carcinoma of urinary bladder, superficial
C1336527|carcinoma of bladder, superficial (diagnosis)
C1336527|bladder malignant carcinoma superficial
C1336527|carcinoma of bladder, superficial
C1336527|Superficial Bladder Carcinoma
C1336527|Superficial Bladder Cancer
C1336527|Superficial Urinary Bladder Cancer
C1336527|Superficial Urinary Bladder Carcinoma
C0280218|stage, bladder cancer
C0280218|bladder cancer stage
C0279879|cellular diagnosis, bladder cancer
C0279879|bladder cancer cellular diagnosis
C1332561|Primary Bladder Lymphoma
C1332561|Lymphoma of Bladder
C1332561|Lymphoma of Urinary Bladder
C1332561|Lymphoma of the Bladder
C1332561|Lymphoma of the Urinary Bladder
C1332561|Urinary Bladder Lymphoma
C1332561|Bladder Lymphoma
C0862326|Malignant neoplasm of bladder recurrent
C0862326|Recurrent Malignant Bladder Neoplasm
C1276593|T3b: Bladder tumor invades perivesical tissue macroscopically (extravesicular mass) (finding)
C1276593|T3b: Bladder tumor invades perivesical tissue macroscopically (extravesicular mass)
C1276593|T3b: Bladder tumour invades perivesical tissue macroscopically (extravesicular mass)
C1276593|T3b: Bladder tumor invades perivesical tissue macroscopically (extravesicular mass) (tumor staging)
C1276588|T2b: Urinary bladder tumor invades deep muscle (outer half) (finding)
C1276588|T2b: Urinary bladder tumor invades deep muscle (outer half)
C1276588|T2b: Urinary bladder tumour invades deep muscle (outer half)
C1276588|T2b: Urinary bladder tumor invades deep muscle (outer half) (tumor staging)
C0349659|rhabdomyosarcoma of bladder (diagnosis)
C0349659|rhabdomyosarcoma of bladder
C0349659|Rhabdomyosarcoma of urinary bladder
C0349659|Rhabdomyosarcoma of bladder (disorder)
C1276587|T2a: Urinary bladder tumor invades superficial muscle (inner half) (finding)
C1276587|T2a: Urinary bladder tumor invades superficial muscle (inner half)
C1276587|T2a: Urinary bladder tumour invades superficial muscle (inner half)
C1276587|T2a: Urinary bladder tumor invades superficial muscle (inner half) (tumor staging)
C1276592|T3a: Bladder tumor invades perivesical tissue microscopically (finding)
C1276592|T3a: Bladder tumor invades perivesical tissue microscopically
C1276592|T3a: Bladder tumour invades perivesical tissue microscopically
C1276592|T3a: Bladder tumor invades perivesical tissue microscopically (tumor staging)
C1276591|T3: Urinary bladder tumor invades perivesical tissue (finding)
C1276591|T3: Urinary bladder tumor invades perivesical tissue
C1276591|T3: Urinary bladder tumour invades perivesical tissue
C1276591|T3: Urinary bladder tumor invades perivesical tissue (tumor staging)
C2212650|grade 3 follicular lymphoma of bladder
C2212650|grade 3 follicular lymphoma of bladder (diagnosis)
C2212657|NK/T-cell lymphoma of bladder
C2212657|NK/T-cell lymphoma of bladder (diagnosis)
C2212631|mixed cellularity Hodgkin's lymphoma of bladder (diagnosis)
C2212631|mixed cellularity Hodgkin's lymphoma of bladder
C2046544|Hodgkin's granuloma of bladder (diagnosis)
C2046544|Hodgkin's granuloma of bladder
C2046684|Hodgkin's sarcoma of bladder (diagnosis)
C2046684|Hodgkin's sarcoma of bladder
C2212640|small B-cell lymphocytic lymphoma of bladder
C2212640|small B-cell lymphocytic lymphoma of bladder (diagnosis)
C2212649|grade 2 follicular lymphoma of bladder
C2212649|grade 2 follicular lymphoma of bladder (diagnosis)
C2212651|marginal zone B-cell lymphoma of bladder
C2212651|marginal zone B-cell lymphoma of bladder (diagnosis)
C2212653|angioimmunoblastic T-cell lymphoma of bladder (diagnosis)
C2212653|angioimmunoblastic T-cell lymphoma of bladder
C2212653|angioimmunoblastic lymphadenopathy with dysproteinemia (AILD) of bladder
C2212662|Sezary syndrome of bladder
C2212662|Sezary syndrome of bladder (diagnosis)
C2046471|bladder malignant lymphoma Hodgkin's and non-Hodgkin's
C2046471|composite Hodgkin's and non-Hodgkin's lymphoma of bladder
C2046471|composite Hodgkin's and non-Hodgkin's lymphoma of bladder (diagnosis)
C2212644|large B-cell diffuse lymphoma of bladder (diagnosis)
C2212644|large B-cell diffuse lymphoma of bladder
C2113746|precursor T-cell lymphoblastic lymphoma of bladder (diagnosis)
C2113746|precursor T-cell lymphoblastic lymphoma of bladder
C2212614|mast cell sarcoma of bladder (diagnosis)
C2212614|mast cell sarcoma of bladder
C2212656|anaplastic large cell lymphoma, null cell type of bladder
C2212656|anaplastic large cell lymphoma, null cell type of bladder (diagnosis)
C2212641|lymphoplasmacytic lymphoma of bladder (diagnosis)
C2212641|lymphoplasmacytic lymphoma of bladder
C2212652|mature T-cell lymphoma of bladder (diagnosis)
C2212652|mature T-cell lymphoma of bladder
C2113675|precursor cell lymphoblastic lymphoma of bladder
C2113675|precursor cell lymphoblastic lymphoma of bladder (diagnosis)
C2212630|lymphocyte-rich Hodgkin's lymphoma of bladder (diagnosis)
C2212630|lymphocyte-rich Hodgkin's lymphoma of bladder
C2212642|mantle cell lymphoma of bladder
C2212642|mantle cell lymphoma of bladder (diagnosis)
C2212643|mixed small and large cell diffuse lymphoma of bladder
C2212643|mixed small and large cell diffuse lymphoma of bladder (diagnosis)
C2212647|follicular lymphoma of bladder (diagnosis)
C2212647|follicular lymphoma of bladder
C2212648|grade 1 follicular lymphoma of bladder
C2212648|grade 1 follicular lymphoma of bladder (diagnosis)
C2113606|precursor B-cell lymphoblastic lymphoma of bladder
C2113606|precursor B-cell lymphoblastic lymphoma of bladder (diagnosis)
C2212658|malignant histiocytosis of bladder (diagnosis)
C2212658|malignant histiocytosis of bladder
C0279565|Invasive Lobular Breast Carcinoma
C0279565|Lobular breast carcinoma invasive
C0279565|lobular invasive breast carcinoma
C0279565|carcinoma; infiltrating lobular, unspecified site
C0279565|infiltrating; lobular carcinoma, unspecified site
C0279565|Classic Invasive Lobular Carcinoma
C0279565|Infiltrating Lobular Adenocarcinoma
C0279565|Infiltrating Lobular Breast Carcinoma
C0279565|Infiltrating Lobular Carcinoma of Breast
C0279565|Infiltrating Lobular Carcinoma of the Breast
C0279565|Invasive Lobular Adenocarcinoma
C0279565|Invasive Lobular Carcinoma of Breast
C0279565|Invasive Lobular Carcinoma of the Breast
C0279565|Invasive Lobular Carcinoma, Classic Type
C0279565|Invasive Lobular Carcinoma
C0281267|bilateral breast cancer
C0281267|Bilateral Breast Carcinoma
C0242787|Malignant neoplasm of male breast
C0242787|malignant neoplasm of male breast (diagnosis)
C0242787|malignant male breast neoplasm
C0242787|malignant tumor of male breast
C0242787|Malignant neoplasm of male breast (disorder)
C0242787|Malignant neoplasm of male breast NOS
C0242787|Malignant neoplasm of male breast NOS (disorder)
C0242787|Breast neoplasm malignant male
C0242787|Malignant breast neoplasm male
C0242787|Malignant neoplasm of male breast, NOS
C0242787|Neoplasm malig;breast:M
C0242787|malignant neosplasm of the male breast
C0496812|Axillary tail of breast
C0496812|Malignant neoplasm of axillary tail of breast
C0496812|breast neoplasm malignant axillary tail
C0496812|malignant neoplasm of axillary tail of breast (diagnosis)
C0496812|Ca breast - axillary tail (disorder)
C0496812|Ca breast - axillary tail
C0496812|Malignant neoplasm of axillary tail of breast (disorder)
C0496807|Central portion of breast
C0496807|Malignant neoplasm of central portion of breast
C0496807|malignant neoplasm of central portion of breast (diagnosis)
C0496807|breast neoplasm malignant central portion
C0006142|Cancer, Breast
C0006142|Malignant neoplasm of breast
C0006142|Breast, unspecified
C0006142|Malignant neoplasm of breast, unspecified
C0006142|Breast cancer
C0006142|malignant neoplasm of breast (diagnosis)
C0006142|breast cancer (diagnosis)
C0006142|malignant breast neoplasm
C0006142|Ca breast
C0006142|cancer of breast
C0006142|malignant tumor of breast
C0006142|Malignant neoplasms of breast (C50)
C0006142|Ca breast - NOS
C0006142|Ca breast - NOS (disorder)
C0006142|[X]Malignant neoplasm of breast (disorder)
C0006142|[X]Malignant neoplasm of breast
C0006142|Breast--Cancer
C0006142|-- Breast Cancer
C0006142|Breast cancer stage unspecified
C0006142|Breast cancer NOS
C0006142|Breast tumor malignant
C0006142|Breast tumour malignant
C0006142|Mammary Cancer
C0006142|Cancer of the Breast
C0006142|Breast Carcinoma
C0006142|CA - Breast cancer
C0006142|Malignant tumour of breast
C0006142|Malignant tumor of breast (disorder)
C0006142|Malignant Breast Tumor
C0006142|Malignant Neoplasm of the Breast
C0006142|Malignant Tumor of the Breast
C0496809|Lower-inner quadrant of breast
C0496809|Malignant neoplasm of lower-inner quadrant of breast
C0496809|malignant neoplasm of lower inner quadrant of breast (diagnosis)
C0496809|breast neoplasm malignant lower inner quadrant
C0496809|malignant neoplasm of lower inner quadrant of breast
C0496809|Malignant neoplasm of breast lower inner quadrant (disorder)
C0496809|Malignant neoplasm of breast lower inner quadrant
C0496811|Lower-outer quadrant of breast
C0496811|Malignant neoplasm of lower-outer quadrant of breast
C0496811|malignant neoplasm of lower outer quadrant of breast
C0496811|malignant neoplasm of lower outer quadrant of breast (diagnosis)
C0496811|breast neoplasm malignant lower outer quadrant
C0496811|Malignant neoplasm of breast lower outer quadrant (disorder)
C0496811|Malignant neoplasm of breast lower outer quadrant
C0496806|Malignant neoplasm of nipple and areola
C0496806|Nipple and areola
C0496806|malignant neoplasm of nipple and areola (diagnosis)
C0496806|breast neoplasm malignant nipple / areola
C0348912|Malignant neoplasm overlapping breast site
C0348912|Overlapping lesion of breast
C0348912|Malignant neoplasm of overlapping sites of breast
C0348912|breast neoplasm malignant overlapping sites
C0348912|malignant neoplasm of overlapping sites of breast (diagnosis)
C0348912|Malignant neoplasm, overlapping lesion of breast
C0348912|Malignant neoplasm, overlapping lesion of breast (disorder)
C0496808|Malignant neoplasm of upper-inner quadrant of breast
C0496808|Upper-inner quadrant of breast
C0496808|breast neoplasm malignant upper inner quadrant
C0496808|malignant neoplasm of upper inner quadrant of breast
C0496808|malignant neoplasm of upper inner quadrant of breast (diagnosis)
C0496808|Malignant neoplasm of breast upper inner quadrant (disorder)
C0496808|Malignant neoplasm of breast upper inner quadrant
C0496810|Malignant neoplasm of upper-outer quadrant of breast
C0496810|Upper-outer quadrant of breast
C0496810|malignant neoplasm of upper outer quadrant of breast (diagnosis)
C0496810|breast neoplasm malignant upper outer quadrant
C0496810|malignant neoplasm of upper outer quadrant of breast
C0496810|Malignant neoplasm of breast upper outer quadrant (disorder)
C0496810|Malignant neoplasm of breast upper outer quadrant
C0678222|CARCINOMA OF BREAST
C0678222|Breast carcinoma
C0678222|carcinoma of breast (diagnosis)
C0678222|breast cancer diagnosis
C0678222|Carcinoma of breast NOS (disorder)
C0678222|Carcinoma of breast (disorder)
C0678222|Carcinoma of breast NOS
C0678222|Breast cancer, NOS
C0678222|breast cancer
C0678222|Cancer, Breast
C0678222|Breast carcinoma NOS
C0678222|Carcinoma breast
C0678222|CA - Carcinoma of breast
C0678222|Cancer of Breast
C0678222|Cancer of the Breast
C0678222|Mammary Carcinoma
C0678222|Carcinoma of the Breast
C2842134|Malignant neoplasm of breast of unspecified site
C0030185|Paget's Disease, Mammary
C0030185|Pagets Disease, Breast
C0030185|Disease, Mammary Paget
C0030185|Disease, Mammary Paget's
C0030185|Mammary Pagets Disease
C0030185|Pagets Disease, Mammary
C0030185|Paget's disease of breast
C0030185|Mammary Paget's Disease
C0030185|PAGETS DIS BREAST
C0030185|PAGET DIS MAMMARY
C0030185|PAGETS DIS MAMMARY
C0030185|MAMMARY PAGETS DIS
C0030185|PAGET DIS BREAST
C0030185|MAMMARY PAGET DIS
C0030185|Paget Disease of the Breast
C0030185|Paget's Disease of the Breast
C0030185|Paget's disease (mammary)
C0030185|Paget's disease of breast (diagnosis)
C0030185|Paget disease, mammary
C0030185|Paget's Disease, Mammary [Disease/Finding]
C0030185|Mammary Paget Disease
C0030185|Paget Disease of Breast
C0030185|Paget's Disease of the Nipple and Areola
C0030185|Paget's Disease of the Nipple
C0030185|Paget Disease, Breast
C0030185|Paget's disease, mammary (morphologic abnormality)
C0030185|breast; Paget
C0030185|breast; disorder, Paget
C0030185|Paget; breast
C2211687|breast neoplasm malignant small cell type
C2211687|malignant small cell neoplasm of breast (diagnosis)
C2211687|malignant small cell neoplasm of breast
C2011353|giant cell type neoplasm of breast
C2011353|giant cell type neoplasm of breast (diagnosis)
C2011353|breast neoplasm malignant giant cell type
C2018637|breast neoplasm malignant spindle cell type
C2018637|spindle cell type neoplasm of breast
C2018637|spindle cell type neoplasm of breast (diagnosis)
C2075596|breast neoplasm malignant clear cell type
C2075596|clear cell type neoplasm of breast (diagnosis)
C2075596|clear cell type neoplasm of breast
C0349667|sarcoma of breast
C0349667|sarcoma of breast (diagnosis)
C0349667|Breast sarcoma
C0349667|Sarcoma of breast (disorder)
C0349667|Sarcoma of the Breast
C2211725|myosarcoma of breast (diagnosis)
C2211725|myosarcoma of breast
C2211725|breast neoplasm malignant myosarcoma
C2007063|carcinosarcoma of breast
C2007063|carcinosarcoma of breast (diagnosis)
C2211730|malignant mesenchymoma of breast
C2211730|malignant mesenchymoma of breast (diagnosis)
C2211731|malignant hemangioendothelioma of breast
C2211731|malignant hemangioendothelioma of breast (diagnosis)
C0346154|Malignant Cystosarcoma Phyllodes of the Breast
C0346154|malignant phyllodes tumor of breast
C0346154|malignant phyllodes tumor of breast (diagnosis)
C0346154|Malignant cystosarcoma phyllodes of breast
C0346154|Malignant phyllodes tumour of breast
C0346154|Malignant phyllodes tumor of breast (disorder)
C0346154|Malignant Breast Phyllodes Neoplasm
C0346154|Malignant Mammary Phyllodes Neoplasm
C0346154|Malignant Mammary Phyllodes Tumor
C0346154|Malignant Phyllodes Breast Neoplasm
C0346154|Malignant Phyllodes Neoplasm of Breast
C0346154|Malignant Phyllodes Neoplasm of the Breast
C0346154|Malignant Phyllodes Tumor of the Breast
C0346154|Malignant Breast Phyllodes Tumor
C2211733|malignant granular cell tumor of breast
C2211733|malignant granular cell tumor of breast (diagnosis)
C2211755|malignant plasmacytoma of breast (diagnosis)
C2211755|malignant plasmacytoma of breast
C2211757|malignant mastocytosis of breast
C2211757|malignant mastocytosis of breast (diagnosis)
C2216702|malignant neoplasm of breast staging (diagnosis)
C2216702|malignant neoplasm of breast staging
C2216702|malignant breast neoplasm staging
C2216702|malignant tumor of breast staging
C2216702|breast cancer staging
C2216702|stage, breast cancer
C2216702|breast cancer stage
C0677776|Hereditary Breast and Ovarian Cancer Syndrome
C0677776|HBOC Syndromes
C0677776|Syndrome, HBOC
C0677776|Syndromes, HBOC
C0677776|HBOC Syndrome
C0677776|Hereditary Breast and Ovarian Cancer Syndrome [Disease/Finding]
C0677776|Familial Breast and Ovarian Cancer Syndrome
C0677776|familial breast-ovarian cancer syndrome
C0677776|familial breast-ovarian cancer syndrome (diagnosis)
C0677776|hereditary breast/ovarian cancer (BRCA1, BRCA2)
C0677776|Familial Breast/Ovarian Cancer (BRCA1, BRCA2)
C0677776|Hereditary Breast and Ovarian Cancer
C0858252|adenocarcinoma of breast (diagnosis)
C0858252|adenocarcinoma of breast
C0858252|breast adenocarcinoma
C0858252|Adenocarcinoma of the Breast
C1332630|fibrosarcoma of breast (diagnosis)
C1332630|fibrosarcoma of breast
C1332630|Fibrosarcoma of the Breast
C1332630|Breast Fibrosarcoma
C2062549|epithelioma of nipple (diagnosis)
C2062549|epithelioma of nipple
C2062549|breast nipple epithelioma
C1332632|liposarcoma of breast (diagnosis)
C1332632|liposarcoma of breast
C1332632|Liposarcoma of the Breast
C1332632|Breast Liposarcoma
C0235653|Malignant neoplasm of breast (female), unspecified
C0235653|Malignant neoplasm of female breast
C0235653|malignant neoplasm of female breast (diagnosis)
C0235653|cancer of female breast
C0235653|malignant female breast neoplasm
C0235653|malignant tumor of female breast
C0235653|Malign neopl breast NOS
C0235653|Malignant neoplasm of female breast (disorder)
C0235653|Malignant neoplasm of female breast NOS
C0235653|Malignant neoplasm of female breast NOS (disorder)
C0235653|Breast cancer female
C0235653|Female breast cancer
C0235653|Malignant neoplasm of female breast, unspecified
C0235653|Breast neoplasm malignant female
C0235653|Breast cancer female NOS
C0235653|Breast cancer, female
C0235653|Malignant neoplasm of female breast, NOS
C0235653|Neoplasm malig;breast;F
C0235653|malignant neosplasm of the female breast
C2211688|malignant epithelioma of breast
C2211688|malignant epithelioma of breast (diagnosis)
C2111593|large cell carcinoma of breast
C2111593|large cell carcinoma of breast (diagnosis)
C1511316|large cell neuroendocrine carcinoma of breast
C1511316|large cell neuroendocrine carcinoma of breast (diagnosis)
C1511316|Breast Large Cell Neuroendocrine Carcinoma
C2111594|large cell carcinoma of breast with rhabdoid phenotype (diagnosis)
C2111594|breast malignant carcinoma large cell w/ rhabdoid phenotype
C2111594|large cell carcinoma of breast with rhabdoid phenotype
C2012071|glassy cell carcinoma of breast
C2012071|glassy cell carcinoma of breast (diagnosis)
C1336854|undifferentiated carcinoma of breast
C1336854|undifferentiated carcinoma of breast (diagnosis)
C2211689|anaplastic carcinoma of breast (diagnosis)
C2211689|anaplastic carcinoma of breast
C2211689|Anaplastic Breast Carcinoma
C1514169|pleomorphic carcinoma of breast
C1514169|pleomorphic carcinoma of breast (diagnosis)
C1514169|Pleomorphic Breast Carcinoma
C2011243|giant cell carcinoma of breast (diagnosis)
C2011243|giant cell carcinoma of breast
C2018385|spindle cell carcinoma of breast
C2018385|spindle cell carcinoma of breast (diagnosis)
C2011208|giant cell and spindle cell carcinoma of breast (diagnosis)
C2011208|giant cell and spindle cell carcinoma of breast
C2142913|pseudosarcomatous carcinoma of breast
C2142913|pseudosarcomatous carcinoma of breast (diagnosis)
C2111795|polygonal cell carcinoma of breast (diagnosis)
C2111795|polygonal cell carcinoma of breast
C2007022|carcinoma of breast with osteoclast-like giant cells (diagnosis)
C2007022|carcinoma of breast with osteoclast-like giant cells
C2007022|breast carcinoma with osteoclast-like giant cells
C3812899|papillary carcinoma of breast
C3812899|papillary carcinoma of breast (diagnosis)
C3812899|Papillary carcinoma of the breast (morphologic abnormality)
C3812899|Papillary carcinoma of the breast
C3812899|Papillary breast carcinoma
C2033277|papillary squamous cell carcinoma of breast (diagnosis)
C2033277|papillary squamous cell carcinoma of breast
C2189332|verrucous carcinoma of breast (diagnosis)
C2189332|verrucous carcinoma of breast
C1336079|Primary Squamous Cell Carcinoma of Breast
C1336079|Primary Squamous Cell Breast Carcinoma
C1336079|Primary Squamous Cell Carcinoma of the Breast
C1336079|squamous cell carcinoma of breast (diagnosis)
C1336079|squamous cell carcinoma of breast
C1336079|SCC of Breast
C1336079|SCC of the Breast
C1336079|Squamous Breast Carcinoma
C1336079|Squamous Carcinoma of Breast
C1336079|Squamous Carcinoma of the Breast
C1336079|Squamous Cell Breast Carcinoma
C1336079|Squamous Cell Carcinoma of the Breast
C2109290|keratinizing squamous cell carcinoma of breast
C2109290|keratinizing squamous cell carcinoma of breast (diagnosis)
C2211690|nonkeratinizing large cell squamous carcinoma cell of breast
C2211690|nonkeratinizing large cell squamous carcinoma cell of breast (diagnosis)
C2211690|breast malignant carcinoma squamous cell large cell nonkeratinizing
C2018534|spindle cell squamous cell carcinoma of breast
C2018534|spindle cell squamous cell carcinoma of breast (diagnosis)
C2211692|adenoid squamous cell carcinoma of breast (diagnosis)
C2211692|adenoid squamous cell carcinoma of breast
C2211693|microinvasive squamous cell carcinoma of breast (diagnosis)
C2211693|microinvasive squamous cell carcinoma of breast
C2019466|squamous cell carcinoma of breast with horn formation
C2019466|squamous cell carcinoma of breast with horn formation (diagnosis)
C2019466|squamous cell carcinoma with horn formation of breast
C1332638|Oat Cell Carcinoma of Breast
C1332638|small cell carcinoma of breast
C1332638|small cell carcinoma of breast (diagnosis)
C1332638|Mammary Small Cell Carcinoma
C1332638|Oat Cell Carcinoma of the Breast
C1332638|Small Cell Carcinoma of the Breast
C1332638|Small Cell Neuroendocrine Carcinoma of Breast
C1332638|Small Cell Neuroendocrine Carcinoma of the Breast
C1332638|Breast Small Cell Carcinoma
C2009874|fusiform type small cell carcinoma of breast (diagnosis)
C2009874|fusiform type small cell carcinoma of breast
C1332167|adenoid cystic carcinoma of breast
C1332167|adenoid cystic carcinoma of breast (diagnosis)
C1332167|Adenoid cystic breast carcinoma
C1332167|Adenocystic Breast Carcinoma
C1332167|Adenocystic Carcinoma of Breast
C1332167|Adenocystic Carcinoma of the Breast
C1332167|Adenoid Cystic Carcinoma of the Breast
C1332167|Mammary Adenocystic Carcinoma
C2007046|carcinoma simplex of breast
C2007046|carcinoma simplex of breast (diagnosis)
C1517894|lipid-rich carcinoma of breast
C1517894|lipid-rich carcinoma of breast (diagnosis)
C1517894|Lipid Secreting Breast Carcinoma
C1517894|Lipid-Rich Breast Carcinoma
C2012538|granular cell carcinoma of breast (diagnosis)
C2012538|granular cell carcinoma of breast
C1335964|signet ring cell carcinoma of breast
C1335964|signet ring cell carcinoma of breast (diagnosis)
C1335964|Mammary Signet Ring Cell Carcinoma
C1335964|Primary Mammary Signet Ring Cell Carcinoma
C1335964|Primary SRC Breast Carcinoma
C1335964|Primary SRC Carcinoma of Breast
C1335964|Primary SRC Carcinoma of the Breast
C1335964|Primary Signet Ring Cell Breast Carcinoma
C1335964|Primary Signet Ring Cell Carcinoma of Breast
C1335964|Primary Signet Ring Cell Carcinoma of the Breast
C1335964|SRC Breast Carcinoma
C1335964|SRC Carcinoma of Breast
C1335964|SRC Carcinoma of the Breast
C1335964|Signet Ring Cell Breast Carcinoma
C1335964|Signet Ring Cell Carcinoma of the Breast
C1334002|comedocarcinoma of breast (diagnosis)
C1334002|comedocarcinoma of breast
C1334002|High Grade Ductal Breast Carcinoma In Situ
C1334002|comedo carcinoma
C1334002|DIN 3
C1334002|Ductal intraepithelial neoplasia 3
C1334002|DCIS Grade 3
C1334002|Ductal Intraepithelial Neoplasia, Grade 3
C1334002|High-Grade DCIS of Breast
C1334002|High-Grade DCIS of the Breast
C1334002|High-Grade Ductal Carcinoma In Situ of Breast
C1334002|Breast Comedocarcinoma
C0334371|Cystic Hypersecretory Carcinoma of Breast
C0334371|Cystic Hypersecretory Breast Carcinoma
C0334371|Secretory Carcinoma
C0334371|Cystic Hypersecretory Carcinoma of the Breast
C0334371|secretory carcinoma of breast (diagnosis)
C0334371|secretory carcinoma of breast
C0334371|hypersecretory cystic carcinoma of breast (diagnosis)
C0334371|hypersecretory cystic carcinoma of breast
C0334371|Secretory breast carcinoma
C0334371|Juvenile carcinoma of the breast
C0334371|Secretory carcinoma of the breast
C0334371|Juvenile carcinoma of the breast (morphologic abnormality)
C0334371|Infiltrating Cystic Hypersecretory Duct Breast Carcinoma
C0334371|Invasive Cystic Hypersecretory Duct Breast Carcinoma
C0334371|Juvenile Breast Carcinoma
C0334371|Juvenile Carcinoma of Breast
C0334371|Juvenile Secretory Breast Carcinoma
C0334371|Juvenile Secretory Carcinoma of Breast
C0334371|Juvenile Secretory Carcinoma of the Breast
C0334376|intracystic carcinoma of breast (diagnosis)
C0334376|intracystic carcinoma of breast
C0334376|Intracystic Papillary Breast Carcinoma
C0334376|[M] Intracystic carcinoma NOS
C0334376|[M] Intracystic carcinoma NOS (morphologic abnormality)
C0334376|Intracystic carcinoma
C0334376|Intracystic carcinoma (morphologic abnormality)
C0334376|Intracystic papillary adenocarcinoma
C0334376|Intracystic carcinoma, NOS
C0334376|Intracystic Breast Carcinoma
C0334376|Noninfiltrating Intracystic Breast Carcinoma
C0860580|medullary carcinoma of breast (diagnosis)
C0860580|medullary carcinoma of breast
C0860580|medullary breast carcinoma
C0860580|Infiltrating Medullary Carcinoma of Breast
C0860580|Infiltrating Medullary Carcinoma of the Breast
C0860580|Invasive Medullary Breast Carcinoma
C0860580|Invasive Medullary Carcinoma of Breast
C0860580|Invasive Medullary Carcinoma of the Breast
C0860580|Medullary Breast Carcinoma with Lymphoid Stroma
C0860580|Medullary Carcinoma of the Breast
C2211694|medullary carcinoma with lymphoid stroma of breast (diagnosis)
C2211694|medullary carcinoma with lymphoid stroma of breast
C1879758|Atypical Medullary Breast Carcinoma
C1879758|Infiltrating Ductal Breast Carcinoma with Medullary Features
C1879758|atypical medullary carcinoma of breast (diagnosis)
C1879758|atypical medullary carcinoma of breast
C2182973|desmoplastic type ductal carcinoma of breast
C2182973|desmoplastic type ductal carcinoma of breast (diagnosis)
C2076522|infiltrating ductal and lobular carcinoma of breast (diagnosis)
C2076522|infiltrating ductal and lobular carcinoma of breast
C2146658|acinar cell carcinoma of breast (diagnosis)
C2146658|acinar cell carcinoma of breast
C2146670|acinar cell cystadenocarcinoma of breast
C2146670|acinar cell cystadenocarcinoma of breast (diagnosis)
C1510796|adenosquamous carcinoma of breast
C1510796|adenosquamous carcinoma of breast (diagnosis)
C1510796|Adenosquamous Breast Carcinoma
C2211695|epithelial-myoepithelial carcinoma of breast (diagnosis)
C2211695|epithelial-myoepithelial carcinoma of breast
C1334708|metaplastic carcinoma of breast (diagnosis)
C1334708|metaplastic carcinoma of breast
C1334708|Metaplastic breast carcinoma
C1334708|Metaplastic Carcinoma of the Breast
C2211696|scirrhous adenocarcinoma of breast
C2211696|scirrhous adenocarcinoma of breast (diagnosis)
C2037312|superficial spreading adenocarcinoma of breast
C2037312|superficial spreading adenocarcinoma of breast (diagnosis)
C2211697|basal cell adenocarcinoma of breast
C2211697|basal cell adenocarcinoma of breast (diagnosis)
C2145023|trabecular adenocarcinoma of breast (diagnosis)
C2145023|trabecular adenocarcinoma of breast
C2033109|papillary adenocarcinoma of breast (diagnosis)
C2033109|papillary adenocarcinoma of breast
C2211698|apocrine adenocarcinoma of breast (diagnosis)
C2211698|apocrine adenocarcinoma of breast
C2211699|intraductal papillary adenocarcinoma of breast with invasion
C2211699|intraductal papillary adenocarcinoma of breast with invasion (diagnosis)
C2211700|mixed cell adenocarcinoma of breast (diagnosis)
C2211700|mixed cell adenocarcinoma of breast
C2211701|polymorphous low grade adenocarcinoma of breast (diagnosis)
C2211701|polymorphous low grade adenocarcinoma of breast
C2075524|clear cell adenocarcinoma of breast (diagnosis)
C2075524|clear cell adenocarcinoma of breast
C2211702|mucinous adenocarcinoma of breast (diagnosis)
C2211702|mucinous adenocarcinoma of breast
C2211703|mucin-producing adenocarcinoma of breast (diagnosis)
C2211703|mucin-producing adenocarcinoma of breast
C2211704|breast adenocarcinoma with metaplasia
C2211704|adenocarcinoma of breast with metaplasia (diagnosis)
C2211704|adenocarcinoma of breast with metaplasia
C1332613|adenocarcinoma of breast with squamous metaplasia (diagnosis)
C1332613|adenocarcinoma of breast with squamous metaplasia
C1332613|breast adenocarcinoma with squamous metaplasia
C1332613|Adenoacanthoma of Breast
C1332613|Adenoacanthoma of the Breast
C1332613|Adenocarcinoma of the Breast with Squamous Metaplasia
C1332613|Breast Adenoacanthoma
C2211705|adenocarcinoma with cartilaginous or osseous metaplasia of breast
C2211705|adenocarcinoma of breast with cartilaginous and osseous metaplasia
C2211705|breast adenocarcinoma with cartilaginous or osseous metaplasia
C2211705|adenocarcinoma of breast with cartilaginous and osseous metaplasia (diagnosis)
C2211705|breast adenocarcinoma with cartilaginous and osseous metaplasia
C1511281|breast adenocarcinoma with spindle cell metaplasia
C1511281|adenocarcinoma of breast with spindle cell metaplasia
C1511281|adenocarcinoma of breast with spindle cell metaplasia (diagnosis)
C2211706|adenocarcinoma of breast with apocrine metaplasia
C2211706|breast adenocarcinoma with apocrine metaplasia
C2211706|adenocarcinoma of breast with apocrine metaplasia (diagnosis)
C2211707|adenocarcinoma of breast with neuroendocrine differentiation (diagnosis)
C2211707|adenocarcinoma of breast with neuroendocrine differentiation
C2211707|breast adenocarcinoma with neuroendocrine differentiation
C2170817|tubular adenocarcinoma of breast (diagnosis)
C2170817|tubular adenocarcinoma of breast
C2211708|alveolar adenocarcinoma of breast
C2211708|alveolar adenocarcinoma of breast (diagnosis)
C2163806|cystadenocarcinoma of breast (diagnosis)
C2163806|cystadenocarcinoma of breast
C2211732|malignant epithelioid hemangioendothelioma of breast
C2211732|malignant epithelioid hemangioendothelioma of breast (diagnosis)
C0334386|Paget's disease and infiltrating duct carcinoma of breast
C0334386|Paget's disease and infiltrating duct carcinoma of breast (diagnosis)
C0334386|Paget disease and infiltrating duct carcinoma of breast
C0334386|Paget's disease and infiltrating duct carcinoma of breast (morphologic abnormality)
C0279566|Paget Disease and Intraductal Carcinoma of the Breast
C0279566|Paget's Disease and Intraductal Carcinoma of the Breast
C0279566|Paget's disease and intraductal carcinoma of breast (diagnosis)
C0279566|Paget's disease and intraductal carcinoma of breast
C0279566|Paget disease and intraductal carcinoma of breast
C0279566|Paget's disease and intraductal carcinoma of breast (disorder)
C0279566|[M]Paget's disease and intraductal carcinoma of breast
C0279566|[M] Paget's disease and intraductal carcinoma of breast
C0279566|Paget's disease and intraductal carcinoma of breast (morphologic abnormality)
C0279566|Paget's disease of the breast with intraductal carcinoma
C0279566|Paget's Disease of Breast with Intraductal Carcinoma
C2211718|malignant solitary fibrous tumor of breast
C2211718|malignant solitary fibrous tumor of breast (diagnosis)
C2211729|embryonal carcinosarcoma of breast
C2211729|embryonal carcinosarcoma of breast (diagnosis)
C1518167|malignant myoepithelioma of breast (diagnosis)
C1518167|malignant myoepithelioma of breast
C1518167|Breast Myoepithelial Carcinoma
C1518167|Malignant Breast Myoepithelioma
C2216703|malignant neoplasm of breast TNM staging
C2216703|malignant neoplasm of breast TNM staging (diagnosis)
C2216703|malignant breast neoplasm TNM staging
C2216703|malignant tumor of breast TNM staging
C2216703|breast cancer TNM staging
C2216694|malignant neoplasm of breast stage 0
C2216694|malignant neoplasm of breast stage 0 (diagnosis)
C2216694|malignant breast neoplasm stage 0
C2216694|breast cancer stage 0
C2216694|malignant tumor of breast stage 0
C2216695|malignant neoplasm of breast stage I (diagnosis)
C2216695|malignant neoplasm of breast stage I
C2216695|malignant breast neoplasm stage I
C2216695|malignant tumor of breast stage I
C2216695|breast cancer stage I
C2216695|Stage I Breast Cancer
C2216695|Stage I Breast Cancer AJCC v7
C2216696|malignant neoplasm of breast stage IIa (diagnosis)
C2216696|malignant neoplasm of breast stage IIa
C2216696|malignant breast neoplasm stage IIa
C2216696|breast cancer stage IIa
C2216696|malignant tumor of breast stage IIa
C2216697|malignant neoplasm of breast stage IIb (diagnosis)
C2216697|malignant neoplasm of breast stage IIb
C2216697|malignant breast neoplasm stage IIb
C2216697|malignant tumor of breast stage IIb
C2216697|breast cancer stage IIb
C2216698|malignant neoplasm of breast stage IIIa (diagnosis)
C2216698|malignant neoplasm of breast stage IIIa
C2216698|malignant breast neoplasm stage IIIa
C2216698|malignant tumor of breast stage IIIa
C2216698|breast cancer stage IIIa
C2216699|malignant neoplasm of breast stage IIIb (diagnosis)
C2216699|malignant neoplasm of breast stage IIIb
C2216699|malignant breast neoplasm stage IIIb
C2216699|breast cancer stage IIIb
C2216699|malignant tumor of breast stage IIIb
C2216700|malignant neoplasm of breast stage IIIc
C2216700|malignant neoplasm of breast stage IIIc (diagnosis)
C2216700|malignant breast neoplasm stage IIIc
C2216700|malignant tumor of breast stage IIIc
C2216700|breast cancer stage IIIc
C2216700|Stage IIIC Breast Cancer AJCC v6
C2216700|Stage IIIC Breast Carcinoma AJCC v6
C2216700|stage IIIC breast cancer
C2216701|malignant neoplasm of breast stage IV
C2216701|malignant neoplasm of breast stage IV (diagnosis)
C2216701|malignant breast neoplasm stage IV
C2216701|breast cancer stage IV
C2216701|malignant tumor of breast stage IV
C2062550|neurosarcoma of breast (diagnosis)
C2062550|neurosarcoma of breast
C2211754|malignant histiocytosis of breast (diagnosis)
C2211754|malignant histiocytosis of breast
C3665394|Malignant neoplasm of skin of breast
C3665394|Malignant neoplasm of skin of breast (disorder)
C3665394|skin neoplasm malignant breast
C3665394|malignant skin neoplasm of breast
C3665394|malignant skin neoplasm of breast (diagnosis)
C3469450|susceptibility to familial breast-ovarian cancer syndrome (diagnosis)
C3469450|susceptibility to familial breast-ovarian cancer syndrome
C3469522|breast cancer susceptibility (diagnosis)
C3469522|breast cancer susceptibility
C3469522|BREAST CANCER, SUSCEPTIBILITY TO
C1306469|Primary malignant neoplasm of male breast (diagnosis)
C1306469|breast neoplasm malignant male primary
C1306469|Primary malignant neoplasm of male breast
C1306469|Primary malignant neoplasm of male breast (disorder)
C0559019|Ca breast-upper,inner quadrant (disorder)
C0559019|Ca breast-upper,inner quadrant
C0559020|Ca breast-upper,outer quadrant
C0559020|Ca breast-upper,outer quadrant (disorder)
C1304708|Primary malignant neoplasm of female breast
C1304708|breast neoplasm malignant female primary
C1304708|Primary malignant neoplasm of female breast (diagnosis)
C1304708|Primary malignant neoplasm of female breast (disorder)
C0346860|malignant male breast tissue neoplasm
C0346860|malignant male breast ectopic tissue neoplasm
C0346860|malignant male breast neoplasm of ectopic breast tissue
C0346860|malignant neoplasm of ectopic tissue of male breast
C0346860|malignant male breast neoplasm of ectopic breast tissue (diagnosis)
C0346860|Malignant neoplasm of ectopic site of male breast
C0346860|Malignant neoplasm of ectopic site of male breast (disorder)
C0559021|Ca breast-lower,outer quadrant
C0559021|Ca breast-lower,outer quadrant (disorder)
C0559062|Ca breast-lower,inner quadrant
C0559062|Ca breast-lower,inner quadrant (disorder)
C0948966|Malignant nipple neoplasm female
C0948966|breast neoplasm malignant female nipple
C0948966|malignant neoplasm of female nipple (diagnosis)
C0948966|malignant neoplasm of female nipple
C0948966|Malignant neoplasm of nipple of female breast
C0948966|Female Malignant Nipple Neoplasm
C0346858|Malignant neoplasm of areola of male breast
C0346858|Malignant neoplasm of areola of male breast (disorder)
C0346858|breast neoplasm malignant male areola primary
C0346858|malignant neoplasm of areola of male breast (diagnosis)
C0346858|primary malignant neoplasm of areola of male breast (diagnosis)
C0346858|breast neoplasm malignant male areola
C0346858|primary malignant neoplasm of areola of male breast
C0346858|Primary malignant neoplasm of areola of male breast (disorder)
C0346857|Malignant neoplasm of nipple of male breast
C0346857|Malignant neoplasm of nipple of male breast (disorder)
C0346857|breast neoplasm malignant male nipple
C0346857|malignant neoplasm of nipple of male breast (diagnosis)
C0346857|primary malignant neoplasm of nipple of male breast (diagnosis)
C0346857|breast neoplasm malignant male nipple primary
C0346857|primary malignant neoplasm of nipple of male breast
C0346857|Primary malignant neoplasm of nipple of male breast (disorder)
C0346862|Malignant neoplasm of areola of female breast
C0346862|Malignant neoplasm of areola of female breast (disorder)
C0346862|breast neoplasm malignant female areola
C0346862|breast neoplasm malignant female areola primary
C0346862|Primary malignant neoplasm of areola of female breast
C0346862|Primary malignant neoplasm of areola of female breast (diagnosis)
C0346862|malignant neoplasm of areola of female breast (diagnosis)
C0346862|Primary malignant neoplasm of areola of female breast (disorder)
C3649897|malignant breast tissue neoplasm
C3649897|malignant breast tissue neoplasm (diagnosis)
C3649897|breast neoplasm malignant breast tissue
C1299258|Primary malignant neoplasm of breast
C1299258|Primary malignant neoplasm of breast (diagnosis)
C1299258|breast neoplasm malignant primary
C1299258|Primary malignant neoplasm of breast (disorder)
C2216720|malignant neoplasm of breast TNM staging regional lymph node (N) NX (diagnosis)
C2216720|malignant neoplasm of breast TNM staging regional lymph node (N) NX
C2216720|malignant breast neoplasm NX
C2216720|breast cancer TNM staging regional lymph node (N) NX
C2216720|malignant tumor of breast TNM staging regional lymph node (N) NX
C2216707|malignant neoplasm of breast TNM staging distant metastasis (M) MX (diagnosis)
C2216707|malignant neoplasm of breast TNM staging distant metastasis (M) MX
C2216707|malignant breast neoplasm MX
C2216707|malignant tumor of breast TNM staging distant metastasis (M) MX
C2216707|breast cancer TNM staging distant metastasis (M) MX
C2216718|malignant neoplasm of breast TNM staging regional lymph node (N) N2
C2216718|malignant neoplasm of breast TNM staging regional lymph node (N) N2 (diagnosis)
C2216718|malignant breast neoplasm N2
C2216718|malignant tumor of breast TNM staging regional lymph node (N) N2
C2216718|breast cancer TNM staging regional lymph node (N) N2
C2216716|malignant neoplasm of breast TNM staging regional lymph node (N) N0 (diagnosis)
C2216716|malignant neoplasm of breast TNM staging regional lymph node (N) N0
C2216716|malignant breast neoplasm N0
C2216716|malignant tumor of breast TNM staging regional lymph node (N) N0
C2216716|breast cancer TNM staging regional lymph node (N) N0
C2216719|malignant neoplasm of breast TNM staging regional lymph node (N) N3
C2216719|malignant neoplasm of breast TNM staging regional lymph node (N) N3 (diagnosis)
C2216719|malignant breast neoplasm N3
C2216719|breast cancer TNM staging regional lymph node (N) N3
C2216719|malignant tumor of breast TNM staging regional lymph node (N) N3
C2216721|malignant neoplasm of breast TNM staging regional lymph nodes (N)
C2216721|malignant neoplasm of breast TNM staging regional lymph nodes (N) (diagnosis)
C2216721|malignant breast neoplasm TNM staging of regional lymph nodes (N)
C2216721|breast cancer TNM staging regional lymph nodes (N)
C2216721|malignant tumor of breast TNM staging regional lymph nodes (N)
C2216706|malignant neoplasm of breast TNM staging distant metastasis (M) M1 (diagnosis)
C2216706|malignant neoplasm of breast TNM staging distant metastasis (M) M1
C2216706|malignant breast neoplasm M1
C2216706|breast cancer TNM staging distant metastasis (M) M1
C2216706|malignant tumor of breast TNM staging distant metastasis (M) M1
C2216705|malignant neoplasm of breast TNM staging distant metastasis (M) M0
C2216705|malignant neoplasm of breast TNM staging distant metastasis (M) M0 (diagnosis)
C2216705|malignant breast neoplasm M0
C2216705|breast cancer TNM staging distant metastasis (M) M0
C2216705|malignant tumor of breast TNM staging distant metastasis (M) M0
C2216717|malignant neoplasm of breast TNM staging regional lymph node (N) N1 (diagnosis)
C2216717|malignant neoplasm of breast TNM staging regional lymph node (N) N1
C2216717|malignant breast neoplasm N1
C2216717|malignant tumor of breast TNM staging regional lymph node (N) N1
C2216717|breast cancer TNM staging regional lymph node (N) N1
C2216704|malignant neoplasm of breast TNM staging distant metastasis (M)
C2216704|malignant neoplasm of breast TNM staging distant metastasis (M) (diagnosis)
C2216704|malignant breast neoplasm TNM staging of distant metastasis (M)
C2216704|breast cancer TNM staging distant metastasis (M)
C2216704|malignant tumor of breast TNM staging distant metastasis (M)
C3694291|metastasis from malignant neoplasm of breast
C3694291|metastasis from malignant neoplasm of breast (diagnosis)
C0346153|Breast Cancer, Familial
C0346153|familial breast cancer
C0346153|familial breast cancer (diagnosis)
C0346153|Familial cancer of breast
C0346153|Familial cancer of breast (disorder)
C0346153|Familial Cancer of the Breast
C0346153|Hereditary Breast Cancer
C0346153|Hereditary Breast Carcinoma
C0346153|Familial Breast Carcinoma
C1562029|breast neoplasm malignant hormone receptor positive
C1562029|Hormone receptor positive malignant neoplasm of breast
C1562029|Hormone receptor positive malignant neoplasm of breast (diagnosis)
C1562029|Hormone receptor positive malignant neoplasm of breast (disorder)
C3695123|local recurrence of malignant breast neoplasm
C3695123|local recurrence of malignant breast neoplasm (diagnosis)
C3695123|breast neoplasm malignant local recurrence
C3695122|breast neoplasm malignant staging tnm pathologic (pn)
C3695122|malignant breast neoplasm pathologic (pN) staging
C3695122|malignant breast neoplasm pathologic (pN) staging (diagnosis)
C0349669|malignant lymphoma of breast
C0349669|Malignant lymphoma of breast (disorder)
C4031559|biopsy of breast showed carcinoma medullary atypical
C4031559|biopsy of breast showed atypical medullary carcinoma
C4031559|biopsy of breast showed atypical medullary carcinoma (procedure)
C4031545|biopsy of breast showed signet ring cell carcinoma (procedure)
C4031545|biopsy of breast showed signet ring cell carcinoma
C4031545|biopsy of breast showed carcinoma signet ring cell
C4031466|biopsy of breast showed precursor cell lymphoblastic lymphoma
C4031466|biopsy of breast showed lymphoma precursor cell lymphoblastic
C4031466|biopsy of breast showed precursor cell lymphoblastic lymphoma (procedure)
C4031512|biopsy of breast showed epithelioid hemangioendothelioma
C4031512|biopsy of breast showed hemangioendothelioma epithelioid
C4031512|biopsy of breast showed epithelioid hemangioendothelioma (procedure)
C4031503|biopsy of breast showed Hodgkin's lymphoma with grade 1 nodular sclerosis
C4031503|biopsy of breast showed Hodgkin's lymphoma with grade 1 nodular sclerosis (procedure)
C4031503|biopsy of breast showed Hodgkin's lymphoma with nodular sclerosis grade 1
C4031490|biopsy of breast showed pleomorphic liposarcoma (procedure)
C4031490|biopsy of breast showed liposarcoma pleomorphic
C4031490|biopsy of breast showed pleomorphic liposarcoma
C4031482|biopsy of breast showed lymphoma composite Hodgkin's and non-Hodgkin's
C4031482|biopsy of breast showed lymphoma composite Hodgkin's and non-Hodgkin's (procedure)
C4031526|biopsy of breast showed duct carcinoma, desmoplastic type
C4031526|biopsy of breast showed duct carcinoma, desmoplastic type (procedure)
C4031526|biopsy of breast showed carcinoma duct, desmoplastic type
C4031523|biopsy of breast showed fibrosarcoma (procedure)
C4031523|biopsy of breast showed fibrosarcoma
C4031505|biopsy of breast showed Hodgkin's lymphoma with lymphocytic depletion with diffuse fibrosis
C4031505|biopsy of breast showed Hodgkin's lymphoma with lymphocytic depletion with diffuse fibrosis (procedure)
C4031494|biopsy of breast showed liposarcoma dedifferentiated
C4031494|biopsy of breast showed dedifferentiated liposarcoma
C4031494|biopsy of breast showed dedifferentiated liposarcoma (procedure)
C4031489|biopsy of breast showed round cell liposarcoma
C4031489|biopsy of breast showed liposarcoma round cell
C4031489|biopsy of breast showed round cell liposarcoma (procedure)
C4031513|biopsy of breast showed hemangioendothelioma
C4031513|biopsy of breast showed hemangioendothelioma (procedure)
C4031488|biopsy of breast showed well differentiated liposarcoma (procedure)
C4031488|biopsy of breast showed well differentiated liposarcoma
C4031488|biopsy of breast showed liposarcoma well differentiated
C4031479|biopsy of breast showed grade 2 follicular lymphoma
C4031479|biopsy of breast showed grade 2 follicular lymphoma (procedure)
C4031479|biopsy of breast showed lymphoma follicular grade 2
C4031472|biopsy of breast showed mantle cell lymphoma
C4031472|biopsy of breast showed lymphoma mantle cell
C4031472|biopsy of breast showed mantle cell lymphoma (procedure)
C4031465|biopsy of breast showed lymphoma precursor cell lymphoblastic b-cell
C4031465|biopsy of breast showed precursor B-cell lymphoblastic lymphoma (procedure)
C4031465|biopsy of breast showed precursor B-cell lymphoblastic lymphoma
C4031464|biopsy of breast showed lymphoma precursor cell lymphoblastic t-cell
C4031464|biopsy of breast showed precursor T-cell lymphoblastic lymphoma (procedure)
C4031464|biopsy of breast showed precursor T-cell lymphoblastic lymphoma
C4031529|biopsy of breast showed embryonal carcinosarcoma (procedure)
C4031529|biopsy of breast showed carcinosarcoma embryonal
C4031529|biopsy of breast showed embryonal carcinosarcoma
C4031521|biopsy of breast showed fascial fibrosarcoma
C4031521|biopsy of breast showed fascial fibrosarcoma (procedure)
C4031521|biopsy of breast showed fibrosarcoma fascial
C4031506|biopsy of breast showed Hodgkin's lymphoma with lymphocytic depletion
C4031506|biopsy of breast showed Hodgkin's lymphoma with lymphocytic depletion (procedure)
C4031493|biopsy of breast showed fibroblastic liposarcoma (procedure)
C4031493|biopsy of breast showed fibroblastic liposarcoma
C4031493|biopsy of breast showed liposarcoma fibroblastic
C4031483|biopsy of breast showed lymphoma burkitt's
C4031483|biopsy of breast showed Burkitt's lymphoma
C4031483|biopsy of breast showed Burkitt's lymphoma (procedure)
C4031558|biopsy of breast showed medullary carcinoma with lymphoid stroma (procedure)
C4031558|biopsy of breast showed carcinoma medullary with lymphoid stroma
C4031558|biopsy of breast showed medullary carcinoma with lymphoid stroma
C4031502|biopsy of breast showed Hodgkin's lymphoma with grade 2 nodular sclerosis
C4031502|biopsy of breast showed Hodgkin's lymphoma with grade 2 nodular sclerosis (procedure)
C4031502|biopsy of breast showed hodgkin's lymphoma with nodular sclerosis grade 2
C4031474|biopsy of breast showed lymphoplasmacytic lymphoma
C4031474|biopsy of breast showed lymphoma lymphoplasmacytic
C4031474|biopsy of breast showed lymphoplasmacytic lymphoma (procedure)
C4031501|biopsy of breast showed Hodgkin's lymphoma with nodular sclerosis in cellular phase (procedure)
C4031501|biopsy of breast showed Hodgkin's lymphoma with nodular sclerosis in cellular phase
C4031467|biopsy of breast showed non-Hodgkin's lymphoma
C4031467|biopsy of breast showed lymphoma non-hodgkin's
C4031467|biopsy of breast showed non-Hodgkin's lymphoma (procedure)
C4031455|biopsy of breast showed myxoid leiomyosarcoma (procedure)
C4031455|biopsy of breast showed myxoid leiomyosarcoma
C4031455|biopsy of breast showed myosarcoma leiomyosarcoma myxoid
C4031580|biopsy of breast showed comedocarcinoma (procedure)
C4031580|biopsy of breast showed carcinoma comedocarcinoma
C4031580|biopsy of breast showed comedocarcinoma
C4031560|biopsy of breast showed medullary carcinoma (procedure)
C4031560|biopsy of breast showed medullary carcinoma
C4031560|biopsy of breast showed carcinoma medullary
C4031519|biopsy of breast showed infantile fibrosarcoma (procedure)
C4031519|biopsy of breast showed infantile fibrosarcoma
C4031519|biopsy of breast showed fibrosarcoma infantile
C4031511|biopsy of breast showed Hodgkin's lymphoma (procedure)
C4031511|biopsy of breast showed Hodgkin's lymphoma
C4031510|biopsy of breast showed Hodgkin's lymphoma granuloma
C4031510|biopsy of breast showed Hodgkin's lymphoma granuloma (procedure)
C4031463|biopsy of breast showed small b-cell lymphocytic lymphoma
C4031463|biopsy of breast showed small b-cell lymphocytic lymphoma (procedure)
C4031463|biopsy of breast showed lymphoma small b-cell lymphocytic
C4031452|biopsy of breast showed plasmacytoma extramedullary
C4031452|biopsy of breast showed extramedullary plasmacytoma
C4031452|biopsy of breast showed extramedullary plasmacytoma (procedure)
C4031567|biopsy of breast showed infiltrating ductal carcinoma mixed with other types (procedure)
C4031567|biopsy of breast showed carcinoma infiltrating ductal mixed with other types
C4031567|biopsy of breast showed infiltrating ductal carcinoma mixed with other types
C4031518|biopsy of breast showed fibrosarcoma, solitary fibrous tumor (procedure)
C4031518|biopsy of breast showed fibrosarcoma, solitary fibrous tumor
C4031518|biopsy of breast showed fibrosarcoma solitary fibrous tumor
C4031456|biopsy of breast showed epithelioid leiomyosarcoma (procedure)
C4031456|biopsy of breast showed myosarcoma leiomyosarcoma epithelioid
C4031456|biopsy of breast showed epithelioid leiomyosarcoma
C4031453|biopsy of breast showed plasmacytoma (procedure)
C4031453|biopsy of breast showed plasmacytoma
C4031602|biopsy of breast showed adenocarcinoma mucin-producing
C4031602|biopsy of breast showed mucin-producing adenocarcinoma
C4031602|biopsy of breast showed mucin-producing adenocarcinoma (procedure)
C4031527|biopsy of breast showed clear cell type neoplasm (procedure)
C4031527|biopsy of breast showed clear cell type neoplasm
C4031527|biopsy of breast showed clear cell type
C4031481|biopsy of breast showed lymphoma follicular
C4031481|biopsy of breast showed follicular lymphoma
C4031481|biopsy of breast showed follicular lymphoma (procedure)
C4031480|biopsy of breast showed lymphoma follicular grade 1
C4031480|biopsy of breast showed grade 1 follicular lymphoma
C4031480|biopsy of breast showed grade 1 follicular lymphoma (procedure)
C4031473|biopsy of breast showed malt lymphoma
C4031473|biopsy of breast showed lymphoma malt
C4031473|biopsy of breast showed malt lymphoma (procedure)
C4031469|biopsy of breast showed mature t-cell angioimmunoblastic lymphoma (procedure)
C4031469|biopsy of breast showed mature t-cell angioimmunoblastic lymphoma
C4031469|biopsy of breast showed lymphoma mature t-cell angioimmunoblastic
C4031460|biopsy of breast showed mesenchymoma
C4031460|biopsy of breast showed mesenchymoma (procedure)
C4031600|biopsy of breast showed polymorphous adenocarcinoma, low grade
C4031600|biopsy of breast showed polymorphous adenocarcinoma, low grade (procedure)
C4031600|biopsy of breast showed adenocarcinoma polymorphous, low grade
C4031522|biopsy of breast showed adenofibrosarcoma
C4031522|biopsy of breast showed adenofibrosarcoma (procedure)
C4031522|biopsy of breast showed fibrosarcoma adenofibrosarcoma
C4031492|biopsy of breast showed mixed type liposarcoma (procedure)
C4031492|biopsy of breast showed mixed type liposarcoma
C4031492|biopsy of breast showed liposarcoma mixed type
C4031478|biopsy of breast showed grade 3 follicular lymphoma (procedure)
C4031478|biopsy of breast showed grade 3 follicular lymphoma
C4031478|biopsy of breast showed lymphoma follicular grade 3
C4031487|biopsy of breast showed lymphoma
C4031487|biopsy of breast showed lymphoma (procedure)
C4031462|biopsy of breast showed malignant neoplasm (procedure)
C4031462|biopsy of breast showed malignant neoplasm
C4031423|biopsy of breast showed small cell type neoplasm (procedure)
C4031423|biopsy of breast showed small cell type
C4031423|biopsy of breast showed small cell type neoplasm
C4031421|biopsy of breast showed spindle cell type neoplasm
C4031421|biopsy of breast showed spindle cell type
C4031421|biopsy of breast showed spindle cell type neoplasm (procedure)
C4031561|biopsy of breast showed lobular carcinoma mixed with other types of carcinoma (procedure)
C4031561|biopsy of breast showed carcinoma lobular mixed with other types of carcinom
C4031561|biopsy of breast showed lobular carcinoma mixed with other types of carcinoma
C4031528|biopsy of breast showed myoepithelioma carcinosarcoma
C4031528|biopsy of breast showed myoepithelioma carcinosarcoma (procedure)
C4031528|biopsy of breast showed carcinosarcoma myoepithelioma
C4031520|biopsy of breast showed fibromyxosarcoma
C4031520|biopsy of breast showed fibrosarcoma fibromyxosarcoma
C4031520|biopsy of breast showed fibromyxosarcoma (procedure)
C4031509|biopsy of breast showed hodgkin's lymphoma lymphocyte-rich
C4031509|biopsy of breast showed Hodgkin's lymphocyte-rich lymphoma (procedure)
C4031509|biopsy of breast showed Hodgkin's lymphocyte-rich lymphoma
C4031504|biopsy of breast showed Hodgkin's lymphoma with nodular sclerosis
C4031504|biopsy of breast showed Hodgkin's lymphoma with nodular sclerosis (procedure)
C4031471|biopsy of breast showed lymphoma marginal zone b-cell
C4031471|biopsy of breast showed marginal zone b-cell lymphoma
C4031471|biopsy of breast showed marginal zone b-cell lymphoma (procedure)
C4031470|biopsy of breast showed mature t-cell lymphoma
C4031470|biopsy of breast showed lymphoma mature t-cell
C4031470|biopsy of breast showed mature t-cell lymphoma (procedure)
C4031459|biopsy of breast showed myosarcoma (procedure)
C4031459|biopsy of breast showed myosarcoma
C4031546|biopsy of breast showed secretory carcinoma
C4031546|biopsy of breast showed carcinoma secretory
C4031546|biopsy of breast showed secretory carcinoma (procedure)
C4031507|biopsy of breast showed Hodgkin's lymphoma sarcoma
C4031507|biopsy of breast showed Hodgkin sarcoma
C4031507|biopsy of breast showed Hodgkin sarcoma (procedure)
C4031475|biopsy of breast showed diffuse large b-cell immunoblastic lymphoma
C4031475|biopsy of breast showed diffuse large b-cell immunoblastic lymphoma (procedure)
C4031475|biopsy of breast showed lymphoma large b-cell, diffuse immunoblastic
C4031461|biopsy of breast showed mastocytosis
C4031461|biopsy of breast showed mastocytosis (procedure)
C4031429|biopsy of breast showed sarcoma neurosarcoma
C4031429|biopsy of breast showed neurosarcoma
C4031429|biopsy of breast showed neurosarcoma (procedure)
C4031586|biopsy of breast showed acinar cell carcinoma (procedure)
C4031586|biopsy of breast showed acinar cell carcinoma
C4031586|biopsy of breast showed carcinoma acinar cell
C4031496|biopsy of breast showed large cell neuroendocrine carcinoma
C4031496|biopsy of breast showed carcinoma large cell neuroendocrine
C4031496|biopsy of breast showed large cell neuroendocrine carcinoma (procedure)
C4031530|biopsy of breast showed carcinosarcoma
C4031530|biopsy of breast showed carcinosarcoma (procedure)
C4031495|biopsy of breast showed liposarcoma (procedure)
C4031495|biopsy of breast showed liposarcoma
C4031477|biopsy of breast showed histiocytosis lymphoma
C4031477|biopsy of breast showed histiocytosis lymphoma (procedure)
C4031477|biopsy of breast showed lymphoma histiocytosis
C4031476|biopsy of breast showed diffuse large b-cell lymphoma (procedure)
C4031476|biopsy of breast showed diffuse large b-cell lymphoma
C4031476|biopsy of breast showed lymphoma large b-cell, diffuse
C4031457|biopsy of breast showed myosarcoma leiomyosarcoma
C4031457|biopsy of breast showed leiomyosarcoma (procedure)
C4031457|biopsy of breast showed leiomyosarcoma
C4031585|biopsy of breast showed acinar cell cystadenocarcinoma
C4031585|biopsy of breast showed acinar cell cystadenocarcinoma (procedure)
C4031585|biopsy of breast showed carcinoma acinar cell cystadenocarcinoma
C4031515|biopsy of breast showed giant cell type neoplasm (procedure)
C4031515|biopsy of breast showed giant cell type neoplasm
C4031515|biopsy of breast showed giant cell type
C4031508|biopsy of breast showed Hodgkin's mixed cellularity lymphoma
C4031508|biopsy of breast showed hodgkin's lymphoma mixed cellularity
C4031508|biopsy of breast showed Hodgkin's mixed cellularity lymphoma (procedure)
C4031491|biopsy of breast showed myxoid liposarcoma (procedure)
C4031491|biopsy of breast showed myxoid liposarcoma
C4031491|biopsy of breast showed liposarcoma myxoid
C4031458|biopsy of breast showed angiomyosarcoma
C4031458|biopsy of breast showed myosarcoma angiomyosarcoma
C4031458|biopsy of breast showed angiomyosarcoma (procedure)
C0346787|Malignant melanoma of breast
C0346787|Malignant melanoma of breast (disorder)
C0346787|breast; melanoma
C0346787|melanoma; breast
C0346787|Malignant Breast Melanoma
C0346787|Malignant Melanoma of the Breast
C0346787|Breast Melanoma
C0346986|metastasis of malignant neoplasm to skin of breast (diagnosis)
C0346986|metastasis of malignant neoplasm to skin of breast
C0346986|Secondary malignant neoplasm of skin of breast (disorder)
C0346986|Secondary malignant neoplasm of skin of breast
C0346986|skin neoplasm malignant breast secondary
C0346986|secondary malignant skin neoplasm of breast (diagnosis)
C0346986|secondary malignant skin neoplasm of breast
C0346986|Metastatic malignant neoplasm to skin of breast
C1282471|Local recurrence of malignant tumor of breast (disorder)
C1282471|Local recurrence of malignant tumor of breast
C1282471|Local recurrence of malignant tumour of breast
C1134719|Carcinomas, Infiltrating Duct
C1134719|Invasive Ductal Breast Carcinoma
C1134719|infiltrating ductal carcinoma of breast
C1134719|infiltrating ductal carcinoma of breast (diagnosis)
C1134719|Carcinoma, Ductal, Breast
C1134719|Carcinoma, Invasive Ductal, Breast
C1134719|Invasive Ductal Carcinoma, Breast
C1134719|Carcinoma, Ductal, Breast [Disease/Finding]
C1134719|Carcinoma, Infiltrating Duct
C1134719|infiltrating ductal carcinoma
C1134719|Invasive Ductal Carcinoma, Not Otherwise Specified
C1134719|BREAST CANCER, INVASIVE DUCTAL
C1134719|Breast ductal cancer infiltrating
C1134719|Invasive ductal breast cancer
C1134719|Breast ductal cancer invasive
C1134719|Infiltrating ductal breast cancer
C1134719|Infiltrating ductular carcinoma
C1134719|Infiltrating ductular carcinoma (morphologic abnormality)
C1134719|Infiltrating duct carcinoma of breast (disorder)
C1134719|Infiltrating duct carcinoma of breast
C1134719|Invasive duct carcinoma of breast
C1134719|Invasive ductal carcinoma of breast
C1134719|ductal invasive breast carcinoma
C1134719|carcinoma; ductal, infiltrating, unspecified site
C1134719|carcinoma; ductular, infiltrating, unspecified site
C1134719|carcinoma; infiltrating duct, unspecified site
C1134719|carcinoma; infiltrating ductular, unspecified site
C1134719|ductal; carcinoma, infiltrating, unspecified site
C1134719|ductular; carcinoma, infiltrating, unspecified site
C1134719|infiltrating; ductal adenocarcinoma, unspecified site
C1134719|infiltrating; ductal carcinoma, unspecified site
C1134719|infiltrating; ductular carcinoma, unspecified site
C1134719|Infiltrating Ductal Adenocarcinoma
C1134719|Infiltrating Ductal Breast Carcinoma
C1134719|Infiltrating Ductal Carcinoma of the Breast
C1134719|Invasive Ductal Adenocarcinoma
C1134719|Invasive Ductal Carcinoma of the Breast
C1134719|Invasive Ductal Carcinoma, NOS
C1134719|Invasive Ductal Carcinoma, NST
C1134719|Invasive Ductal Carcinoma
C1134719|Invasive Ductal Carcinoma, No Specific Type
C1386255|ductal; infiltrating adenocarcinoma, unspecified site, female
C1386255|adenocarcinoma; ductal infiltrating, unspecified site, female
C1386267|adenocarcinoma; infiltrating duct, unspecified site
C1386268|adenocarcinoma; infiltrating duct, unspecified site, female
C1386269|inflammatory; adenocarcinoma, unspecified site
C1386269|adenocarcinoma; inflammatory, unspecified site
C1386276|adenocarcinoma; intraductal, noninfiltrating, papillary, with invasion, unspecified site
C1386278|adenocarcinoma; intraductal, papillary, with invasion, unspecified site
C1386278|adenocarcinoma; papillary, intraductal, with invasion, unspecified site
C1386278|papillary; adenocarcinoma, intraductal, with invasion, unspecified site
C1386282|lobular; adenocarcinoma, unspecified site
C1386282|adenocarcinoma; lobular, unspecified site
C1391891|breast; carcinoma in situ, lobular with infiltrating duct
C1391891|carcinoma in situ; lobular with infiltrating duct, breast
C1391891|lobular; carcinoma in situ, with infiltrating duct, breast
C1391892|carcinoma in situ; lobular with infiltrating duct, unspecified site
C1391892|lobular; carcinoma in situ, with infiltrating duct, unspecified site
C1391902|carcinoma; ductal with lobular (infiltrating), unspecified site
C1391902|ductal; carcinoma with lobular (infiltrating), unspecified site
C1391903|carcinoma; ductal, infiltrating, with lobular carcinoma in situ, unspecified site
C1391903|ductal; carcinoma, infiltrating, with lobular carcinoma in situ, unspecified site
C1391904|carcinoma; ductal, infiltrating, with lobular carcinoma, unspecified site
C1391904|ductal; carcinoma, infiltrating, with lobular carcinoma, unspecified site
C1391904|infiltrating; ductal carcinoma, with lobular carcinoma, unspecified site
C0334384|Carcinoma of breast with ductal and lobular features (disorder)
C0334384|Carcinoma of breast with ductal and lobular features
C0334384|Mixed ductal and lobular carcinoma of breast
C0334384|Infiltrating duct and lobular carcinoma
C0334384|Infiltrating duct and lobular carcinoma (disorder)
C0334384|breast neoplasm malignant carcinoma with ductal and lobular features
C0334384|Carcinoma of breast with ductal and lobular features (diagnosis)
C0334384|[M] Infiltrating duct and lobular carcinoma
C0334384|[M]Infiltrating duct and lobular carcinoma
C0334384|Mixed ductal lobular breast carcinoma
C0334384|Infiltrating duct and lobular carcinoma in situ
C0334384|Intraductal and lobular carcinoma
C0334384|Lobular and ductal carcinoma
C0334384|Infiltrating duct and lobular carcinoma (morphologic abnormality)
C0334384|Infiltrating lobular carcinoma and ductal carcinoma in situ
C0334384|carcinoma; infiltrating duct with lobular ca, unspecified site
C0334384|DCIS and ILC
C0334384|DCIS and Infiltrating Lobular Carcinoma
C0334384|Ductal Carcinoma in situ and Infiltrating Lobular Carcinoma
C0334384|Ductal and Lobular Carcinoma
C0334384|Infiltrating Ductal and Lobular Carcinoma in situ
C0334384|LCIS and Infiltrating Ductal Carcinoma
C0334384|Lobular Carcinoma in situ and Infiltrating Ductal Carcinoma
C0334384|Lobular Carcinoma in situ and Invasive Ductal Carcinoma
C0334384|Mixed Ductal and Lobular Breast Carcinoma
C0334384|Mixed Ductal and Lobular Carcinoma of the Breast
C0334384|Mixed Lobular and Ductal Breast Carcinoma
C0334384|Mixed Lobular and Ductal Carcinoma of Breast
C0334384|Mixed Lobular and Ductal Carcinoma of the Breast
C0334384|Mixed Lobular and Ductal Carcinoma
C0334384|Non-Infiltrating Ductal Carcinoma and ILC
C0334384|Non-Infiltrating Ductal Carcinoma and Infiltrating Lobular Carcinoma
C0334384|Ductal Breast Carcinoma In Situ and Invasive Lobular Carcinoma
C0334384|Invasive Ductal and Lobular Carcinoma In Situ
C0334385|Inflammatory adenocarcinoma
C0334385|Inflammatory carcinoma
C0334385|Inflammatory carcinoma (morphologic abnormality)
C0334385|carcinoma; inflammatory, unspecified site
C0334385|inflammatory; carcinoma, unspecified site
C1391916|carcinoma; intraductal, papillary with invasion, unspecified site
C1391916|intraductal; carcinoma, papillary with invasion, unspecified site
C0334318|Lipid-rich carcinoma (disorder)
C0334318|Lipid-rich carcinoma
C0334318|[M] Lipid-rich carcinoma
C0334318|[M]Lipid-rich carcinoma
C0334318|Lipid-rich carcinoma (morphologic abnormality)
C0334318|carcinoma; lipid-rich
C0334318|lipid-rich; carcinoma
C1391922|carcinoma; lobular with intraductal, unspecified site
C1391923|carcinoma; lobular, unspecified site
C1391923|lobular; carcinoma, unspecified site
C0334380|Medullary carcinoma with lymphoid stroma
C0334380|Medullary carcinoma with lymphoid stroma (morphologic abnormality)
C0334380|carcinoma; medullary with lymphoid stroma, unspecified site
C0334380|medullary; carcinoma with lymphoid stroma, unspecified site
C1391934|carcinoma; papillary, intraductal (noninfiltrating), with invasion, unspecified site
C1391934|papillary; carcinoma, intraductal (noninfiltrating), with invasion, unspecified site
C1403125|lobular; carcinoma, with intraductal carcinoma, unspecified site
C0279855|cellular diagnosis, breast cancer
C0279855|breast cancer cellular diagnosis
C0281663|breast cancer and pregnancy
C0281663|pregnancy and breast cancer
C0238033|Cancer, Male Breast
C0238033|Carcinoma of Male Breast
C0238033|Breast Cancer, Male
C0238033|Male Breast Cancer
C0238033|Ca breast - male (disorder)
C0238033|Ca breast - male
C0238033|Carcinoma of male breast (diagnosis)
C0238033|breast neoplasm malignant male carcinoma
C0238033|Breast cancer male NOS
C0238033|Cancer of male breast
C0238033|Breast cancer male
C0238033|Breast Carcinoma, Male
C0238033|Carcinoma of male breast (disorder)
C0238033|Male Breast Carcinoma
C0238033|Carcinoma, Male Breast
C0238033|Carcinoma of the Male Breast
C0238033|Carcinoma;breast;M
C0238033|carcinoma of the breast
C0346993|Metastatic Neoplasm to the Breast
C0346993|secondary malignant neoplasm of breast (diagnosis)
C0346993|secondary malignant neoplasm of breast
C0346993|Metastases to breast
C0346993|Second malig neo breast
C0346993|Secondary malignant neoplasm of female breast (diagnosis)
C0346993|Secondary malignant neoplasm of female breast
C0346993|breast neoplasm malignant female secondary
C0346993|Metastatic Malignant Neoplasm to the Breast
C0346993|Metastatic Malignant Neoplasm in the Breast
C0346993|Breast metastases
C0346993|Metastasis to breast
C0346993|Secondary malignant deposit to breast
C0346993|Metastatic malignant neoplasm to female breast
C0346993|Secondary malignant neoplasm of female breast (disorder)
C0346993|Metastatic malignant neoplasm to female breast, NOS
C0346993|Secondary malignant neoplasm of female breast, NOS
C0346993|Metastatic Cancer to the Breast
C0346993|Metastatic Tumor to the Breast
C0346993|Breast Metastasis
C1334565|Malignant Breast Eccrine Spiradenoma
C1334565|Malignant Eccrine Spiradenoma of Breast
C1334565|Malignant Eccrine Spiradenoma of the Breast
C1334564|Malignant Adenomyoepithelioma of Breast
C1334564|Malignant Adenomyoepithelioma of the Breast
C1334564|Malignant Breast Adenomyoepithelioma
C1334564|Breast Adenomyoepithelioma with Malignant Change
C1704251|Primary Breast Lymphoma
C1704251|Breast Lymphoma
C1704251|Lymphoma of Breast
C1704251|Lymphoma of the Breast
C0859086|Malignant nipple neoplasm NOS
C0859086|Malignant nipple neoplasm
C0859086|Malignant Neoplasm of Nipple
C0859086|Malignant Neoplasm of the Nipple
C0859086|Malignant Nipple Tumor
C0859086|Malignant Tumor of Nipple
C0859086|Malignant Tumor of the Nipple
C2211713|mast cell sarcoma of breast (diagnosis)
C2211713|mast cell sarcoma of breast
C0345867|Carcinoma in situ of descending colon
C0345867|Carcinoma in situ of descending colon (disorder)
C0700315|large intestine adenocarcinoma - splenic flexure carcinoma
C0700315|Carcinoma of splenic flexure
C0700315|Carcinoma of splenic flexure (diagnosis)
C0700315|Carcinoma of splenic flexure (disorder)
C0728951|carcinoma of appendix
C0728951|carcinoma of appendix (diagnosis)
C0728951|Appendix Cancer
C0728951|(Ca appendix) or (appendix carcinoma)
C0728951|Appendix carcinoma
C0728951|Ca appendix
C0728951|(Ca appendix) or (appendix carcinoma) (disorder)
C0728951|Carcinoma of the appendix
C0856355|Cancer of sigmoid colon (excluding rectosigmoid)
C0856355|Cancer of sigmoid colon (excl rectosigmoid)
C0153439|Malignant neoplasm of ascending colon
C0153439|Ascending colon
C0153439|malignant neoplasm of ascending colon (diagnosis)
C0153439|cancer of ascending colon
C0153439|malignant tumor of ascending colon
C0153439|Malig neo ascend colon
C0153439|Ca ascending colon (disorder)
C0153439|Ca ascending colon
C0153439|Ascending colon cancer
C0153439|Malignant tumour of ascending colon
C0153439|Malignant tumor of ascending colon (disorder)
C0153439|Malignant neoplasm of right colon
C0496779|Appendix
C0496779|Malignant neoplasm of appendix
C0496779|malignant neoplasm of appendix (diagnosis)
C0496779|malignant appendiceal neoplasm
C0496779|malignant tumor of appendix
C0496779|Malignant neo appendix
C0496779|Appendix cancer
C0496779|Malignant neoplasm of appendix vermiformis
C0496779|Cancer, Appendiceal
C0496779|Cancer of the Appendix
C0496779|Cancer of Appendix
C0496779|Cancer, Appendix
C0496779|Malignant tumour of appendix
C0496779|Malignant tumor of appendix (disorder)
C0496779|Malignant Appendix Neoplasm
C0496779|Malignant Appendix Tumor
C0496779|Malignant Neoplasm of the Appendix
C0496779|Malignant Tumor of the Appendix
C0496779|Appendiceal Cancer
C0349051|Malignant neoplasm overlapping colon site
C0349051|Overlapping lesion of colon
C0349051|Malignant neoplasm of overlapping sites of colon
C0349051|malignant neoplasm, overlapping lesion of colon (diagnosis)
C0349051|malignant neoplasm, overlapping lesion of colon
C0349051|large intestine neoplasm malignant, overlapping lesion of colon
C0349051|Malignant neoplasm, overlapping lesion of colon (disorder)
C0153433|Malignant neoplasm of hepatic flexure
C0153433|Hepatic flexure
C0153433|Malignant neoplasm of hepatic flexure of colon
C0153433|malignant neoplasm of hepatic flexure (diagnosis)
C0153433|malignant tumor of hepatic flexure
C0153433|Mal neo hepatic flexure
C0153433|Ca hepatic flexure - colon (disorder)
C0153433|Ca hepatic flexure - colon
C0153433|Hepatic flexure colon cancer
C0153433|Malignant tumour of hepatic flexure
C0153433|Malignant tumor of hepatic flexure (disorder)
C0153434|Malignant neoplasm of transverse colon
C0153434|Transverse colon
C0153434|malignant neoplasm of transverse colon (diagnosis)
C0153434|malignant tumor of transverse colon
C0153434|Mal neo transverse colon
C0153434|Ca transverse colon
C0153434|Ca transverse colon (disorder)
C0153434|Cancer of transverse colon
C0153434|Transverse colon cancer
C0153434|Malignant tumour of transverse colon
C0153434|Malignant tumor of transverse colon (disorder)
C0153435|Malignant neoplasm of descending colon
C0153435|Descending colon
C0153435|malignant neoplasm of descending colon (diagnosis)
C0153435|malignant tumor of descending colon
C0153435|Mal neo descend colon
C0153435|Ca descending colon
C0153435|Ca descending colon (disorder)
C0153435|Cancer of descending colon
C0153435|Descending colon cancer
C0153435|Malignant tumour of descending colon
C0153435|Malignant tumor of descending colon (disorder)
C0153435|Malignant neoplasm of left colon
C0153436|Malignant neoplasm of sigmoid colon
C0153436|Sigmoid colon
C0153436|malignant neoplasm of sigmoid colon (diagnosis)
C0153436|malignant tumor of sigmoid colon
C0153436|Mal neo sigmoid colon
C0153436|Ca sigmoid colon
C0153436|Ca sigmoid colon (disorder)
C0153436|Sigmoid colon cancer
C0153436|Malignant tumour of sigmoid colon
C0153436|Malignant tumor of sigmoid colon (disorder)
C0153443|Malignant neoplasm of rectosigmoid junction
C0153443|Mal neo rectosigmoid jct
C0153443|Malignant neoplasm of rectosigmoid (colon)
C0153443|rectal neoplasm malignant rectosigmoid junction
C0153443|malignant neoplasm of rectosigmoid junction (diagnosis)
C0153443|Rectosigmoid colon cancer
C0153443|Ca rectosigmoid junction
C0153443|Malignant tumor of rectosigmoid junction
C0153443|Malignant tumour of rectosigmoid junction
C0153443|Malignant tumor of rectosigmoid junction (disorder)
C0153443|Malignant Neoplasm of the Rectosigmoid Junction
C0153443|Malignant Rectosigmoid Neoplasm
C0153443|Malignant Rectosigmoid Tumor
C0153443|Malignant Tumor of the Rectosigmoid Junction
C0153443|Malignant neoplasm of rectosigmoid colon
C0153443|Malignant neoplasm of rectosigmoid
C1096639|mucinous cystadenocarcinoma of appendix (diagnosis)
C1096639|mucinous cystadenocarcinoma of appendix
C1096639|Mucinous cystadenocarcinoma appendix
C1096639|Colloid Cystadenocarcinoma of Appendix
C1096639|Colloid Cystadenocarcinoma of the Appendix
C1096639|Colloidal Cystadenocarcinoma of Appendix
C1096639|Colloidal Cystadenocarcinoma of the Appendix
C1096639|Mucinous Cystadenocarcinoma of the Appendix
C1096639|Appendiceal Colloid Cystadenocarcinoma
C1096639|Appendiceal Colloidal Cystadenocarcinoma
C1096639|Appendiceal Mucinous Cystadenocarcinoma
C1096639|Appendix Colloid Cystadenocarcinoma
C1096639|Appendix Colloidal Cystadenocarcinoma
C1096639|Appendix Mucinous Cystadenocarcinoma
C0153440|Malignant neoplasm of splenic flexure
C0153440|Splenic flexure
C0153440|Malignant neoplasm of splenic flexure of colon
C0153440|malignant neoplasm of splenic flexure (diagnosis)
C0153440|malignant tumor of splenic flexure
C0153440|Mal neo splenic flexure
C0153440|Ca splenic flexure - colon (disorder)
C0153440|Ca splenic flexure - colon
C0153440|Cancer of splenic flexure
C0153440|Splenic flexure colon cancer
C0153440|Malignant tumour of splenic flexure
C0153440|Malignant tumor of splenic flexure (disorder)
C0153437|Cecum
C0153437|Malignant neoplasm of cecum
C0153437|Caecum
C0153437|Malignant neoplasm of caecum
C0153437|malignant neoplasm of cecum (diagnosis)
C0153437|malignant tumor of cecum
C0153437|Malignant neoplasm cecum
C0153437|Ca caecum
C0153437|Ca cecum
C0153437|Cecum--Cancer
C0153437|Cecal cancer
C0153437|Caecal cancer
C0153437|Cancer of the Cecum
C0153437|Cancer, Cecal
C0153437|CA - Cancer of caecum
C0153437|CA - Cancer of cecum
C0153437|Cancer of caecum
C0153437|Cancer of cecum
C0153437|Malignant tumour of caecum
C0153437|Malignant tumor of cecum (disorder)
C0153437|Malignant Cecum Neoplasm
C0153437|Malignant Cecum Tumor
C0153437|Malignant Neoplasm of the Cecum
C0153437|Malignant Tumor of the Cecum
C0007102|Malignant neoplasm of colon
C0007102|colon cancer
C0007102|Cancer of colon
C0007102|Malignant neoplasm of colon, unspecified
C0007102|Malignant tumor of colon
C0007102|Colon, unspecified
C0007102|Cancers, Colon
C0007102|Colon Cancers
C0007102|Cancer, Colonic
C0007102|Cancers, Colonic
C0007102|Colonic Cancers
C0007102|Malignant neo colon NOS
C0007102|Cancer, Colon
C0007102|Malignant neoplasm of colon, unspecified site
C0007102|Colonic cancer
C0007102|Ca colon NOS (disorder)
C0007102|Malignant neoplasm of colon NOS
C0007102|Ca colon NOS
C0007102|Malignant neoplasm of colon (& NOS) (disorder)
C0007102|Malignant neoplasm of colon (& NOS)
C0007102|Malignant neoplasm of colon NOS (disorder)
C0007102|-- Colon Cancer
C0007102|Colon cancer NOS
C0007102|Colonic cancer NOS
C0007102|Cancer of the Colon
C0007102|CA - Cancer of colon
C0007102|Malignant tumour of colon
C0007102|Malignant tumor of colon (disorder)
C0007102|Malignant neoplasm of colon, NOS
C0007102|Colon Neoplasm, Malignant
C0007102|Colon Tumor, Malignant
C0007102|Malignant Colon Neoplasm
C0007102|Malignant Colon Tumor
C0007102|Malignant Colonic Neoplasm
C0007102|Malignant Colonic Tumor
C0007102|Malignant Neoplasm of the Colon
C0007102|Malignant Tumor of the Colon
C1333990|HNPCC
C1333990|hereditary non-polyposis colon cancer
C1333990|hereditary non-polyposis colon cancer (diagnosis)
C1333990|Hereditary Nonpolyposis Colorectal Cancer
C1333990|Lynch Syndrome
C1333990|HNPCC - hereditary nonpolyposis colorectal cancer
C1333990|Hereditary nonpolyposis colon cancer
C1333990|Hereditary Nonpolyposis Colon Cancer (hMSH2, hMLH1, hPMS1, hPMS2)
C1333990|Colon Cancer, Familial Nonpolyposis
C1333990|Colorectal Cancer Hereditary Nonpolyposis
C1333990|Lynch Syndrome I
C1333990|Lynch Cancer Family Syndrome I
C1333990|HNPCC - hereditary nonpolyposis colon cancer
C1333990|Hereditary nonpolyposis colon cancer (disorder)
C1333990|hereditary non-polyposis colon cancer (hMSH2, hMLH1, hPMS1, hPMS2)
C1333990|Familial Non-Polyposis Colon Cancer (hMSH2, hMLH1, hPMS1, hPMS2)
C1333990|Hereditary Colorectal Endometrial Cancer Syndrome
C1333990|Hereditary Defective Mismatch Repair Syndrome
C1333990|Syndrome, Lynch
C3472669|Primary adenocarcinoma of colon
C3472669|Primary adenocarcinoma of colon (disorder)
C0346630|Malignant neoplasm of other specified sites of colon (disorder)
C0346630|Malignant neoplasm of other specified sites of colon
C1304819|Primary malignant neoplasm of colon
C1304819|large intestine neoplasm malignant, colon primary
C1304819|Primary malignant neoplasm of colon (diagnosis)
C1304819|Primary malignant neoplasm of colon (disorder)
C0519037|Primary Colon Lymphoma
C0519037|Colonic lymphoma
C0519037|Lymphoma of colon (disorder)
C0519037|Lymphoma of colon
C0519037|Colon Lymphoma
C0519037|Lymphoma of the Colon
C0346974|Metastatic Neoplasm to the Colon
C0346974|Secondary malignant neoplasm of colon
C0346974|Secondary malignant neoplasm of colon (disorder)
C0346974|secondary malignant neoplasm of colon (diagnosis)
C0346974|Metastatic Malignant Neoplasm in the Colon
C0346974|Metastatic Malignant Neoplasm to the Colon
C0346974|Metastatic malignant neoplasm to colon
C0346974|Metastatic malignant neoplasm to colon, NOS
C0346974|Secondary malignant neoplasm of colon, NOS
C0346974|Metastatic Tumor to the Colon
C1282478|local recurrence of malignant neoplasm of colon (diagnosis)
C1282478|local recurrence of malignant neoplasm of colon
C1282478|Local recurrence of malignant tumor of colon (disorder)
C1282478|Local recurrence of malignant tumor of colon
C1282478|Local recurrence of malignant tumour of colon
C1386266|adenocarcinoma; in polyposis coli
C1391915|carcinoma; in polyposis coli
C1391915|polyposis coli; with carcinoma
C1391940|carcinoma; poliposis coli
C1391940|poliposis coli; carcinoma
C0334293|Adenocarcinoma in adenomatous polyposis coli
C0334293|Adenocarcinoma in adenomatous polyposis coli (morphologic abnormality)
C0334293|polyposis coli; adenocarcinoma, adenomatous (in)
C0279880|cellular diagnosis, colon cancer
C0279880|colon cancer cellular diagnosis
C0280252|stage, colon cancer
C0280252|colon cancer stage
C0699790|CARCINOMA OF COLON
C0699790|Colon carcinoma
C0699790|Colon cancer
C0699790|Carcinoma;colon
C0699790|Carcinoma of colon (disorder)
C0699790|Carcinoma colon
C0699790|Colonic Carcinoma
C0699790|Carcinoma of the Colon
C1333098|Colon Sarcoma
C1333098|Colonic Sarcoma
C1333098|Sarcoma of Colon
C1333098|Sarcoma of the Colon
C0153441|Malignant neoplasm of other specified sites of large intestine
C0153441|Malignant neo colon NEC
C1319315|adenocarcinoma of large intestine (diagnosis)
C1319315|adenocarcinoma of large intestine
C1319315|Colorectal adenocarcinoma
C1319315|large intestine adenocarcinoma
C1319315|Adenocarcinoma of large intestine (disorder)
C1319315|Adenocarcinoma of Large Bowel
C1319315|Adenocarcinoma of the Large Bowel
C1319315|Adenocarcinoma of the Large Intestine
C1319315|Large Bowel Adenocarcinoma
C0809966|Other non-epithelial cancer of skin
C0151779|Malignant melanoma of skin
C0151779|Malignant melanoma of skin, unspecified
C0151779|Melanoma of skin, site unspecified
C0151779|Cutaneous Melanoma
C0151779|CMM
C0151779|malignant melanoma of skin (diagnosis)
C0151779|Malig melanoma skin NOS
C0151779|Melanomas of skin
C0151779|Melanoma (malignant) NOS
C0151779|Skin melanoma
C0151779|Melanoma, Cutaneous Malignant
C0151779|Dysplastic Nevus Syndrome, Hereditary
C0151779|Melanoma, Familial
C0151779|Fammm
C0151779|Familial Atypical Mole-Malignant Melanoma Syndrome
C0151779|[X]Malignant melanoma of skin, unspecified
C0151779|Melanoma of skin
C0151779|[X]Malignant melanoma of skin, unspecified (disorder)
C0151779|Malignant melanoma of skin NOS (disorder)
C0151779|Malignant melanoma of skin NOS
C0151779|Melanoma of skin (disorder)
C0151779|Cutaneous malignant melanoma
C0151779|MELANOMA, MALIGNANT
C0151779|Malignant melanoma of skin stage unspecified
C0151779|Melanoma skin
C0151779|Melanoma of skin (malignant)
C0151779|MM - Malignant melanoma of skin
C0151779|Malignant melanoma of skin (disorder)
C0151779|melanoma, cutaneous
C0151779|Skin cancer, melanoma
C0151779|melanoma; skin
C0151779|skin; melanoma
C0151779|Malignant melanoma of skin, NOS
C0151779|Malignant Cutaneous Melanoma
C0151779|Malignant Melanoma (of Skin), Stage Unspecified
C0151779|Melanoma of the Skin
C0151779|Skin, Melanoma
C0852524|Skin melanomas (excl ocular)
C0852524|Skin melanomas (excluding ocular)
C0852525|Skin neoplasms malignant and unspecified (excl melanoma)
C0852525|Skin neoplasms malignant and unspecified (excluding melanoma)
C0007114|Malignant neoplasm of skin, unspecified
C0007114|Skin cancers
C0007114|Malignant neoplasm of skin
C0007114|skin cancer (diagnosis)
C0007114|skin cancer
C0007114|malignant neoplasm of skin (diagnosis)
C0007114|malignant skin neoplasm
C0007114|Cancer of skin
C0007114|Skin neoplasms malignant and unspecified
C0007114|Cancers, Skin
C0007114|malignant tumor of skin
C0007114|Cancer, Skin
C0007114|Malignant neoplasm of skin NOS
C0007114|Skin Neoplasm, Malignant
C0007114|Malignant tumour of skin (disorder)
C0007114|Malignant neoplasm of skin NOS (disorder)
C0007114|CA - Skin cancer
C0007114|Malignant tumour of skin
C0007114|[X]Malignant neoplasm of skin, unspecified
C0007114|[X]Malignant neoplasm of skin, unspecified (disorder)
C0007114|Skin--Cancer
C0007114|Skin cancer, NOS
C0007114|-- Skin Cancer
C0007114|Skin malignant neoplasm NOS
C0007114|Skin neoplasm malignant
C0007114|Malignant skin neoplasm NOS
C0007114|Skin neoplasm malignant NOS
C0007114|Cancer of the Skin
C0007114|Malignant neoplasm of skin (disorder)
C0007114|Skin cancer, nonmelanomatous (squamous and basal cell)
C0007114|Malignant neoplasm of skin, NOS
C0007114|Malignant Neoplasm of the Skin
C0007114|Malignant Skin Tumor
C0007114|Malignant Tumor of the Skin
C0007114|Melanoma and Non-Melanoma Skin Cancer
C0007114|Skin Cancer, Including Melanoma
C0007114|Neoplasm malig;skin
C0007114|malignant neosplasm of the skin
C2146257|trichilemmocarcinoma of skin (diagnosis)
C2146257|trichilemmocarcinoma of skin
C0699893|CARCINOMA OF SKIN
C0699893|Skin carcinoma
C0699893|carcinoma of skin (diagnosis)
C0699893|Carcinoma;skin
C0699893|nonmelanoma skin cancer
C0699893|Carcinoma skin
C0699893|Skin carcinoma NOS
C0699893|carcinoma of the skin
C0699893|Non-Melanoma Cancer of Skin
C0699893|Non-Melanoma Cancer of the Skin
C0699893|Non-Melanoma Skin Cancer
C0699893|Skin Cancer, Non-Melanoma
C2211421|adenocarcinoma of skin (diagnosis)
C2211421|adenocarcinoma of skin
C2163816|cystadenocarcinoma of skin
C2163816|cystadenocarcinoma of skin (diagnosis)
C0334447|Melanoma Arising from Blue Nevus
C0334447|Blue Nevus-Like Melanoma
C0334447|malignant blue nevus of skin (diagnosis)
C0334447|malignant blue nevus of skin
C0334447|Malignant blue naevus
C0334447|[M]Blue naevus, malignant
C0334447|[M]Blue nevus, malignant
C0334447|Malignant melanoma in blue nevus
C0334447|Malignant melanoma in blue naevus
C0334447|Blue naevus-like melanoma
C0334447|Malignant blue nevus
C0334447|Blue nevus, malignant
C0334447|Blue naevus, malignant
C0334447|Malignant blue naevus of skin
C0334447|Blue nevus, malignant (morphologic abnormality)
C0334447|Malignant blue nevus of skin (disorder)
C0334447|Malignant Blue Nevus of the Skin
C0334447|Malignant Cutaneous Blue Nevus
C0334447|Malignant Skin Blue Nevus
C0856900|sarcoma of skin (diagnosis)
C0856900|sarcoma of skin
C0856900|Cutaneous Sarcoma
C0856900|Sarcoma of the Skin
C0856900|Skin Sarcoma
C2211446|fibrosarcoma of skin (diagnosis)
C2211446|fibrosarcoma of skin
C2182812|dermatofibrosarcoma of skin
C2182812|dermatofibrosarcoma of skin (diagnosis)
C1333175|liposarcoma of skin (diagnosis)
C1333175|liposarcoma of skin
C1333175|Cutaneous Liposarcoma
C1333175|Liposarcoma of the Skin
C1333175|Skin Liposarcoma
C2211457|myosarcoma of skin
C2211457|myosarcoma of skin (diagnosis)
C1275281|carcinosarcoma of skin (diagnosis)
C1275281|carcinosarcoma of skin
C1275281|Carcinosarcoma of skin (disorder)
C2242810|malignant hemangioendothelioma of skin (diagnosis)
C2242810|malignant hemangioendothelioma of skin
C0346085|malignant hemangiopericytoma of skin (diagnosis)
C0346085|malignant hemangiopericytoma of skin
C0346085|Malignant Skin Hemangiopericytoma
C0346085|Malignant Hemangiopericytoma of the Skin
C0346085|Malignant haemangiopericytoma of skin
C0346085|Malignant hemangiopericytoma of skin (disorder)
C2211463|malignant neurilemoma of skin (diagnosis)
C2211463|malignant neurilemoma of skin
C2211464|malignant peripheral nerve sheath tumor (MPNST) of skin
C2211464|malignant peripheral nerve sheath tumor (MPNST) of skin (diagnosis)
C1321781|malignant mixed tumor of skin
C1321781|malignant mixed tumor of skin (diagnosis)
C1321781|Malignant chondroid syringoma
C1321781|Eccrine mixed tumor, malignant
C1321781|Eccrine mixed tumour, malignant
C1321781|Malignant chondroid syringoma (morphologic abnormality)
C1321781|Malignant chondroid syringoma of skin (disorder)
C1321781|Malignant chondroid syringoma of skin
C1321781|Malignant mixed tumor of the skin
C1321781|Malignant mixed tumour of the skin
C2211466|malignant lymphoma of skin (diagnosis)
C2211466|malignant lymphoma of skin
C1707551|Cutaneous Mature B-Cell Lymphocytic Neoplasm
C1707551|Cutaneous Mature B-Cell Neoplasm
C0948976|Leukemia Cutis
C0948976|Leukaemia cutis
C0948976|Leukemic infiltration of skin
C0948976|skin neoplasm malignant secondary leukemic infiltration
C0948976|Leukemic infiltration of skin (diagnosis)
C0948976|Leukaemic infiltration of skin
C0948976|Leukemic infiltration of skin (disorder)
C2211422|scirrhous adenocarcinoma of skin
C2211422|scirrhous adenocarcinoma of skin (diagnosis)
C2037356|superficial spreading adenocarcinoma of skin
C2037356|superficial spreading adenocarcinoma of skin (diagnosis)
C2145030|trabecular adenocarcinoma of skin (diagnosis)
C2145030|trabecular adenocarcinoma of skin
C0346017|adenoid cystic carcinoma of skin (diagnosis)
C0346017|adenoid cystic carcinoma of skin
C0346017|Adenoid cystic eccrine carcinoma of skin
C0346017|Adenoid cystic eccrine carcinoma of skin (diagnosis)
C0346017|skin neop malignant adnexa w/ eccrine differentiation adenoid cystic carcinoma
C0346017|Adenoid cystic eccrine carcinoma
C0346017|Primary cutaneous adenocystic carcinoma
C0346017|Adenoid cystic eccrine carcinoma (morphologic abnormality)
C0346017|Adenoid cystic eccrine carcinoma of skin (disorder)
C0346017|Adenoid cystic eccrine carcinoma (disorder)
C0346017|Adenoid Cystic Carcinoma of the Skin
C0346017|Adenoid Cystic Cutaneous Carcinoma
C0346017|Adenoid Cystic Skin Carcinoma
C2138462|cribriform carcinoma of skin
C2138462|cribriform carcinoma of skin (diagnosis)
C2017457|solid carcinoma of skin (diagnosis)
C2017457|solid carcinoma of skin
C2007050|carcinoma simplex of skin (diagnosis)
C2007050|carcinoma simplex of skin
C2033135|papillary adenocarcinoma of skin (diagnosis)
C2033135|papillary adenocarcinoma of skin
C2189650|villous adenocarcinoma of skin
C2189650|villous adenocarcinoma of skin (diagnosis)
C2211424|adenocarcinoma in villous adenoma of skin (diagnosis)
C2211424|adenocarcinoma in villous adenoma of skin
C2211425|adenocarcinoma in tubulovillous adenoma of skin (diagnosis)
C2211425|adenocarcinoma in tubulovillous adenoma of skin
C2075542|clear cell adenocarcinoma of skin (diagnosis)
C2075542|clear cell adenocarcinoma of skin
C0206697|Carcinoma, Skin Appendage
C0206697|Appendage Carcinoma, Skin
C0206697|Appendage Carcinomas, Skin
C0206697|Carcinomas, Skin Appendage
C0206697|Skin Appendage Carcinomas
C0206697|Skin Appendage Carcinoma
C0206697|skin appendage carcinoma (diagnosis)
C0206697|Carcinoma, Skin Appendage [Disease/Finding]
C0206697|[M]Skin appendage carcinoma
C0206697|[M]Skin appendage carcinoma (morphologic abnormality)
C0206697|CARCINOMA, ADNEXAL, MALIGNANT
C0206697|Carcinoma of Skin Appendage
C0206697|Carcinoma of Adnexa
C0206697|Adnexal carcinoma
C0206697|Skin appendage carcinoma (morphologic abnormality)
C2211430|sebaceous adenocarcinoma of skin (diagnosis)
C2211430|sebaceous adenocarcinoma of skin
C2026730|ceruminous adenocarcinoma of skin
C2026730|ceruminous adenocarcinoma of skin (diagnosis)
C2211431|mucinous adenocarcinoma of skin
C2211431|mucinous adenocarcinoma of skin (diagnosis)
C2211432|mucin-producing adenocarcinoma of skin (diagnosis)
C2211432|mucin-producing adenocarcinoma of skin
C1710103|Skin Adenosquamous Carcinoma
C1710103|adenosquamous carcinoma of skin
C1710103|adenosquamous carcinoma of skin (diagnosis)
C2211433|epithelial-myoepithelial carcinoma of skin
C2211433|epithelial-myoepithelial carcinoma of skin (diagnosis)
C2211434|adenocarcinoma of skin with metaplasia
C2211434|adenocarcinoma of skin with metaplasia (diagnosis)
C2211434|skin adenocarcinoma with metaplasia
C2211436|adenocarcinoma with cartilaginous or osseous metaplasia of skin
C2211436|skin adenocarcinoma with cartilaginous or osseous metaplasia
C2211436|adenocarcinoma of skin with cartilaginous and osseous metaplasia (diagnosis)
C2211436|adenocarcinoma of skin with cartilaginous and osseous metaplasia
C2211437|adenocarcinoma of skin with spindle cell metaplasia (diagnosis)
C2211437|adenocarcinoma of skin with spindle cell metaplasia
C2211438|adenocarcinoma of skin with apocrine metaplasia (diagnosis)
C2211438|adenocarcinoma of skin with apocrine metaplasia
C2211439|adenocarcinoma of skin with neuroendocrine differentiation
C2211439|adenocarcinoma of skin with neuroendocrine differentiation (diagnosis)
C2018514|spindle cell sarcoma of skin
C2018514|spindle cell sarcoma of skin (diagnosis)
C2011328|giant cell sarcoma of skin
C2011328|giant cell sarcoma of skin (diagnosis)
C2211445|small cell sarcoma of skin
C2211445|small cell sarcoma of skin (diagnosis)
C2188151|undifferentiated sarcoma of skin
C2188151|undifferentiated sarcoma of skin (diagnosis)
C2182958|desmoplastic small round cell sarcoma of skin (diagnosis)
C2182958|skin neoplasm malignant sarcoma desmoplastic small round cell
C2182958|desmoplastic small round cell sarcoma of skin
C2211447|fibromyxosarcoma of skin (diagnosis)
C2211447|fibromyxosarcoma of skin
C2211448|fascial fibrosarcoma of skin
C2211448|fascial fibrosarcoma of skin (diagnosis)
C2211449|infantile fibrosarcoma of skin (diagnosis)
C2211449|infantile fibrosarcoma of skin
C2211450|malignant solitary fibrous tumor of skin
C2211450|malignant solitary fibrous tumor of skin (diagnosis)
C2211451|well differentiated liposarcoma of skin
C2211451|well differentiated liposarcoma of skin (diagnosis)
C2211452|myxoid liposarcoma of skin
C2211452|myxoid liposarcoma of skin (diagnosis)
C2211453|round cell liposarcoma of skin
C2211453|round cell liposarcoma of skin (diagnosis)
C2211454|pleomorphic liposarcoma of skin
C2211454|pleomorphic liposarcoma of skin (diagnosis)
C2211455|mixed type liposarcoma of skin (diagnosis)
C2211455|mixed type liposarcoma of skin
C2211456|fibroblastic liposarcoma of skin (diagnosis)
C2211456|fibroblastic liposarcoma of skin
C2164525|dedifferentiated liposarcoma of skin (diagnosis)
C2164525|dedifferentiated liposarcoma of skin
C2200374|rhabdomyosarcoma of skin (diagnosis)
C2200374|rhabdomyosarcoma of skin
C2006989|carcinoma ex pleomorphic adenoma of skin (diagnosis)
C2006989|carcinoma ex pleomorphic adenoma of skin
C2211458|embryonal rhabdomyosarcoma of skin
C2211458|embryonal rhabdomyosarcoma of skin (diagnosis)
C2018456|spindle cell rhabdomyosarcoma of skin
C2018456|spindle cell rhabdomyosarcoma of skin (diagnosis)
C2211459|angiomyosarcoma of skin (diagnosis)
C2211459|angiomyosarcoma of skin
C2211460|embryonal carcinosarcoma of skin (diagnosis)
C2211460|embryonal carcinosarcoma of skin
C2211461|malignant myoepithelioma of skin
C2211461|malignant myoepithelioma of skin (diagnosis)
C0346081|hemangiosarcoma of skin (diagnosis)
C0346081|hemangiosarcoma of skin
C0346081|Skin angiosarcoma
C0346081|Cutaneous hemangiosarcoma
C0346081|Hemangiosarcoma of skin (disorder)
C0346081|malignant neoplasm sarcoma angiosarcoma of skin
C0346081|angiosarcoma of skin (diagnosis)
C0346081|angiosarcoma of skin
C0346081|Angiosarcoma of skin (disorder)
C0346081|Hemangiosarcoma of the Skin
C0346081|Angiosarcoma of the Skin
C0346081|Skin Hemangiosarcoma
C0030186|Extra Mammary Paget Disease
C0030186|Extra Mammary Paget's Disease
C0030186|Extra-Mammary Pagets Disease
C0030186|Extramammary Pagets Disease
C0030186|Paget Disease, Extra Mammary
C0030186|Paget's Disease, Extra Mammary
C0030186|Pagets Disease, Extra-Mammary
C0030186|Pagets Disease, Extramammary
C0030186|Cutaneous Paget's Disease
C0030186|Paget's Disease of Skin
C0030186|Paget's Disease of the Skin
C0030186|Paget's Skin Disease
C0030186|PAGET DISEASE, EXTRAMAMMARY
C0030186|PAGETS DIS EXTRA MAMMARY
C0030186|PAGETS DIS EXTRAMAMMARY
C0030186|EXTRAMAMMARY PAGETS DIS
C0030186|PAGET DIS EXTRA MAMMARY
C0030186|EXTRA MAMMARY PAGET DIS
C0030186|EXTRAMAMMARY PAGET DIS
C0030186|PAGET DIS EXTRAMAMMARY
C0030186|EXTRA MAMMARY PAGETS DIS
C0030186|Extramammary Paget's Disease
C0030186|Extramammary Paget Disease
C0030186|extramammary Paget's disease (diagnosis)
C0030186|Extramammary, Paget Disease
C0030186|Paget Disease Extramammary
C0030186|Paget disease of skin
C0030186|Paget disease, extramammary (except Paget disease of bone)
C0030186|Extra-Mammary Paget Disease
C0030186|Extra-Mammary Paget's Disease
C0030186|Paget Disease, Extra-Mammary
C0030186|Paget's Disease, Extra-Mammary
C0030186|Paget's Disease, Extramammary
C0030186|Paget Disease, Extramammary [Disease/Finding]
C0030186|Extramammary Paget's disease (morphologic abnormality)
C0030186|[M]Paget's disease, extramammary, excluding Paget's disease of bone
C0030186|Paget's disease, extramammary (except Paget's disease of bone)
C0030186|Paget's disease of skin (morphologic abnormality)
C0030186|Paget's disease, extramammary (except Paget's disease of bone) (morphologic abnormality)
C0030186|[M]Paget's disease, extramammary, excluding Paget's disease of bone (morphologic abnormality)
C3251593|skin neoplasm location malignant (diagnosis)
C3251593|skin neoplasm location malignant
C3251594|skin neoplasm location malignant basal cell carcinoma
C3251594|skin neoplasm location malignant basal cell carcinoma (diagnosis)
C3251595|skin neoplasm location malignant squamous cell carcinoma
C3251595|skin neoplasm location malignant squamous cell carcinoma (diagnosis)
C0375068|Other malignant neoplasm of skin, site unspecified
C0553723|Squamous cell carcinoma of skin
C0553723|Squamous cell carcinoma of the skin
C0553723|squamous cell carcinoma of skin (diagnosis)
C0553723|Squamous cell carcinoma - skin
C0553723|Squamous skin carcinoma
C0553723|Spinous cell carcinoma
C0553723|Cutaneous squamous cell carcinoma
C0553723|SCC - Cutaneous squamous cell carcinoma
C0553723|SCC - Squamous cell carcinoma of skin
C0553723|Squamous cell carcinoma of skin (disorder)
C0553723|cancer of the skin, squamous cell
C0553723|carcinoma of the skin, squamous cell
C0553723|carcinoma, epidermoid, skin
C0553723|carcinoma, squamous cell, skin
C0553723|epidermoid carcinoma of the skin
C0553723|skin cancer, epidermoid carcinoma
C0553723|skin cancer, squamous cell
C0553723|Epidermoid Carcinoma of Skin
C0553723|Epidermoid Skin Carcinoma
C0553723|Skin Squamous Cell Carcinoma
C0553723|Squamous Cell Skin Carcinoma
C0007117|Basal cell carcinoma
C0007117|BASAL CELL CARCINOMA OF SKIN
C0007117|Basal Cell Carcinomas
C0007117|Basal Cell Epitheliomas
C0007117|Carcinoma, Basal Cell
C0007117|Carcinomas, Basal Cell
C0007117|Epitheliomas, Basal Cell
C0007117|Basal Cell Epithelioma
C0007117|Rodent Ulcers
C0007117|Ulcers, Rodent
C0007117|basal cell carcinoma of skin (diagnosis)
C0007117|Carcinoma, Basal Cell [Disease/Finding]
C0007117|Epithelioma, Basal Cell
C0007117|Rodent Ulcer
C0007117|Ulcer, Rodent
C0007117|Ulcer;rodent
C0007117|[M]Basal cell carcinoma NOS (morphologic abnormality)
C0007117|[M]Basal cell carcinoma NOS
C0007117|Epithelioma basal cell
C0007117|Basal cell epithelioma (diagnosis)
C0007117|malignant neoplasm carcinoma epithelioma basal cell
C0007117|basal cell cancer
C0007117|Basalioma
C0007117|Cancer of skin, basal cell
C0007117|Carcinoma basal cell
C0007117|BCC - Basal cell carcinoma
C0007117|BCC - Basal cell carcinoma of skin
C0007117|Basiloma
C0007117|RU - Rodent ulcer
C0007117|Epithelioma basal cell (disorder)
C0007117|Basal cell carcinoma (morphologic abnormality)
C0007117|Basal cell carcinoma of skin (disorder)
C0007117|basal cell carcinoma of the skin
C0007117|carcinoma of the skin, basal cell
C0007117|carcinoma, basal cell, skin
C0007117|Basal cell carcinoma, NOS
C0007117|BCC
C0007117|Basal Cell Skin Carcinoma
C0007117|Skin Basal Cell Carcinoma
C1261513|skin neoplasm nose malignant primary
C1261513|Primary malignant neoplasm of skin of nose
C1261513|Primary malignant neoplasm of skin of nose (diagnosis)
C1261513|Primary malignant neoplasm of skin of nose (disorder)
C1314758|Primary malignant neoplasm of skin (diagnosis)
C1314758|Primary malignant neoplasm of skin
C1314758|skin neoplasm malignant primary
C1314758|Primary malignant neoplasm of skin (disorder)
C0348363|Malignant neoplasm overlapping skin site
C0348363|Overlapping lesion of skin
C0348363|malignant neoplasm of overlapping sites of skin (diagnosis)
C0348363|skin neoplasm malignant overlapping sites
C0348363|malignant neoplasm of overlapping sites of skin
C0348363|[X]Malignant neoplasm overlapping lesion of skin
C0348363|[X]Malignant neoplasm overlapping lesion of skin (disorder)
C0153346|Malignant neoplasm of commissure of lip
C0153346|Commissure of lip
C0153346|lip neoplasm malignant labial commissure
C0153346|Mal neo lip, commissure
C0153346|Malignant tumour of commissure of lip
C0153346|Malignant tumor of commissure of lip
C0153346|Malignant tumor of labial commissure
C0153346|Malignant tumour of labial commissure
C0153346|malignant neoplasm of labial commissure
C0153346|malignant neoplasm of commissure of lip (diagnosis)
C0153346|Malignant tumor of commissure of lip (disorder)
C0153346|Malignant neoplasm of labial commissure of lip
C0346735|malignant skin neoplasm of cheek (external)
C0346735|malignant skin neoplasm of cheek (external) (diagnosis)
C0346735|Malignant neoplasm of skin of cheek, external (disorder)
C0346735|Malignant neoplasm of skin of cheek, external
C0346026|Benign Mixed Tumor of the Skin (Chondroid Syringoma)
C0346026|Mixed Tumor of the Skin (Chondroid Syringoma)
C0346026|Eccrine mixed tumor of skin
C0346026|Eccrine mixed tumour of skin
C0346026|Eccrine mixed tumor
C0346026|Eccrine mixed tumour
C0346026|Mixed tumor of skin
C0346026|Mixed tumour of skin
C0346026|Eccrine mixed tumor (morphologic abnormality)
C0346026|Eccrine mixed tumor of skin (disorder)
C0346026|Eccrine mixed tumor (disorder)
C0346026|Chondroid Syringoma
C0346026|Benign Mixed Tumor of Skin (Chondroid Syringoma)
C0346026|Benign Mixed Tumor of Skin
C0346026|Benign Mixed Tumor of the Skin
C1275323|Primary cutaneous plasmacytoma (diagnosis)
C1275323|Primary cutaneous plasmacytoma
C1275323|skin malignant lymphoma non-hodgkin's primary cutaneous plasmacytoma
C1275323|Primary cutaneous plasmacytic B-cell lymphoma
C1275323|Primary cutaneous plasmacytoma (disorder)
C1275323|Primary cutaneous plasmacytoma (morphologic abnormality)
C1275318|Angiocentric natural killer/T-cell malignant lymphoma involving skin
C1275318|Angiocentric NK/T-cell malignant lymphoma involving skin (disorder)
C1275318|Angiocentric natural killer/T-cell malignant lymphoma involving skin (disorder)
C1275318|Angiocentric NK/T-cell malignant lymphoma involving skin
C1275318|skin malignant lymphoma non-hodgkin's angiocentric nk/t-cell
C1275318|Angiocentric NK/T-cell malignant lymphoma involving skin (diagnosis)
C1275318|Angiocentric lymphoma involving skin
C3489398|NEUROEPITHELIOMA, PERIPHERAL
C3489398|PNE
C3489398|skin neoplasm malignant primary peripheral neuroepithelioma
C3489398|Peripheral neuroepithelioma
C3489398|Peripheral neuroepithelioma (diagnosis)
C3489398|PNE - Peripheral neuroepithelioma
C3489398|Peripheral neuroepithelioma (disorder)
C0346770|Malignant skin tumour with adnexal differentiation
C0346770|Malignant skin tumor with adnexal differentiation
C0346770|Malignant tumor of epidermal appendage
C0346770|Malignant tumour of epidermal appendage
C0346770|Malignant skin tumor with adnexal differentiation (disorder)
C0346770|Malignant tumor of epidermal appendage (disorder)
C0346770|Malignant Cutaneous Adnexal Neoplasm
C0346770|Malignant Epidermal Appendage Neoplasm
C0346770|Malignant Epidermal Appendage Tumor
C0346770|Malignant Neoplasm of Epidermal Appendage
C0346770|Malignant Neoplasm of the Epidermal Appendage
C0346770|Malignant Skin Adnexal Neoplasm
C0346770|Malignant Skin Adnexal Tumor
C0346770|Malignant Skin Appendage Neoplasm
C0346770|Malignant Tumor of the Epidermal Appendage
C0346728|Malignant neoplasm of skin of external auditory meatus
C0346728|Malignant neoplasm of skin of external auditory meatus (disorder)
C0346079|Proliferating angioendotheliomatosis
C0346079|non-hodgkin's lymphoma of skin proliferating angioendotheliomatosis
C0346079|Proliferating angioendotheliomatosis (diagnosis)
C0346079|Proliferating angioendotheliomatosis (disorder)
C0346024|Eccrine Dermal Duct Neoplasm
C0346024|Dermal Duct Tumor
C0346024|Eccrine dermal duct tumour of skin
C0346024|Eccrine dermal duct tumor of skin
C0346024|Dermal duct tumor (morphologic abnormality)
C0346024|Dermal duct tumour
C0346024|Eccrine dermal duct tumor
C0346024|Eccrine dermal duct tumour
C0346024|Eccrine dermal duct tumor of skin (disorder)
C0346024|Eccrine dermal duct tumor (disorder)
C0346024|Dermal Duct Neoplasm
C0684352|Malignant neoplasm of adnexa of skin
C0684352|Primary malignant neoplasm of skin with adnexal differentiation
C0684352|primary malignant neoplasm of skin adnexa
C0684352|primary malignant neoplasm of skin adnexa (diagnosis)
C0684352|skin neoplasm malignant adnexa
C0684352|malignant neoplasm of skin adnexa (diagnosis)
C0684352|malignant neoplasm of skin adnexa
C0684352|skin neoplasm malignant adnexa primary
C0684352|Primary malignant neoplasm of adnexa of skin
C0684352|Primary malignant neoplasm of skin with adnexal differentiation (disorder)
C0684352|Primary malignant neoplasm of adnexa of skin (disorder)
C1304523|Aggressive natural killer-cell leukemia involving skin
C1304523|Aggressive NK-cell leukemia involving skin (disorder)
C1304523|Aggressive natural killer-cell leukemia involving skin (disorder)
C1304523|Aggressive NK-cell leukemia involving skin (diagnosis)
C1304523|malignant neoplasm lymphoma agressive nk-cell involving skin
C1304523|Aggressive NK-cell leukemia involving skin
C1304523|Aggressive natural killer-cell leukaemia involving skin
C1304523|Aggressive NK-cell leukaemia involving skin
C2314897|Skin Squamous Cell Carcinoma In Situ
C2314897|Squamous cell carcinoma in situ of skin
C2314897|Squamous cell carcinoma in situ of skin (disorder)
C2314897|Cancer in situ skin, squamous cell
C2314897|Intraepidermal squamous cell carcinoma
C2314897|Squamous cell carcinoma of skin in situ
C2314897|IEC - Intraepidermal carcinoma of skin
C2314897|Intraepidermal carcinoma of skin
C2314897|SCC - Squamous cell carcinoma in situ of skin
C2314897|Squamous Cell Carcinoma in situ of the Skin
C0346734|malignant neoplasm of skin of temple (diagnosis)
C0346734|malignant neoplasm of skin of temple
C0346734|skin neoplasm temple malignant
C0346734|Malignant neoplasm of skin of temple (disorder)
C0346082|Stewart-Treves syndrome
C0346082|Postmastectomy extremity angiosarcoma
C0346082|Angiosarcoma associated with chronic lymphedema
C0346082|Lymphangiosarcoma following mastectomy
C0346082|Stewart Treves syndrome
C0346082|Stewart-Treves syndrome (diagnosis)
C0346082|benign neoplasm stewart-treves syndrome
C0346082|Postmastectomy lymphangiosarcoma syndrome
C0346082|Lymphangiosarcoma of Stewart and Treves
C0346082|Lymphangiosarcoma of skin
C0346082|Stewart-Treves syndrome (disorder)
C0346082|Lymphangiosarcoma of the Skin
C0346082|Skin Lymphangiosarcoma
C0346769|Malignant neoplasm of other specified skin sites (disorder)
C0346769|Malignant neoplasm of other specified skin sites
C0559018|Ca skin - other
C0559018|Ca skin - other NOS (disorder)
C0559018|Ca skin - other NOS
C3665499|Malignant neoplasm of skin of elbow
C3665499|skin neoplasm elbow malignant
C3665499|malignant neoplasm of skin of elbow (diagnosis)
C3665401|Malignant neoplasm of skin of thigh (disorder)
C3665401|Malignant neoplasm of skin of thigh
C3665401|malignant neoplasm of skin of thigh (diagnosis)
C2210570|skin biopsy specimen malignant neoplasm (procedure)
C2210570|skin biopsy specimen malignant neoplasm
C3665399|Malignant neoplasm of skin of hand
C3665399|Malignant neoplasm of skin of hand (disorder)
C3665399|skin neoplasm hand malignant
C3665399|malignant skin neoplasm of hand
C3665399|malignant skin neoplasm of hand (diagnosis)
C1282486|skin neoplasm malignant, local recurrence
C1282486|local recurrence of malignant skin neoplasm
C1282486|local recurrence of malignant skin neoplasm (diagnosis)
C1282486|Local recurrence of malignant tumor of skin (disorder)
C1282486|Local recurrence of malignant tumor of skin
C1282486|Local recurrence of malignant tumour of skin
C1304404|malignant vascular neoplasm of skin (diagnosis)
C1304404|malignant vascular neoplasm of skin
C1304404|skin malignant neoplasm vascular
C1304404|Malignant vascular tumor of skin (disorder)
C1304404|Malignant vascular tumor of skin
C1304404|Malignant vascular tumour of skin
C1304404|Malignant Cutaneous Vascular Neoplasm
C1304404|Malignant Cutaneous Vascular Tumor
C1304404|Malignant Skin Vascular Neoplasm
C1304404|Malignant Skin Vascular Tumor
C1282490|metastasis from malignant neoplasm of skin (diagnosis)
C1282490|metastasis from malignant neoplasm of skin
C1282490|skin neoplasm malignant metastasis
C1282490|Metastasis from malignant tumor of skin (disorder)
C1282490|Metastasis from malignant tumor of skin
C1282490|Metastasis from malignant tumour of skin
C0346031|malignant neoplasm of skin with apocrine differentiation
C0346031|skin neoplasm malignant with apocrine differentiation
C0346031|malignant neoplasm of skin with apocrine differentiation (diagnosis)
C0346031|Malignant skin tumor with apocrine differentiation
C0346031|Malignant skin tumour with apocrine differentiation
C0346031|Malignant skin tumor with apocrine differentiation (disorder)
C1304452|malignant fibrohistiocytic neoplasm of skin
C1304452|malignant fibrohistiocytic neoplasm of skin (diagnosis)
C1304452|skin neoplasm malignant fibrohistiocytic
C1304452|Malignant fibrohistiocytic tumor of skin (disorder)
C1304452|Malignant fibrohistiocytic tumor of skin
C1304452|Malignant fibrohistiocytic tumour of skin
C0346811|skin neoplasm malignant dermis
C0346811|malignant neoplasm of dermis
C0346811|malignant neoplasm of dermis (diagnosis)
C0346811|Malignant tumor of dermis
C0346811|Malignant tumour of dermis
C0346811|Malignant tumor of dermis (disorder)
C0346811|Malignant Dermal Neoplasm
C0346811|Malignant Dermis Neoplasm
C0346811|Malignant Dermis Tumor
C0346811|Malignant Neoplasm of the Dermis
C0346811|Malignant Tumor of the Dermis
C1275031|PUVA therapy-associated skin malignancy (disorder)
C1275031|Psoralen and long-wave ultraviolet radiation (PUVA) therapy-associated skin malignancy
C1275031|Psoralen and long-wave ultraviolet radiation (PUVA) therapy-associated skin malignancy (disorder)
C1275031|Psoralen and long-wave ultraviolet radiation therapy-associated skin malignancy (disorder)
C1275031|Psoralen and long-wave ultraviolet radiation therapy-associated skin malignancy
C1275031|Psoralen and long-wave ultraviolet radiation therapy-associated skin malignancy (diagnosis)
C1275031|skin neoplasm malignant psoralen/long-wave ultraviolet radiation therapy assoc
C1275031|PUVA therapy-associated skin malignancy
C1275046|Radiation-induced skin malignancy
C1275046|skin neoplasm malignant radiation-induced
C1275046|Radiation-induced skin malignancy (diagnosis)
C1275046|Radiation-induced skin malignancy (disorder)
C1275056|arsenic-induced malignancy
C1275056|skin neoplasm malignant arsenic-induced
C1275056|arsenic-induced malignancy (diagnosis)
C1275056|Arsenic-induced skin malignancy (disorder)
C1275056|Arsenic-induced skin malignancy
C1998037|Malignant basal cell tumor of skin
C1998037|Malignant basal cell neoplasm of skin
C1998037|Malignant basal cell tumour of skin
C1998037|Malignant basal cell neoplasm of skin (disorder)
C1998037|malignant basal cell neoplasm of skin (diagnosis)
C1998037|skin malignant neoplasm basal cell
C0153687|Secondary malignant neoplasm of skin
C0153687|Metastatic Neoplasm to the Skin
C0153687|metastasis of malignant neoplasm to skin (diagnosis)
C0153687|metastasis to the skin
C0153687|metastasis of malignant neoplasm to skin
C0153687|Metastases to skin
C0153687|Secondary malig neo skin
C0153687|secondary malignant neoplasm of skin (diagnosis)
C0153687|secondary malignant neoplasm skin
C0153687|Secondary malignant neoplasm of skin NOS (disorder)
C0153687|Metastasis to skin (disorder)
C0153687|Skin cancer metastatic
C0153687|Metastasis to skin
C0153687|Secondary malignant neoplasm of skin NOS
C0153687|Metastases to skin, NOS
C0153687|Metastatic Malignant Neoplasm to the Skin
C0153687|Metastatic Malignant Neoplasm in the Skin
C0153687|Cancer metastatic to skin
C0153687|Skin metastases
C0153687|Cutaneous metastasis
C0153687|Dermal metastasis
C0153687|Malignant infiltration of skin
C0153687|Skin secondaries
C0153687|Secondary cancer of skin
C0153687|Metastatic malignant neoplasm to skin
C0153687|Secondary malignant neoplasm of skin (disorder)
C0153687|cancer, metastatic to skin
C0153687|metastatic cancer to skin
C0153687|skin, metastatic cancer to
C0153687|Metastatic malignant neoplasm to skin, NOS
C0153687|Secondary malignant neoplasm of skin, NOS
C0153687|Metastatic Tumor to the Skin
C0153687|Skin Metastasis
C0349513|skin neoplasm malignant with pilar differentiation (diagnosis)
C0349513|skin neoplasm malignant with pilar differentiation
C0349513|Malignant tumor of skin with pilar differentiation
C0349513|Malignant tumour of skin with pilar differentiation
C0349513|Malignant tumor of skin with pilar differentiation (disorder)
C0547064|Malignant skin tumor with eccrine differentiation
C0547064|malignant skin neoplasm with eccrine differentiation
C0547064|skin neoplasm malignant adnexa with eccrine differentiation
C0547064|malignant skin neoplasm with eccrine differentiation (diagnosis)
C0547064|Malignant skin tumour with eccrine differentiation
C0547064|Malignant sweat gland tumor
C0547064|Malignant sweat gland tumour
C0547064|Malignant skin tumor with eccrine differentiation (disorder)
C0496797|Skin of trunk
C0496797|Malignant neoplasm of skin of trunk
C0496797|malignant neoplasm of skin of trunk (diagnosis)
C0496797|skin neoplasm trunk malignant
C0496797|Ca skin - trunk (disorder)
C0496797|Ca skin - trunk
C0496797|Malignant neoplasm of skin of trunk (disorder)
C0496797|Malignant neoplasm of skin of trunk, NOS
C0345977|Malignant tumor of surface epithelium
C0345977|Malignant tumour of surface epithelium
C0345977|Malignant epithelial neoplasm of skin (disorder)
C0345977|Malignant epithelial neoplasm of skin
C0345977|Malignant tumor of surface epithelium (disorder)
C1269827|malignant skin neoplasm of head and neck (diagnosis)
C1269827|malignant skin neoplasm of head and neck
C1269827|skin neoplasm head and neck malignant
C1269827|Ca skin - head/neck
C1269827|Malignant neoplasm of skin head and neck (disorder)
C1269827|Malignant neoplasm of skin head and neck
C0559017|skin neoplasm lower extremities malignant
C0559017|malignant neoplasm of skin of lower extremities (diagnosis)
C0559017|malignant neoplasm of skin of lower extremities
C0559017|Ca skin - lower limb (disorder)
C0559017|Ca skin - lower limb
C0559017|Malignant neoplasm of skin of lower limb (disorder)
C0559017|Malignant neoplasm of skin of lower limb
C0684431|Malignant neoplasm of skin of upper limb
C0684431|Malignant neoplasm of skin of arm
C0684431|skin neoplasm upper extremities malignant
C0684431|malignant neoplasm of skin of upper extremities (diagnosis)
C0684431|malignant neoplasm of skin of upper extremities
C0684431|Ca skin - upper limb
C0684431|Ca skin - upper limb (disorder)
C0684431|Malignant neoplasm of skin of upper limb (disorder)
C0684431|Malignant neoplasm of skin of upper limb, NOS
C1274311|Hodgkin disease affecting skin
C1274311|Hodgkin's disease affecting skin (diagnosis)
C1274311|Hodgkin's disease affecting skin
C1274311|Hodgkin's disease affecting skin (disorder)
C1275320|small B-cell lymphocytic lymphoma of skin (diagnosis)
C1275320|small B-cell lymphocytic lymphoma of skin
C1275320|Small lymphocytic B-cell lymphoma involving skin (disorder)
C1275320|Small lymphocytic B-cell lymphoma involving skin
C0334346|apocrine adenocarcinoma
C0334346|apocrine adenocarcinoma (diagnosis)
C0334346|Apocrine adenocarcinoma (morphologic abnormality)
C0334346|adenocarcinoma; apocrine, unspecified site
C0334346|apocrine; adenocarcinoma, unspecified site
C1388303|carcinoma; apocrine, unspecified site
C1388303|apocrine; carcinoma, unspecified site
C1395263|dermatofibrosarcoma; (site of skin not specified)
C0392784|dermatofibrosarcoma protuberans
C0392784|Dermatofibrosarcoma protuberans (disorder)
C0392784|Dermatofibrosarcoma
C0392784|Dermatofibrosarcoma protuberans (diagnosis)
C0392784|soft tissue malignant neoplasm dermatofibrosarcoma protuberans
C0392784|[M]Dermatofibroma protuberans
C0392784|DFSP - Dermatofibrosarcoma protruberans
C0392784|Dermatofibrosarcoma (morphologic abnormality)
C0392784|dermatofibrosarcoma; protuberans
C0392784|protuberans; dermatofibrosarcoma
C0392784|Dermatofibrosarcoma protuberans, NOS
C0392784|DFSP
C0280247|stage/cell type, skin cancer
C0280247|skin cancer stage
C1302772|Primary Cutaneous Lymphoma
C1302772|skin malignant lymphoma primary cutaneous
C1302772|Primary cutaneous lymphoma (diagnosis)
C1302772|Primary cutaneous lymphoma (disorder)
C1302772|Cutaneous Lymphoma
C1302772|Skin Lymphoma
C1302772|Primary cutaneous lymphoma (morphologic abnormality)
C0153604|Scrotum
C0153604|Malignant neoplasm of scrotum
C0153604|malignant neoplasm of scrotum (diagnosis)
C0153604|Scrotal cancer
C0153604|malignant tumor of scrotum
C0153604|Malign neopl scrotum
C0153604|Malignant tumour of scrotum
C0153604|Malignant tumour of scrotum (disorder)
C0153604|CA - Cancer of scrotum
C0153604|Cancer of scrotum
C0153604|Scrotal Ca
C0153604|Malignant scrotal tumor
C0153604|Malignant scrotal tumour
C0153604|Malignant tumor of scrotum (disorder)
C0153604|Malignant Neoplasm of the Scrotum
C0153604|Malignant Scrotal Neoplasm
C0153604|Malignant Tumor of the Scrotum
C1707590|Cutaneous Precursor Lymphoblastic Lymphoma/Leukemia
C1707590|Cutaneous Precursor Lymphoid Neoplasm
C1301363|Blastic NK-Cell Lymphoma
C1301363|Early Plasmacytoid Dendritic Cell Leukemia/Lymphoma
C1301363|Primary Cutaneous CD4+/CD56+ Hematolymphoid Neoplasm
C1301363|Blastic Natural Killer Leukemia/Lymphoma
C1301363|CD4+/CD56+ Hematodermic Neoplasm
C1301363|Agranular CD4+ CD56+ Hematodermic Neoplasm/Tumor
C1301363|Blastic Plasmacytoid Dendritic Cell Neoplasm
C1301363|Agranular CD4+ Natural Killer Cell Leukemia
C1301363|Blastic plasmacytoid dendritic cell neoplasm (morphologic abnormality)
C1301363|Blastic plasmacytoid dendritic cell neoplasm (disorder)
C1301363|malignant neoplasm lymphoma nk-cell blastic
C1301363|Blastic NK-cell lymphoma (diagnosis)
C1301363|Blastic NK-cell lymphoma (morphologic abnormality)
C1301363|neoplasm of hematopoietic cell type blastic plasmacytoid dendritic cell
C1301363|Blastic plasmacytoid dendritic cell neoplasm (diagnosis)
C1301363|Monomorphic NK-Cell Lymphoma
C2211472|nodular sclerosing Hodgkin's lymphoma of skin (diagnosis)
C2211472|nodular sclerosing Hodgkin's lymphoma of skin
C2211475|grade 2 nodular sclerosing Hodgkin's lymphoma of skin
C2211475|grade 2 nodular sclerosing Hodgkin's lymphoma of skin (diagnosis)
C2046521|skin malignant lymphoma Hodgkin's and non-Hodgkin's
C2046521|composite Hodgkin's and non-Hodgkin's lymphoma of skin
C2046521|composite Hodgkin's and non-Hodgkin's lymphoma of skin (diagnosis)
C2211476|lymphoplasmacytic lymphoma of skin (diagnosis)
C2211476|lymphoplasmacytic lymphoma of skin
C2211477|mantle cell lymphoma of skin
C2211477|mantle cell lymphoma of skin (diagnosis)
C2211483|grade 2 follicular lymphoma of skin (diagnosis)
C2211483|grade 2 follicular lymphoma of skin
C2211486|angioimmunoblastic T-cell lymphoma of skin (diagnosis)
C2211486|angioimmunoblastic T-cell lymphoma of skin
C2211486|angioimmunoblastic lymphadenopathy with dysproteinemia (AILD) of skin
C2211471|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of skin (diagnosis)
C2211471|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of skin
C2211474|grade 1 nodular sclerosing Hodgkin's lymphoma of skin (diagnosis)
C2211474|grade 1 nodular sclerosing Hodgkin's lymphoma of skin
C2211479|immunoblastic large B-cell diffuse lymphoma of skin (diagnosis)
C2211479|immunoblastic large B-cell diffuse lymphoma of skin
C2211484|grade 3 follicular lymphoma of skin
C2211484|grade 3 follicular lymphoma of skin (diagnosis)
C2046594|Hodgkin's granuloma of skin
C2046594|Hodgkin's granuloma of skin (diagnosis)
C1367653|Primary Cutaneous Marginal Zone B Cell Lymphoma of Mucosa-Associated Lymphoid Tissue
C1367653|marginal zone B-cell lymphoma of skin (diagnosis)
C1367653|marginal zone B-cell lymphoma of skin
C1367653|Primary Cutaneous Marginal Zone Lymphoma of Mucosa-Associated Lymphoid Tissue
C1367653|Primary Cutaneous Marginal Zone B-Cell Lymphoma of Mucosa-Associated Lymphoid Tissue
C1367653|SALT lymphoma
C1367653|Skin-associated lymphoid tissue lymphoma
C1367653|Cutaneous Immunocytoma
C1367653|Marginal Zone B Cell Lymphoma of Skin
C1367653|Marginal Zone B Cell Lymphoma of the Skin
C1367653|C-MALT
C2211488|subcutaneous panniculitis-like T-cell lymphoma of skin (diagnosis)
C2211488|subcutaneous panniculitis-like T-cell lymphoma of skin
C2211469|mixed cellularity Hodgkin's lymphoma of skin
C2211469|mixed cellularity Hodgkin's lymphoma of skin (diagnosis)
C2211473|nodular sclerosing Hodgkin's lymphoma in cellular phase of skin
C2211473|nodular sclerosing Hodgkin's lymphoma in cellular phase of skin (diagnosis)
C2211485|mature T-cell lymphoma of skin (diagnosis)
C2211485|mature T-cell lymphoma of skin
C2211470|Hodgkin's disease, lymphocytic depletion of skin
C2211470|Hodgkin's disease, lymphocytic depletion of skin (diagnosis)
C2046734|Hodgkin's sarcoma of skin
C2046734|Hodgkin's sarcoma of skin (diagnosis)
C2211482|grade 1 follicular lymphoma of skin (diagnosis)
C2211482|grade 1 follicular lymphoma of skin
C2211468|lymphocyte-rich Hodgkin's lymphoma of skin (diagnosis)
C2211468|lymphocyte-rich Hodgkin's lymphoma of skin
C2211478|large B-cell diffuse lymphoma of skin (diagnosis)
C2211478|large B-cell diffuse lymphoma of skin
C0238461|Anaplastic Thyroid Carcinoma
C0238461|Thyroid Gland Carcinosarcoma
C0238461|Thyroid Gland Undifferentiated (Anaplastic) Carcinoma
C0238461|Undifferentiated (Anaplastic) Thyroid Gland Carcinoma
C0238461|Dedifferentiated Thyroid Gland Carcinoma
C0238461|Metaplastic Thyroid Gland Carcinoma
C0238461|Pleomorphic Thyroid Gland Carcinoma
C0238461|Sarcomatoid Thyroid Gland Carcinoma
C0238461|carcinosarcoma of thyroid gland
C0238461|carcinosarcoma of thyroid gland (diagnosis)
C0238461|Anaplastic thyroid cancer
C0238461|undifferentiated carcinoma of thyroid gland
C0238461|anaplastic carcinoma of thyroid gland
C0238461|anaplastic thyroid carcinoma (diagnosis)
C0238461|undifferentiated carcinoma of the thyroid gland
C0238461|undifferentiated carcinoma of the thyroid gland (diagnosis)
C0238461|Anaplastic Thyroid Carcinomas
C0238461|Cancers, Anaplastic Thyroid
C0238461|Thyroid Cancers, Anaplastic
C0238461|Thyroid Carcinoma, Anaplastic
C0238461|Carcinoma, Anaplastic Thyroid
C0238461|Anaplastic Thyroid Cancers
C0238461|Thyroid Carcinomas, Anaplastic
C0238461|Cancer, Anaplastic Thyroid
C0238461|Carcinomas, Anaplastic Thyroid
C0238461|Thyroid Carcinoma, Anaplastic [Disease/Finding]
C0238461|Thyroid Cancer, Anaplastic
C0238461|Anaplastic thyroid carcinoma (disorder)
C0238461|anaplastic carcinoma of the thyroid
C0238461|thyroid cancer, anaplastic carcinoma
C0238461|thyroid cancer, undifferentiated carcinoma
C0238461|undifferentiated carcinoma of the thyroid
C0238461|undifferentiated thyroid cancer
C0238461|Anaplastic Carcinoma of Thyroid
C0238461|Anaplastic Carcinoma of the Thyroid Gland
C0238461|Anaplastic Thyroid Gland Carcinoma
C0238461|Undifferentiated Carcinoma of Thyroid
C0238461|Undifferentiated Thyroid Carcinoma
C0238461|Undifferentiated Thyroid Gland Carcinoma
C0206682|Adenocarcinoma, Follicular
C0206682|Adenocarcinomas, Follicular
C0206682|Follicular Adenocarcinomas
C0206682|Follicular Adenocarcinoma
C0206682|Follicular Thyroid Carcinoma
C0206682|Thyroid Gland Follicular Carcinoma
C0206682|Follicular Thyroid Gland Carcinoma
C0206682|THYROID CARCINOMA, FOLLICULAR
C0206682|FTC
C0206682|follicular adenocarcinoma of thyroid gland
C0206682|follicular adenocarcinoma of thyroid gland (diagnosis)
C0206682|Follicular thyroid cancer
C0206682|Adenocarcinoma, Follicular [Disease/Finding]
C0206682|Carcinoma, Follicular Thyroid
C0206682|Carcinomas, Follicular Thyroid
C0206682|Follicular Thyroid Carcinomas
C0206682|Thyroid Carcinomas, Follicular
C0206682|[M]Follicular adenocarcinoma NOS (morphologic abnormality)
C0206682|[M]Follicular adenocarcinoma NOS
C0206682|[M]Follicular carcinoma
C0206682|CARCINOMA, FOLLICULAR CELL, MALIGNANT
C0206682|follicular thyroid carcinoma (diagnosis)
C0206682|thyroid malignant carcinoma follicualr
C0206682|Follicular Carcinoma of Thyroid Gland
C0206682|Follicular Cancer of Thyroid
C0206682|Follicular Carcinoma of the Thyroid Gland
C0206682|Follicular Carcinoma
C0206682|Follicular Carcinoma of the Thyroid
C0206682|Well-differentiated Follicular Adenocarcinoma
C0206682|Well-differentiated Follicular Carcinoma
C0206682|Follicular Carcinoma of Thyroid
C0206682|Follicular Cancer of the Thyroid
C0206682|Thyroid Follicular Carcinoma
C0206682|Follicular Cancer of Thyroid Gland
C0206682|Follicular Cancer of the Thyroid Gland
C0206682|Follicular adenocarcinoma - well differentiated
C0206682|Follicular adenocarcinoma, well differentiated
C0206682|Follicular carcinoma - well differentiated
C0206682|Follicular carcinoma, well differentiated
C0206682|FTC - Follicular thyroid carcinoma
C0206682|Follicular adenocarcinoma (morphologic abnormality)
C0206682|Follicular adenocarcinoma, well differentiated (morphologic abnormality)
C0206682|Follicular thyroid carcinoma (disorder)
C0206682|thyroid cancer, follicular
C0206682|carcinoma; follicular, pure
C0206682|carcinoma; follicular, well differentiated
C0206682|follicular; adenocarcinoma, well differentiated
C0206682|follicular; carcinoma, well differentiated
C0206682|adenocarcinoma; follicular, well differentiated
C0206682|Follicular adenocarcinoma, NOS
C0206682|Follicular carcinoma, NOS
C0238462|medullary thyroid carcinoma
C0238462|Thyroid Gland Medullary Carcinoma
C0238462|Thyroid Gland Neuroendocrine Carcinoma
C0238462|Medullary Thyroid Gland Carcinoma
C0238462|Medullary Carcinoma
C0238462|MTC
C0238462|Medullary thyroid cancer
C0238462|Thyroid cancer, medullary
C0238462|Thyroid carcinoma, medullary
C0238462|Medullary thyroid cancer (MTC)
C0238462|CARCINOMA, C-CELL, MALIGNANT
C0238462|solid carcinoma of the thyroid gland
C0238462|solid carcinoma of thyroid gland
C0238462|medullary thyroid carcinoma (diagnosis)
C0238462|solid carcinoma of the thyroid gland (diagnosis)
C0238462|medullary carcinoma of thyroid gland
C0238462|Medullary Carcinoma of the Thyroid
C0238462|C Cell Carcinoma
C0238462|Medullary Carcinoma of Thyroid
C0238462|Medullary Carcinoma of the Thyroid Gland
C0238462|Thyroid Medullary Carcinoma
C0238462|Parafollicular Cell Carcinoma
C0238462|Ultimobranchial thyroid tumor
C0238462|Ultimobranchial thyroid tumour
C0238462|MTC - Medullary thyroid carcinoma
C0238462|Medullary thyroid carcinoma (disorder)
C0238463|Papillary Thyroid Carcinoma
C0238463|Thyroid Gland Papillary Carcinoma
C0238463|Papillary Thyroid Gland Carcinoma
C0238463|THYROID CARCINOMA, PAPILLARY
C0238463|TPC
C0238463|PTC
C0238463|Thyroid papillary carcinoma
C0238463|PACT
C0238463|Papillary carcinoma of thyroid
C0238463|Papillary thyroid cancer
C0238463|Thyroid cancer, papillary
C0238463|papillary carcinoma of the thyroid gland (diagnosis)
C0238463|papillary carcinoma of the thyroid gland
C0238463|papillary carcinoma of thyroid gland
C0238463|Carcinoma papillary thyroid
C0238463|PTC - Papillary thyroid carcinoma
C0238463|Papillary thyroid carcinoma (disorder)
C0238463|Papillary Cancer of Thyroid Gland
C0238463|Papillary Cancer of Thyroid
C0238463|Papillary Cancer of the Thyroid Gland
C0238463|Papillary Cancer of the Thyroid
C0238463|Papillary Carcinoma of the Thyroid
C1096666|Thyroid cancer metastatic
C2116054|carcinoma simplex of the thyroid gland (diagnosis)
C2116054|carcinoma simplex of thyroid gland
C2116054|carcinoma simplex of the thyroid gland
C2213252|malignant small cell neoplasm of thyroid gland
C2213252|malignant small cell neoplasm of thyroid gland (diagnosis)
C2011415|giant cell type neoplasm of thyroid gland
C2011415|giant cell type neoplasm of thyroid gland (diagnosis)
C2018696|spindle cell type neoplasm of thyroid gland (diagnosis)
C2018696|spindle cell type neoplasm of thyroid gland
C2075656|clear cell type neoplasm of thyroid gland (diagnosis)
C2075656|clear cell type neoplasm of thyroid gland
C0549473|Thyroid Carcinoma
C0549473|Thyroid Gland Carcinoma
C0549473|Thyroid cancer
C0549473|thyroid cancer (diagnosis)
C0549473|Cancers, Thyroid
C0549473|Thyroid Cancers
C0549473|Thyroid Gland Cancer
C0549473|Carcinoma;thyroid gland
C0549473|Cancer, Thyroid
C0549473|Thyroid gland--Cancer
C0549473|Thyroid cancer, NOS
C0549473|carcinoma of thyroid gland
C0549473|thyroid carcinoma (diagnosis)
C0549473|Thyroid Carcinomas
C0549473|Carcinomas, Thyroid
C0549473|Carcinoma thyroid
C0549473|Thyroid carcinoma NOS
C0549473|Cancer of Thyroid
C0549473|Cancer of the Thyroid
C0549473|Head and Neck Cancer, Thyroid
C0549473|Carcinoma of Thyroid
C0549473|Carcinoma of the Thyroid Gland
C0549473|Carcinoma of the Thyroid
C0549473|Carcinoma, Thyroid
C1704228|Thyroid Adenocarcinoma
C1704228|Thyroid Gland Adenocarcinoma
C1704228|Adenocarcinoma of thyroid gland (disorder)
C1704228|Adenocarcinoma of thyroid gland
C1704228|Adenocarcinoma of thyroid
C1704228|thyroid adenocarcinoma (diagnosis)
C1704228|Adenocarcinoma thyroid
C2213264|malignant fibrous histiocytoma of thyroid gland
C2213264|malignant fibrous histiocytoma of thyroid gland (diagnosis)
C1336756|Thyroid Gland Sarcoma
C1336756|Thyroid Sarcoma
C1336756|sarcoma of thyroid gland (diagnosis)
C1336756|sarcoma of thyroid gland
C1336756|Sarcoma of Thyroid
C1336756|Sarcoma of the Thyroid Gland
C1336756|Sarcoma of the Thyroid
C0349668|malignant lymphoma of thyroid gland (diagnosis)
C0349668|malignant lymphoma of thyroid gland
C0349668|Malignant lymphoma of thyroid gland (disorder)
C2213268|malignant plasmacytoma of thyroid gland (diagnosis)
C2213268|malignant plasmacytoma of thyroid gland
C2213270|malignant mastocytosis of thyroid gland (diagnosis)
C2213270|malignant mastocytosis of thyroid gland
C2217675|malignant neoplasm of thyroid gland staging
C2217675|malignant neoplasm of thyroid gland staging (diagnosis)
C2217675|malignant thyroid neoplasm staging
C2217675|malignant tumor of thyroid gland staging
C2217675|thyroid cancer staging
C0347023|Metastatic Malignant Neoplasm to the Thyroid
C0347023|metastasis to thyroid
C0347023|metastasis to thyroid (diagnosis)
C0347023|Metastases to thyroid
C0347023|thyroid malignant neoplasm secondary
C0347023|Secondary malignant neoplasm of thyroid gland
C0347023|Secondary malignant neoplasm of thyroid gland (diagnosis)
C0347023|Metastatic Malignant Neoplasm in the Thyroid Gland
C0347023|Cancer metastatic to thyroid
C0347023|Metastatic malignant neoplasm to thyroid gland
C0347023|Secondary malignant neoplasm of thyroid gland (disorder)
C0347023|Metastasis to the Thyroid Gland
C0347023|Metastasis to the Thyroid
C0347023|Metastatic Malignant Neoplasm to the Thyroid Gland
C0347023|Metastatic Malignant Tumor to the Thyroid Gland
C0347023|Metastatic Malignant Tumor to the Thyroid
C0347023|Metastatic Neoplasm to the Thyroid Gland
C0347023|Metastatic Neoplasm to the Thyroid
C0347023|Metastatic Tumor to the Thyroid Gland
C0347023|Metastatic Tumor to the Thyroid
C0347023|Secondary Malignant Neoplasm to the Thyroid Gland
C0347023|Secondary Malignant Neoplasm to the Thyroid
C0347023|Secondary Malignant Tumor to the Thyroid Gland
C0347023|Secondary Malignant Tumor to the Thyroid
C2062941|differentiated malignant neoplasm of thyroid recurrence after ablation
C2062941|differentiated malignant neoplasm of thyroid recurrence after ablation (diagnosis)
C2062941|malignant thyroid neoplasm recurrence after ablation (differentiated)
C2938921|Thyroid cancer stage 0
C2082467|pleomorphic carcinoma of thyroid gland
C2082467|pleomorphic carcinoma of the thyroid gland
C2082467|pleomorphic carcinoma of the thyroid gland (diagnosis)
C2011267|giant cell carcinoma of thyroid gland
C2011267|giant cell carcinoma of the thyroid gland (diagnosis)
C2011267|giant cell carcinoma of the thyroid gland
C2142937|pseudosarcomatous carcinoma of the thyroid gland (diagnosis)
C2142937|pseudosarcomatous carcinoma of the thyroid gland
C2142937|pseudosarcomatous carcinoma of thyroid gland
C2111819|polygonal cell carcinoma of thyroid gland
C2111819|polygonal cell carcinoma of the thyroid gland (diagnosis)
C2111819|polygonal cell carcinoma of the thyroid gland
C2116055|thyroid carcinoma with osteoclast-like giant cells
C2116055|carcinoma of the thyroid gland with osteoclast-like giant cells (diagnosis)
C2116055|carcinoma of the thyroid gland with osteoclast-like giant cells
C2116055|carcinoma of thyroid gland with osteoclast-like giant cells
C2213254|small cell carcinoma of the thyroid gland (diagnosis)
C2213254|small cell carcinoma of the thyroid gland
C2213254|small cell carcinoma of thyroid gland
C2009891|small cell fusiform cell carcinoma of the thyroid gland
C2009891|fusiform type small cell carcinoma of thyroid gland
C2009891|small cell fusiform cell carcinoma of the thyroid gland (diagnosis)
C2146668|acinar cell carcinoma of thyroid
C2146668|acinar cell carcinoma of the thyroid gland
C2146668|acinar cell carcinoma of the thyroid gland (diagnosis)
C2146668|acinar cell carcinoma of thyroid gland
C1710177|Thyroid Gland Squamous Cell Carcinoma
C1710177|Squamous Cell Thyroid Gland Carcinoma
C1710177|squamous cell carcinoma of thyroid gland
C1710177|squamous cell carcinoma of the thyroid gland (diagnosis)
C1710177|squamous cell carcinoma of the thyroid gland
C2109326|keratinizing squamous cell carcinoma of thyroid gland
C2109326|keratinizing squamous cell carcinoma of the thyroid gland (diagnosis)
C2109326|keratinizing squamous cell carcinoma of the thyroid gland
C2213255|large cell, nonkeratinizing squamous cell carcinoma of the thyroid gland
C2213255|nonkeratinizing large cell squamous carcinoma cell of thyroid gland
C2213255|large cell, nonkeratinizing squamous cell carcinoma of the thyroid gland (diagnosis)
C2213256|small cell, nonkeratinizing squamous cell carcinoma of the thyroid gland (diagnosis)
C2213256|nonkeratinizing small cell squamous cell carcinoma of thyroid gland
C2213256|small cell, nonkeratinizing squamous cell carcinoma of the thyroid gland
C2018573|spindle cell squamous cell carcinoma of the thyroid gland
C2018573|spindle cell squamous cell carcinoma of the thyroid gland (diagnosis)
C2018573|spindle cell squamous cell carcinoma of thyroid gland
C2213257|adenoid squamous cell carcinoma of thyroid gland
C2213257|adenoid squamous cell carcinoma of the thyroid gland (diagnosis)
C2213257|adenoid squamous cell carcinoma of the thyroid gland
C2213258|microinvasive squamous cell carcinoma of the thyroid gland (diagnosis)
C2213258|microinvasive squamous cell carcinoma of thyroid gland
C2213258|microinvasive squamous cell carcinoma of the thyroid gland
C2019459|squamous cell carcinoma with horn formation of thyroid
C2019459|squamous cell carcinoma of the thyroid gland with horn formation (diagnosis)
C2019459|squamous cell carcinoma of the thyroid gland with horn formation
C2019459|squamous cell carcinoma of thyroid gland with horn formation
C1883338|Thyroid Gland Follicular Carcinoma, Minimally Invasive
C1883338|minimally invasive follicular carcinoma of thyroid gland
C1883338|minimally invasive follicular carcinoma of the thyroid gland
C1883338|minimally invasive follicular carcinoma of the thyroid gland (diagnosis)
C2116051|insular carcinoma of the thyroid gland (diagnosis)
C2116051|insular carcinoma of thyroid gland
C2116051|insular carcinoma of the thyroid gland
C0334379|Medullary Carcinoma with Amyloid Stroma
C0334379|Thyroid Gland Medullary Carcinoma with Amyloid Stroma
C0334379|Medullary Thyroid Gland Carcinoma with Amyloid Stroma
C0334379|Medullary carcinoma with amyloid stroma -RETIRED-
C0334379|Medullary carcinoma with amyloid stroma (morphologic abnormality)
C0334379|medullary thyroid carcinoma with amyloid stroma
C0334379|medullary thyroid carcinoma with amyloid stroma (diagnosis)
C0334379|medullary carcinoma of thyroid with amyloid stroma
C0334379|medullary carcinoma of thyroid gland with amyloid stroma
C0334379|carcinoma; medullary with amyloid stroma, unspecified site
C0334379|medullary; carcinoma with amyloid stroma, unspecified site
C0334379|Medullary Adenocarcinoma with Amyloid Stroma
C0334379|Parafollicular Cell Adenocarcinoma with Amyloid Stroma
C0334379|Parafollicular Cell Carcinoma with Amyloid Stroma
C0334379|C Cell Adenocarcinoma with Amyloid Stroma
C0334379|C Cell Carcinoma with Amyloid Stroma
C2116052|mixed medullary-follicular carcinoma of thyroid gland
C2116052|mixed medullary-follicular thyroid carcinoma
C2116052|mixed medullary-follicular thyroid carcinoma (diagnosis)
C1710414|Thyroid Gland Mixed Medullary and Follicular Cell Carcinoma
C1710414|Thyroid Gland Mixed Medullary and Papillary Carcinoma
C1710414|mixed medullary-papillary thyroid carcinoma
C1710414|mixed medullary-papillary carcinoma of thyroid gland
C1710414|mixed medullary-papillary thyroid carcinoma (diagnosis)
C2116053|nonencapsulated sclerosing carcinoma of the thyroid gland
C2116053|nonencapsulated sclerosing carcinoma of thyroid gland
C2116053|nonencapsulated sclerosing carcinoma of the thyroid gland (diagnosis)
C2033139|papillary adenocarcinoma of thyroid gland
C2033139|papillary adenocarcinoma of thyroid gland (diagnosis)
C2116009|adenocarcinoma in villous adenoma of thyroid gland (diagnosis)
C2116009|adenocarcinoma in villous adenoma of thyroid gland
C2116008|adenocarcinoma in tubulovillous adenoma of thyroid gland (diagnosis)
C2116008|adenocarcinoma in tubulovillous adenoma of thyroid gland
C2163817|cystadenocarcinoma of thyroid gland
C2163817|cystadenocarcinoma of the thyroid gland
C2163817|cystadenocarcinoma of the thyroid gland (diagnosis)
C2033251|papillary cystadenocarcinoma of the thyroid gland
C2033251|papillary cystadenocarcinoma of thyroid gland
C2033251|papillary cystadenocarcinoma of the thyroid gland (diagnosis)
C2146680|acinar cell cystadenocarcinoma of thyroid
C2146680|acinar cell cystadenocarcinoma of thyroid gland
C2146680|acinar cell cystadenocarcinoma of the thyroid gland
C2146680|acinar cell cystadenocarcinoma of the thyroid gland (diagnosis)
C3714651|Follicular Variant Papillary Carcinoma
C3714651|Follicular Variant Papillary Thyroid Gland Carcinoma
C3714651|Follicular Variant Thyroid Gland Papillary Carcinoma
C3714651|follicular variant papillary carcinoma of the thyroid gland
C3714651|follicular variant papillary carcinoma of thyroid gland
C3714651|follicular variant papillary carcinoma of the thyroid gland (diagnosis)
C3714651|Follicular Variant Papillary Adenocarcinoma
C3714651|Papillary Carcinoma Follicular Variant
C1709457|Thyroid Gland Papillary Microcarcinoma
C1709457|Papillary Microcarcinoma of the Thyroid Gland
C1709457|Papillary Microcarcinoma of the Thyroid
C1709457|Papillary Thyroid Gland Microcarcinoma
C1709457|Papillary Thyroid Microcarcinoma
C1709457|papillary microcarcinoma of thyroid gland
C1709457|papillary microcarcinoma of the thyroid gland (diagnosis)
C2016175|papillary oxyphilic cell carcinoma of the thyroid gland
C2016175|papillary oxyphilic cell carcinoma of thyroid gland
C2016175|papillary oxyphilic cell carcinoma of the thyroid gland (diagnosis)
C1880498|Encapsulated Thyroid Gland Papillary Carcinoma
C1880498|encapsulated papillary carcinoma of the thyroid gland
C1880498|encapsulated papillary carcinoma of thyroid gland
C1880498|encapsulated papillary carcinoma of the thyroid gland (diagnosis)
C2106521|papillary columnar cell carcinoma of the thyroid gland
C2106521|columnar cell papillary carcinoma of thyroid gland
C2106521|papillary columnar cell carcinoma of the thyroid gland (diagnosis)
C2033239|thyroid malignant carcinoma papillary metastatic to regional lymph node
C2033239|papillary carcinoma of thyroid metastatic to regional lymph node
C2033239|papillary thyroid carcinoma with metastasis to regional lymph nodes (diagnosis)
C2033239|papillary thyroid carcinoma with metastasis to regional lymph nodes
C2033240|thyroid malignant carcinoma papillary metastatic to supraclavicular lymph node
C2033240|papillary thyroid carcinoma with metastasis to supraclavicular lymph nodes
C2033240|papillary thyroid carcinoma with metastasis to supraclavicular lymph nodes (diagnosis)
C2033240|papillary carcinoma of thyroid metastatic to supraclavicular lymph node
C2217676|malignant neoplasm of thyroid stage I
C2217676|malignant neoplasm of thyroid stage I (diagnosis)
C2217676|malignant tumor of thyroid stage I
C2217676|thyroid cancer stage I
C2217677|malignant neoplasm of thyroid stage II
C2217677|malignant neoplasm of thyroid stage II (diagnosis)
C2217677|thyroid cancer stage II
C2217677|malignant tumor of thyroid stage II
C2217678|malignant neoplasm of thyroid stage III
C2217678|malignant neoplasm of thyroid stage III (diagnosis)
C2217678|thyroid cancer stage III
C2217678|malignant tumor of thyroid stage III
C3160834|Thyroid cancer stage IV
C2213253|malignant epithelioma of the thyroid gland
C2213253|malignant epithelioma of thyroid gland
C2213253|malignant epithelioma of the thyroid gland (diagnosis)
C2111684|large cell carcinoma of the thyroid gland (diagnosis)
C2111684|large cell carcinoma of thyroid gland
C2111684|large cell carcinoma of the thyroid gland
C2111754|large cell neuroendocrine carcinoma of thyroid gland
C2111754|large cell neuroendocrine carcinoma of the thyroid gland (diagnosis)
C2111754|large cell neuroendocrine carcinoma of the thyroid gland
C2111685|thyroid malignant carcinoma large cell with rhabdoid phenotype
C2111685|large cell carcinoma of the thyroid gland with rhabdoid phenotype
C2111685|large cell carcinoma of the thyroid gland with rhabdoid phenotype (diagnosis)
C2111685|large cell carcinoma of thyroid gland with rhabdoid phenotype
C2012119|glassy cell carcinoma of thyroid gland
C2012119|glassy cell carcinoma of the thyroid gland (diagnosis)
C2012119|glassy cell carcinoma of the thyroid gland
C2018407|spindle cell carcinoma of thyroid gland
C2018407|spindle cell carcinoma of the thyroid gland (diagnosis)
C2018407|spindle cell carcinoma of the thyroid gland
C2011232|giant cell and spindle cell carcinoma of the thyroid gland
C2011232|giant cell and spindle cell carcinoma of the thyroid gland (diagnosis)
C2011232|giant cell and spindle cell carcinoma of thyroid gland
C2213259|scirrhous adenocarcinoma of thyroid gland (diagnosis)
C2213259|scirrhous adenocarcinoma of thyroid gland
C2037361|superficial spreading adenocarcinoma of thyroid gland (diagnosis)
C2037361|superficial spreading adenocarcinoma of thyroid gland
C2213260|basal cell adenocarcinoma of thyroid gland
C2213260|basal cell adenocarcinoma of thyroid gland (diagnosis)
C2213260|basal cell adenocarcinoma of thyroid
C2145031|trabecular adenocarcinoma of thyroid gland (diagnosis)
C2145031|trabecular adenocarcinoma of thyroid gland
C2189655|villous adenocarcinoma of thyroid gland
C2189655|villous adenocarcinoma of thyroid gland (diagnosis)
C2016174|oxyphilic adenocarcinoma of thyroid gland
C2016174|oxyphilic adenocarcinoma of thyroid gland (diagnosis)
C2075544|clear cell adenocarcinoma of thyroid gland
C2075544|clear cell adenocarcinoma of thyroid gland (diagnosis)
C2116005|alveolar adenocarcinoma of thyroid gland (diagnosis)
C2116005|alveolar adenocarcinoma of thyroid gland
C2203046|well differentiated follicular adenocarcinoma of thyroid gland (diagnosis)
C2203046|well differentiated follicular adenocarcinoma of thyroid gland
C2213261|follicular trabecular adenocarcinoma of thyroid gland (diagnosis)
C2213261|follicular trabecular adenocarcinoma of thyroid gland
C2116050|fetal adenocarcinoma of thyroid gland
C2116050|fetal adenocarcinoma of thyroid gland (diagnosis)
C2213262|embryonal carcinosarcoma of thyroid gland (diagnosis)
C2213262|embryonal carcinosarcoma of thyroid gland
C2213263|malignant myoepithelioma of thyroid gland
C2213263|malignant myoepithelioma of thyroid gland (diagnosis)
C2046351|histiocytic sarcoma of thyroid gland (diagnosis)
C2046351|histiocytic sarcoma of thyroid gland
C2111188|Langerhans cell sarcoma of thyroid gland (diagnosis)
C2111188|Langerhans cell sarcoma of thyroid gland
C2077774|interdigitating dendritic cell sarcoma of thyroid gland (diagnosis)
C2077774|interdigitating dendritic cell sarcoma of thyroid gland
C2213266|follicular dendritic cell sarcoma of thyroid gland (diagnosis)
C2213266|follicular dendritic cell sarcoma of thyroid gland
C2033237|thyroid malignant carcinoma papillary metastatic to cervical lymph node
C2033237|papillary thyroid carcinoma with metastasis to cervical lymph nodes (diagnosis)
C2033237|papillary thyroid carcinoma with metastasis to cervical lymph nodes
C2033237|papillary carcinoma of thyroid metastatic to cervical lymph node
C3163939|Carcinoma of thyroid
C3163939|Malignant epithelial neoplasm of thyroid
C3163939|Malignant epithelial neoplasm of thyroid (disorder)
C2116063|malignant histiocytosis of thyroid gland (diagnosis)
C2116063|malignant histiocytosis of thyroid gland
C2098465|thyroid biopsy showing malignant neoplasm
C2098465|thyroid biopsy malignant neoplasm (procedure)
C2098465|thyroid biopsy malignant neoplasm
C0278861|Recurrent Thyroid Carcinoma
C0278861|Recurrent Thyroid Gland Carcinoma
C0278861|Thyroid cancer recurrent
C0278861|recurrent thyroid cancer
C0278861|thyroid cancer, recurrent
C0278861|Recurrent Cancer of Thyroid Gland
C0278861|Recurrent Cancer of Thyroid
C0278861|Recurrent Cancer of the Thyroid Gland
C0278861|Recurrent Cancer of the Thyroid
C0278861|Relapsed Cancer of Thyroid Gland
C0278861|Relapsed Cancer of Thyroid
C0278861|Relapsed Cancer of the Thyroid Gland
C0278861|Relapsed Cancer of the Thyroid
C0278861|Relapsed Thyroid Cancer
C0278861|Relapsed Thyroid Gland Cancer
C0205642|Adenocarcinomas, Oxyphilic
C0205642|Oxyphilic Adenocarcinomas
C0205642|Oxyphilic Adenocarcinoma
C0205642|oxyphilic adenocarcinoma (diagnosis)
C0205642|Oxyphilic adenocarcinoma (disorder)
C0205642|Huerthle cell carcinoma
C0205642|ONCOCYTOMA, MALIGNANT
C0205642|Hurthle Cell Adenocarcinoma
C0205642|Oncocytic Adenocarcinoma
C0205642|Oncocytic Carcinoma
C0205642|Hurthle Cell Carcinoma
C0205642|Follicular carcinoma, oxyphilic cell
C0205642|Oxyphilic adenocarcinoma (morphologic abnormality)
C0205642|Hurthle cell; adenocarcinoma
C0205642|Hurthle cell; carcinoma
C0205642|carcinoma; Hurthle cell
C0205642|adenocarcinoma; Hurthle cell
C0205642|Adenocarcinoma, Oxyphilic
C1306310|Primary malignant neoplasm of thyroid gland (diagnosis)
C1306310|Primary malignant neoplasm of thyroid gland
C1306310|thyroid malignant neoplasm primary
C1306310|Primary malignant neoplasm of thyroid gland (disorder)
C1282509|metastasis from malignant neoplasm of thyroid
C1282509|metastasis from malignant neoplasm of thyroid (diagnosis)
C1282509|Metastasis from malignant tumor of thyroid (disorder)
C1282509|Metastasis from malignant tumor of thyroid
C1282509|Metastasis from malignant tumour of thyroid
C1282469|local recurrence of malignant neoplasm of thyroid gland
C1282469|thyroid malignant neoplasm local recurrence
C1282469|local recurrence of malignant neoplasm of thyroid gland (diagnosis)
C1282469|Local recurrence of malignant tumor of thyroid gland (disorder)
C1282469|Local recurrence of malignant tumor of thyroid gland
C1282469|Local recurrence of malignant tumour of thyroid gland
C4038608|Diffuse sclerosing papillary thyroid carcinoma (disorder)
C4038608|Diffuse sclerosing papillary thyroid carcinoma
C1266050|Poorly Differentiated Thyroid Carcinoma
C1266050|Thyroid Gland Poorly Differentiated Carcinoma
C1266050|Poorly Differentiated Thyroid Gland Carcinoma
C1266050|Insular carcinoma (morphologic abnormality)
C1266050|Insular carcinoma
C1266050|Poorly Differentiated Carcinoma of Thyroid Gland
C1266050|Poorly Differentiated Carcinoma of the Thyroid Gland
C0206683|Carcinoma, Papillary, Follicular
C0206683|Thyroid Gland Papillary and Follicular Carcinoma
C0206683|Carcinoma, Papillary, Follicular [Disease/Finding]
C0206683|Papillary and Follicular Adenocarcinoma
C0206683|Papillary and Follicular Carcinoma
C0206683|Follicular Variant Thyroid Gland Papillary Carcinoma
C0206683|Papillary adenocarcinoma - follicular variant
C0206683|Papillary adenocarcinoma, follicular variant
C0206683|Papillary carcinoma - follicular variant
C0206683|Papillary carcinoma, follicular variant
C0206683|Papillary and follicular adenocarcinoma (morphologic abnormality)
C0206683|Papillary carcinoma, follicular variant (morphologic abnormality)
C0206683|carcinoma; follicular with papillary
C0206683|carcinoma; papillary with follicular
C0206683|carcinoma; papillary, follicular variant
C0206683|follicular; adenocarcinoma with papillary
C0206683|follicular; carcinoma, with papillary
C0206683|adenocarcinoma; follicular with papillary
C0206683|adenocarcinoma; papillary with follicular
C0206683|adenocarcinoma; papillary, follicular variant
C0206683|papillary; adenocarcinoma with follicular
C0206683|papillary; adenocarcinoma, follicular variant
C0206683|papillary; carcinoma, follicular variant
C0206683|papillary; carcinoma, with follicular
C1386262|follicular; adenocarcinoma, intermediate differentiation
C1386262|adenocarcinoma; follicular, intermediate differentiation
C1386263|follicular; adenocarcinoma, unspecified site
C1386263|adenocarcinoma; follicular, unspecified site
C0334327|Follicular adenocarcinoma - moderately differentiated
C0334327|Follicular adenocarcinoma - trabecular
C0334327|Follicular adenocarcinoma, moderately differentiated
C0334327|Follicular adenocarcinoma, trabecular
C0334327|Follicular carcinoma - moderately differentiated
C0334327|Follicular carcinoma - trabecular
C0334327|Follicular carcinoma, moderately differentiated
C0334327|Follicular carcinoma, trabecular
C0334327|Follicular adenocarcinoma, trabecular (morphologic abnormality)
C0334327|carcinoma; follicular, trabecular
C0334327|carcinoma; trabecular, follicular
C0334327|Langhans; wuchernde Struma
C0334327|follicular; adenocarcinoma, trabecular
C0334327|follicular; carcinoma, trabecular
C0334327|adenocarcinoma; follicular, trabecular
C0334327|adenocarcinoma; trabecular follicular
C0334327|trabecular; follicular adenocarcinoma
C0334327|wuchernde Struma Langhans
C0334327|Trabecular Follicular Adenocarcinoma
C0334330|Nonencapsulated sclerosing adenocarcinoma
C0334330|Nonencapsulated sclerosing carcinoma
C0334330|Nonencapsulated sclerosing carcinoma (morphologic abnormality)
C0334330|Papillary carcinoma, diffuse sclerosing
C0334330|carcinoma; nonencapsulated sclerosing
C0334330|adenocarcinoma; nonencapsulated sclerosing
C0334330|nonencapsulated sclerosing; carcinoma
C0334330|nonencapsulated; sclerosing adenocarcinoma
C0334330|Nonencapsulated Sclerosing Neoplasm
C1541839|carcinoma; C-cell, unspecified site
C1541839|C-cell; carcinoma, unspecified site
C1391909|carcinoma; follicular, intermediate differentiation
C1391909|follicular; carcinoma, intermediate differentiation
C1391910|carcinoma; follicular, unspecified site
C1391910|follicular; carcinoma, unspecified site
C1391938|carcinoma; parafollicular cell, unspecified site
C1391938|parafollicular cell; carcinoma, unspecified site
C1397650|follicular; carcinoma, pure follicle
C1399823|Hurthle cell; tumor, malignant
C1399823|tumor; Hurthle cell, malignant
C1321862|Nonencapsulated Sclerosing Papillary Thyroid Carcinoma
C1321862|Thyroid Gland Diffuse Sclerosing Papillary Carcinoma
C1321862|Nonencapsulated sclerosing tumor
C1321862|Nonencapsulated sclerosing tumour
C1321862|nonencapsulated; sclerosing tumor
C1321862|tumor; nonencapsulated sclerosing
C1410366|struma; toxic, tumor, malignant
C1410366|toxic; goiter, tumor, malignant
C1522358|Mouse Thyroid Carcinoma
C0280258|stage/cell type, thyroid cancer
C0280258|thyroid cancer stage
C1336753|Thyroid Gland Lymphoma
C1336753|Thyroid Lymphoma
C1336753|Primary Thyroid Gland Lymphoma
C1336753|Lymphoma of Thyroid Gland
C1336753|Lymphoma of Thyroid
C1336753|Lymphoma of the Thyroid Gland
C1336753|Lymphoma of the Thyroid
C0686505|Malignant neoplasm of thyroglossal duct
C0686505|Primary malignant neoplasm of thyroglossal duct
C0686505|thyroid neoplasm location: ectopic thyroglossal duct malignant primary
C0686505|Primary malignant neoplasm of thyroglossal duct (diagnosis)
C0686505|Primary malignant neoplasm of thyroglossal duct (disorder)
C1302463|pT4b: Extrathyroidal anaplastic carcinoma - surgically unresectable (anaplastic carcinoma) (thyroid) (finding)
C1302463|pT4b: Extrathyroidal anaplastic carcinoma - surgically unresectable (anaplastic carcinoma) (thyroid)
C1276616|T2: Tumor > 1 cm but < 4 cm, limited to thyroid (finding)
C1276616|T2: Tumor > 1 cm but < 4 cm, limited to thyroid
C1276616|T2: Tumour > 1 cm but < 4 cm, limited to thyroid
C1276616|T2: Tumor > 1 cm but < 4 cm, limited to thyroid (tumor staging)
C1276617|T3: Thyroid tumor > 4 cm, limited to thyroid (finding)
C1276617|T3: Thyroid tumor > 4 cm, limited to thyroid
C1276617|T3: Thyroid tumour > 4 cm, limited to thyroid
C1276617|T3: Thyroid tumor > 4 cm, limited to thyroid (tumor staging)
C1276618|T4: Thyroid tumor of any size extending beyond the thyroid capsule (finding)
C1276618|T4: Thyroid tumor of any size extending beyond the thyroid capsule
C1276618|T4: Thyroid tumour of any size extending beyond the thyroid capsule
C1276618|T4: Thyroid tumor of any size extending beyond the thyroid capsule (tumor staging)
C0346398|Mixed follicular and papillary thyroid carcinoma
C0346398|thyroid malignant carcinoma mixed follicular and papillary
C0346398|Mixed follicular and papillary thyroid carcinoma (diagnosis)
C0346398|Mixed follicular and papillary thyroid carcinoma (disorder)
C0749424|Thyroid Hurthle Cell Carcinoma
C0749424|Thyroid Gland Oncocytic Follicular Carcinoma
C0749424|Hurthle Cell Thyroid Gland Carcinoma
C0749424|Hurthle cell carcinoma of thyroid
C0749424|Hurthle cell carcinoma of thyroid (disorder)
C0749424|THYROID CARCINOMA, HURTHLE CELL
C0749424|Thyroid cancer, follicular, Hurthle cell type
C0749424|Follicular thyroid cancer, Hurthle cell type
C0749424|Hurthle cell carcinoma of the thyroid
C0749424|Thyroid cancer, Hurthle cell
C0749424|Hurthle cell carcinoma of thyroid (diagnosis)
C0749424|thyroid malignant carcinoma hurthle cell
C0749424|Hurthle Cell Thyroid Neoplasia
C0749424|Cancer of thyroid, Hurthle cell
C0749424|Hurthle cell neoplasm of the thyroid
C0749424|Hurthle Cell Carcinoma of Thyroid Gland
C0749424|Hurthle Cell Carcinoma of the Thyroid Gland
C0749424|Oncocytic Carcinoma of Thyroid
C0749424|Oncocytic Carcinoma of the Thyroid
C0749424|Thyroid Gland Hurthle Cell Carcinoma
C0749424|Thyroid Oncocytic Carcinoma
C1302519|pT4a: Intrathyroidal anaplastic carcinoma - surgically resectable (anaplastic carcinoma) (thyroid) (finding)
C1302519|pT4a: Intrathyroidal anaplastic carcinoma - surgically resectable (anaplastic carcinoma) (thyroid)
C2213271|Sezary syndrome of thyroid gland (diagnosis)
C2213271|Sezary syndrome of thyroid gland
C2113733|precursor cell lymphoblastic lymphoma of thyroid gland (diagnosis)
C2113733|precursor cell lymphoblastic lymphoma of thyroid gland
C2213265|mast cell sarcoma of thyroid gland
C2213265|mast cell sarcoma of thyroid gland (diagnosis)
C0346643|Malignant neoplasm of hepatic duct
C0346643|malignant extrahepatic neoplasm hepatic duct
C0346643|malignant neoplasm of hepatic duct (diagnosis)
C0346643|Malignant neoplasm of hepatic duct (disorder)
C0546835|Malignant neoplasm of intrahepatic biliary passages
C0546835|Malignant neoplasm of intrahepatic bile ducts
C0546835|malignant neoplasm of intrahepatic bile duct (diagnosis)
C0546835|malignant neoplasm of intrahepatic bile duct
C0546835|malignant tumor of intrahepatic bile duct
C0546835|Mal neo intrahepat ducts
C0546835|Ca intrahepatic bile ducts
C0546835|Malignant neoplasm of intrahepatic bile ducts NOS (disorder)
C0546835|Ca intrahepatic bile ducts (disorder)
C0546835|Malignant neoplasm of intrahepatic bile ducts NOS
C0546835|Malignant neoplasm of intrahepatic biliary passages (disorder)
C0546835|Malignant neoplasm of intrahepatic bile ducts (disorder)
C0546835|Intrahepatic bile duct cancer
C0546835|Intrahepatic bile duct cancer NOS
C0546835|Malignant neoplasm of intrahepatic gall duct
C0546835|Malignant neoplasm of intrahepatic gall duct (disorder)
C2239176|Liver cell carcinoma
C2239176|Carcinoma, Hepatocellular
C2239176|Carcinomas, Hepatocellular
C2239176|Hepatocellular Carcinomas
C2239176|Hepatoma
C2239176|Hepatomas
C2239176|hepatocellular carcinoma
C2239176|LCC
C2239176|carcinoma of liver (diagnosis)
C2239176|hepatocellular carcinoma of liver (diagnosis)
C2239176|hepatocellular carcinoma of liver
C2239176|liver neoplasm malignant carcinoma
C2239176|carcinoma of liver
C2239176|Liver carcinoma
C2239176|Liver Cell Cancer (Hepatocellular Carcinoma)
C2239176|Carcinoma, Hepatocellular [Disease/Finding]
C2239176|Cancers, Adult Liver
C2239176|Adult Liver Cancer
C2239176|Cancer, Adult Liver
C2239176|Adult Liver Cancers
C2239176|Liver Cancers, Adult
C2239176|Liver Cancer, Adult
C2239176|Liver Cell Carcinoma, Adult
C2239176|Liver Cell Carcinomas
C2239176|Cell Carcinoma, Liver
C2239176|Cell Carcinomas, Liver
C2239176|Carcinoma, Liver Cell
C2239176|Carcinomas, Liver Cell
C2239176|Hepatic cell carcinoma
C2239176|Primary carcinoma of liver
C2239176|liver neoplasm malignant carcinoma primary
C2239176|Primary carcinoma of liver (diagnosis)
C2239176|HCC
C2239176|CARCINOMA, HEPATOCELLULAR, MALIGNANT
C2239176|[M]Hepatocellular carcinoma NOS
C2239176|Carcinoma of the Liver Cells
C2239176|Primary Carcinoma of the Liver Cells
C2239176|Carcinoma of Liver Cells
C2239176|Primary Carcinoma of Liver Cells
C2239176|Liver cell carcinoma (clinical)
C2239176|Hepatocellular carcinoma (clinical)
C2239176|Carcinoma liver
C2239176|Carcinoma hepatocellular
C2239176|Hepatocarcinoma
C2239176|Hepatoma, malignant
C2239176|Malignant hepatoma
C2239176|LCC - Liver cell carcinoma
C2239176|HCC - Hepatocellular carcinoma
C2239176|Hepatocellular carcinoma (morphologic abnormality)
C2239176|Liver cell carcinoma (disorder)
C2239176|Primary carcinoma of liver (disorder)
C2239176|carcinoma; hepatic cell
C2239176|carcinoma; hepatocellular
C2239176|hepatic cell; carcinoma
C2239176|hepatocellular; carcinoma
C2239176|Hepatocellular carcinoma, NOS
C2239176|Hepatoma, NOS
C2239176|Carcinoma of liver, specified as primary
C2239176|Carcinoma of liver cell
C0206624|Hepatoblastoma
C0206624|Hepatoblastomas
C0206624|hepatoblastoma of liver
C0206624|hepatoblastoma of liver (diagnosis)
C0206624|Hepatoblastoma [Disease/Finding]
C0206624|HBL
C0206624|HEPATOBLASTOMA, MALIGNANT
C0206624|Pediatric Hepatoblastoma
C0206624|Pediatric Embryonal Hepatoma
C0206624|Hepatoblastoma NOS
C0206624|Embryonal hepatoma
C0206624|HBL - Hepatoblastoma
C0206624|Hepatoblastoma (clinical)
C0206624|Hepatoblastoma (disorder)
C0206624|Hepatoblastoma (morphologic abnormality)
C0206624|childhood hepatoblastoma
C0206624|hepatoblastoma, childhood
C0206624|embryonal; hepatoma
C0206624|hepatoma; embryonal
C0345907|Angiosarcoma of liver
C0345907|Hepatic angiosarcoma
C0345907|hemangiosarcoma of liver
C0345907|hemangiosarcoma of liver (diagnosis)
C0345907|hepatic hemangiosarcoma
C0345907|Liver Angiosarcoma
C0345907|Angiosarcoma of liver (disorder)
C0345907|Hemangiosarcoma of liver (disorder)
C0345907|liver neoplasm malignant angiosarcoma
C0345907|Angiosarcoma of liver (diagnosis)
C0345907|Primary angiosarcoma of liver
C0345907|liver; angiosarcoma
C0345907|angiosarcoma; liver
C0345907|Hemangiosarcoma of the Liver
C0345907|Liver Hemangiosarcoma
C0345907|Angiosarcoma of the Liver
C0345907|Primary Angiosarcoma of the Liver
C0345905|Intrahepatic bile duct carcinoma
C0345905|cholangiocarcinoma of intrahepatic bile duct (diagnosis)
C0345905|cholangiocarcinoma of intrahepatic bile duct
C0345905|carcinoma of intrahepatic bile duct
C0345905|carcinoma of intrahepatic bile duct (diagnosis)
C0345905|CHOLANGIOCARCINOMA, INTRAHEPATIC, MALIGNANT
C0345905|Intrahepatic Carcinoma of the Bile Duct
C0345905|Intrahepatic Carcinoma of Bile Duct
C0345905|Cholangiocarcinomas, Intrahepatic
C0345905|Intrahepatic Cholangiocarcinomas
C0345905|Cholangiocarcinoma, Intrahepatic
C0345905|Intrahepatic cholangiocarcinoma
C0345905|Intrahepatic bile duct carcinoma (disorder)
C0345905|ICC
C0345905|Intrahepatic Cholangiocellular Carcinoma
C0348340|Other specified carcinomas of liver
C0348340|[X]Other specified carcinomas of liver
C0348340|Other specified carcinoma of liver
C0348340|Other specified carcinoma of liver (disorder)
C0348340|[X]Other specified carcinomas of liver (disorder)
C0345904|Liver, unspecified
C0345904|Malignant neoplasm of liver, unspecified
C0345904|malignant neoplasm of liver
C0345904|liver cancer
C0345904|liver cancer (diagnosis)
C0345904|liver neoplasm malignant
C0345904|malignant neoplasm of liver (diagnosis)
C0345904|Hepatic neoplasms malignant
C0345904|Cancer, Hepatic
C0345904|Cancers, Hepatic
C0345904|Hepatic Cancers
C0345904|Cancers, Liver
C0345904|Liver Cancers
C0345904|malignant tumor of liver
C0345904|Malignant neo liver NOS
C0345904|Malignant neoplasm of liver, not specified as primary or secondary
C0345904|hepatic cancer
C0345904|Cancer, Liver
C0345904|Malig neoplasm of liver, not specified as primary or sec
C0345904|Cancers, Hepatocellular
C0345904|Hepatocellular Cancers
C0345904|Malignant neoplasm of liver unspecified (disorder)
C0345904|Malignant tumor of liver (disorder)
C0345904|Malignant neoplasm of liver unspecified
C0345904|Malignant tumour of liver
C0345904|Liver--Cancer
C0345904|CANCER, HEPATOCELLULAR
C0345904|Hepatic neoplasm malignant NOS
C0345904|Malignant hepatic neoplasm
C0345904|Malignant liver tumor
C0345904|Hepatic tumour malignant
C0345904|Liver, cancer of
C0345904|Malignant liver tumour
C0345904|Hepatic neoplasm malignant
C0345904|Hepatic tumor malignant
C0345904|Hepatocellular Cancer
C0345904|Cancer of the Liver
C0345904|CA - Liver cancer
C0345904|Malignant neoplasm of liver (disorder)
C0345904|Malignant neoplasm of liver, NOS
C0345904|Cancer of Liver
C0345904|Neoplasm malig;liver
C0345904|malignant neosplasm of the liver
C0348339|Other sarcomas of liver
C0348339|Other sarcoma of liver
C0348339|[X]Other sarcomas of the liver (disorder)
C0348339|[X]Other sarcomas of the liver
C0348339|Other sarcoma of liver (disorder)
C0153448|Malignant neoplasm of liver and intrahepatic bile ducts
C0153448|Cancer of liver and intrahepatic bile duct
C0153448|Malignant neoplasm of liver and intrahepatic bile ducts NOS
C0153448|Malignant neoplasm of liver and intrahepatic bile ducts NOS (disorder)
C0153448|malignant neoplasm of liver and intrahepatic bile ducts (diagnosis)
C0153448|Malignant neoplasm of liver and intrahepatic bile ducts (disorder)
C2837938|Malignant neoplasm of liver, primary, unspecified as to type
C2188066|undifferentiated carcinoma of intrahepatic bile duct
C2188066|undifferentiated carcinoma of intrahepatic bile duct (diagnosis)
C2078126|undifferentiated sarcoma of intrahepatic bile duct (diagnosis)
C2078126|undifferentiated sarcoma of intrahepatic bile duct
C0279000|Liver and Intrahepatic Bile Duct Carcinoma
C0279000|Liver and Intrahepatic Biliary Tract Carcinoma
C0279000|Liver and hepatobiliary cancer, NOS
C0279000|Liver/hepatobiliary cancer
C0279000|liver cancer
C0279000|liver and intrahepatic biliary tract cancer
C0279000|Hepatic Cancer
C0279000|Cancer of Liver
C0279000|Cancer of the Liver
C0279000|Liver and Intrahepatic Bile Duct Cancer
C0279000|Primary Liver Carcinoma
C0279000|Cancer of Liver and Intrahepatic Biliary Tract
C0279000|Cancer of the Liver and Intrahepatic Biliary Tract
C0024620|Primary liver cancer
C0024620|Primary malignant neoplasm of liver
C0024620|Mal neo liver, primary
C0024620|Primary Malignant Liver Neoplasm
C0024620|primary malignant neoplasm of liver (diagnosis)
C0024620|liver neoplasm malignant primary
C0024620|Ca liver - primary (disorder)
C0024620|Primary malignant neoplasm of liver NOS (disorder)
C0024620|Primary malignant neoplasm of liver (disorder)
C0024620|Ca liver - primary
C0024620|Primary malignant neoplasm of liver NOS
C0024620|Malignant neoplasm of liver, primary
C0024620|Liver, cancer of, primary
C0024620|Primary cancer of liver
C0024620|Cancer of liver, primary
C0206630|Sarcoma, Endometrial Stromal
C0206630|Endometrial Stromal Sarcomas
C0206630|Sarcomas, Endometrial Stromal
C0206630|Stromal Sarcoma, Endometrial
C0206630|Stromal Sarcomas, Endometrial
C0206630|Sarcoma, Endometrial Stromal [Disease/Finding]
C0206630|Endometrial Stromal Sarcoma
C0206630|Endometrioid Stromal Sarcoma
C0206630|Endometrial stromal sarcoma (disorder)
C0206630|STROMAL SARCOMA, ENDOMETRIAL, MALIGNANT
C0206630|ESS
C0206630|Primary malignant stromal sarcoma of endometrium
C0206630|Endometrial sarcoma
C0206630|Endometrial sarcoma, NOS
C0206630|Stromal sarcoma, NOS
C0346191|Endometrium
C0346191|Carcinoma in situ of endometrium
C0346191|Ca endometrium stage 0
C0346191|Endometrial cancer stage 0
C0346191|Carcinoma in situ of endometrium (disorder)
C0346191|Cancer of endometrium stage 0
C0346191|Endometrial carcinoma stage 0
C0346191|Carcinoma endometrial stage 0
C0346191|stage 0 endometrial cancer
C0346191|cancer of the endometrium, stage 0
C0346191|carcinoma of the endometrium, stage 0
C0346191|endometrial cancer, stage 0
C0346191|endometrial carcinoma, stage 0
C0346191|stage 0 cancer of the endometrium
C0346191|stage 0 carcinoma of the endometrium
C0346191|stage 0 uterine cancer
C0346191|uterine cancer, stage 0
C0476089|CARCINOMA OF ENDOMETRIUM
C0476089|Cancer, Endometrial
C0476089|Cancers, Endometrial
C0476089|Endometrial Cancers
C0476089|ENDOMETRIAL CANCER
C0476089|Ca endometrium
C0476089|Endometrial carcinoma (NOS)
C0476089|Cancers, Endometrium
C0476089|Endometrium Cancers
C0476089|Cancer, Endometrium
C0476089|Endometrial carcinoma
C0476089|Endometrial Ca
C0476089|uterine neoplasm, malignant - of endometrium carcinoma
C0476089|Endometrial carcinoma (diagnosis)
C0476089|Carcinoma, Endometrial
C0476089|Carcinomas, Endometrial
C0476089|Endometrial Carcinomas
C0476089|Endometrium Carcinoma
C0476089|Endometrium Carcinomas
C0476089|Endometrium--Cancer
C0476089|CARCINOMA, ENDOMETRIAL, MALIGNANT
C0476089|Carcinoma of the Endometrium
C0476089|Cancer of endometrium
C0476089|Carcinoma endometrial
C0476089|Endometrial cancer NOS
C0476089|Endometrium Cancer
C0476089|Cancer of the Endometrium
C0476089|Endometrial carcinoma (disorder)
C0476089|Carcinoma;endometrial
C0813216|Corpus uteri carcinoma
C0813216|Carcinoma of corpus uteri
C0813216|Malignant epithelial neoplasm of body of uterus (disorder)
C0813216|Malignant epithelial neoplasm of body of uterus
C0813216|Carcinoma body of uterus
C0813216|uterine neoplasm, malignant - of corpus uteri carcinoma
C0813216|Carcinoma of corpus uteri (diagnosis)
C0813216|Carcinoma corpus uteri
C1153706|Uterine adenocarcinoma
C1153706|adenocarcinoma of uterus
C1153706|adenocarcinoma of uterus (diagnosis)
C1153706|Endometrial adenocarcinoma
C1153706|[M]Endometrioid adenomas and carcinomas
C1153706|[M]Endometrioid adenomas and carcinomas (morphologic abnormality)
C1153706|[M]Endometrioid adenoma or carcinoma NOS (morphologic abnormality)
C1153706|[M]Endometrioid adenoma or carcinoma NOS
C1153706|ADENOCARCINOMA, ENDOMETRIAL, MALIGNANT
C1153706|Adenocarcinoma of endometrium (diagnosis)
C1153706|Adenocarcinoma of endometrium
C1153706|uterine adenocarcinoma endometrium
C1153706|Adenocarcinoma of the Endometrium
C1153706|Adenocarcinoma endometrial
C1153706|Adenocarcinoma of endometrium (disorder)
C1153706|Adenocarcinoma of uterus (disorder)
C1153706|adenocarcinoma of the uterus
C1153706|uterine cancer, adenocarcinoma
C1153706|uterus cancer, adenocarcinoma
C0153574|Corpus uteri, unspecified
C0153574|Malignant neoplasm of corpus uteri
C0153574|Malignant neoplasm of corpus uteri, unspecified
C0153574|Malignant neoplasm of body of uterus
C0153574|malignant neoplasm of corpus uteri (diagnosis)
C0153574|malignant tumor of corpus uteri
C0153574|Malignant neoplasm of corpus uteri NOS
C0153574|Malignant tumor of body of uterus
C0153574|Body of uterus Ca
C0153574|Malignant neoplasm of body of uterus NOS
C0153574|Uterus body Ca
C0153574|Malignant neoplasm of corpus uteri NOS (disorder)
C0153574|Malignant tumour of body of uterus
C0153574|Malignant tumour of body of uterus (disorder)
C0153574|Malignant neoplasm of body of uterus NOS (disorder)
C0153574|Cancer of uterine body
C0153574|Uterine cancer, body
C0153574|Cancer of body of uterus
C0153574|Malignant neoplasm of body of uterus (disorder)
C0153574|uterine corpus cancer
C0153574|Malignant Corpus Uteri Neoplasm
C0153574|Malignant Corpus Uteri Tumor
C0153574|Malignant Neoplasm of Uterine Body
C0153574|Malignant Neoplasm of the Uterine Body
C0153574|Malignant Tumor of Uterine Body
C0153574|Malignant Tumor of the Uterine Body
C0153574|Malignant Uterine Body Neoplasm
C0153574|Malignant Uterine Body Tumor
C0153574|Malignant Uterine Corpus Neoplasm
C0153574|Malignant Uterine Corpus Tumor
C0338113|sarcoma of uterus (diagnosis)
C0338113|sarcoma of uterus
C0338113|uterine sarcoma
C0338113|Sarcoma uterus
C0338113|Uterine sarcoma NOS
C0338113|Sarcoma of uterus (disorder)
C0338113|sarcoma of the uterus
C0338113|uterine cancer, sarcoma
C0338113|uterine corpus cancer, sarcoma
C0338113|uterus cancer, sarcoma
C0338113|Corpus Uteri Sarcoma
C0338113|Sarcoma of Body of Uterus
C0338113|Sarcoma of Corpus Uteri
C0338113|Sarcoma of Uterine Body
C0338113|Sarcoma of Uterine Corpus
C0338113|Sarcoma of the Body of Uterus
C0338113|Sarcoma of the Corpus Uteri
C0338113|Sarcoma of the Uterine Body
C0338113|Sarcoma of the Uterine Corpus
C0338113|Uterine Body Sarcoma
C0338113|Uterine Corpus Sarcoma
C0338113|Uterus Sarcoma
C0338113|Body of Uterus Sarcoma
C1297960|uterine neoplasm, malignant corpus uteri, by direct extension from bladder
C1297960|malignant neoplasm involving uterine corpus by direct extension from bladder (diagnosis)
C1297960|malignant neoplasm involving uterine corpus by direct extension from bladder
C1297960|Malignant tumor involving uterine corpus by direct extension from bladder (disorder)
C1297960|Malignant tumor involving uterine corpus by direct extension from bladder
C1297960|Malignant tumour involving uterine corpus by direct extension from bladder
C1297961|malignant neoplasm involving uterine corpus by direct extension from ovary (diagnosis)
C1297961|uterine neoplasm, malignant corpus uteri, by direct extension from ovary
C1297961|malignant neoplasm involving uterine corpus by direct extension from ovary
C1297961|Malignant tumor involving uterine corpus by direct extension from ovary (disorder)
C1297961|Malignant tumor involving uterine corpus by direct extension from ovary
C1297961|Malignant tumour involving uterine corpus by direct extension from ovary
C1297962|malignant neoplasm involving uterine corpus by direct extension from uterine cervix
C1297962|malignant neoplasm involving uterine corpus by direct extension from uterine cervix (diagnosis)
C1297962|uterine neoplasm, malignant corpus uteri by direct extension from uterine cervix
C1297962|Malignant tumor involving uterine corpus by direct extension from uterine cervix (disorder)
C1297962|Malignant tumor involving uterine corpus by direct extension from uterine cervix
C1297962|Malignant tumour involving uterine corpus by direct extension from uterine cervix
C1297963|uterine neoplasm, malignant corpus uteri, by direct extension from vagina
C1297963|malignant neoplasm involving uterine corpus by direct extension from vagina (diagnosis)
C1297963|malignant neoplasm involving uterine corpus by direct extension from vagina
C1297963|Malignant tumor involving uterine corpus by direct extension from vagina (disorder)
C1297963|Malignant tumor involving uterine corpus by direct extension from vagina
C1297963|Malignant tumour involving uterine corpus by direct extension from vagina
C1298046|uterine neoplasm, malignant corpus uteri by direct extension from fallopian tube
C1298046|malignant neoplasm involving uterine corpus by direct extension from fallopian tube (diagnosis)
C1298046|malignant neoplasm involving uterine corpus by direct extension from fallopian tube
C1298046|Malignant tumor involving uterine corpus by direct extension from fallopian tube (disorder)
C1298046|Malignant tumor involving uterine corpus by direct extension from fallopian tube
C1298046|Malignant tumour involving uterine corpus by direct extension from fallopian tube
C0153567|uterine cancer
C0153567|Malignant neoplasm of uterus, part unspecified
C0153567|malignant neoplasm of uterus (diagnosis)
C0153567|cancer of uterus
C0153567|malignant neoplasm of uterus
C0153567|uterine cancer (diagnosis)
C0153567|Cancer, Uterine
C0153567|Cancers, Uterine
C0153567|Uterine Cancers
C0153567|Cancers, Uterus
C0153567|Uterus Cancers
C0153567|malignant tumor of uterus
C0153567|Malig neopl uterus NOS
C0153567|Cancer, Uterus
C0153567|Malignant neoplasm of uterus, part unspecified (disorder)
C0153567|Malignant neoplasm of uterus (disorder)
C0153567|CA - Cancer of uterus
C0153567|Malignant tumour of uterus
C0153567|Uterine Ca NOS
C0153567|Ca uterus NOS
C0153567|Uterus--Cancer
C0153567|Uterine cancer, NOS
C0153567|-- Uterine Cancer
C0153567|Uterine cancer NOS
C0153567|Uterus Cancer
C0153567|Cancer of the Uterus
C0153567|Malignant neoplasm of uterus, NOS
C0153567|Malignant Neoplasm of the Uterus
C0153567|Malignant Tumor of the Uterus
C0153567|Malignant Uterine Neoplasm
C0153567|Malignant Uterine Tumor
C0153567|Neoplasm malig;uterus
C0153567|malignant neosplasm of the uterus
C0153569|Malignant neoplasm of endocervix
C0153569|Endocervix
C0153569|malignant neoplasm of cervical canal (diagnosis)
C0153569|malignant neoplasm of endocervical canal
C0153569|malignant neoplasm of endocervical canal (diagnosis)
C0153569|malignant neoplasm of cervical canal
C0153569|malignant tumor of endocervical canal
C0153569|malignant tumor of cervical canal
C0153569|Malig neo endocervix
C0153569|cervical neoplasm malignant endocervix
C0153569|malignant neoplasm of endocervix (diagnosis)
C0153569|Malignant neoplasm of endocervix (disorder)
C0153569|Malignant neoplasm of endocervix NOS (disorder)
C0153569|Malignant neoplasm of endocervix NOS
C0153569|Malignant neoplasm of endocervical canal (disorder)
C0153569|Malignant Endocervical Neoplasm
C0153569|Malignant Endocervical Tumor
C0153569|Malignant Endocervix Neoplasm
C0153569|Malignant Endocervix Tumor
C0153569|Malignant Neoplasm of Uterine Endocervix
C0153569|Malignant Neoplasm of the Endocervix
C0153569|Malignant Neoplasm of the Uterine Endocervix
C0153569|Malignant Tumor of Endocervix
C0153569|Malignant Tumor of Uterine Endocervix
C0153569|Malignant Tumor of the Endocervix
C0153569|Malignant Tumor of the Uterine Endocervix
C0153569|Malignant Uterine Endocervix Neoplasm
C0153569|Malignant Uterine Endocervix Tumor
C0153569|Malignant neoplasm of cervical canal NOS
C0153570|Malignant neoplasm of exocervix
C0153570|Exocervix
C0153570|malignant neoplasm of exocervix (diagnosis)
C0153570|malignant tumor of exocervix
C0153570|Malig neo exocervix
C0153570|Malignant neoplasm of exocervix (disorder)
C0153570|Ca cervix uteri - exocervix (disorder)
C0153570|Ca cervix uteri - exocervix
C0153570|Cancer of exocervix
C0153570|Malignant Exocervical Neoplasm
C0153570|Malignant Exocervical Tumor
C0153570|Malignant Exocervix Neoplasm
C0153570|Malignant Exocervix Tumor
C0153570|Malignant Neoplasm of Uterine Exocervix
C0153570|Malignant Neoplasm of the Exocervix
C0153570|Malignant Neoplasm of the Uterine Exocervix
C0153570|Malignant Tumor of Uterine Exocervix
C0153570|Malignant Tumor of the Exocervix
C0153570|Malignant Tumor of the Uterine Exocervix
C0153570|Malignant Uterine Exocervix Neoplasm
C0153570|Malignant Uterine Exocervix Tumor
C0269193|anaplasia of cervix (diagnosis)
C0269193|dysplasia of cervix (uteri) anaplasia
C0269193|anaplasia of cervix
C0269193|Anaplasia of cervix (disorder)
C0269193|anaplasia; cervix
C2211948|malignant small cell neoplasm of uterus
C2211948|uterine neoplasm malignant small cell type
C2211948|malignant small cell neoplasm of uterus (diagnosis)
C2011421|uterine neoplasm malignant giant cell type
C2011421|giant cell type neoplasm of uterus (diagnosis)
C2011421|giant cell type neoplasm of uterus
C2018702|uterine neoplasm malignant spindle cell type
C2018702|spindle cell type neoplasm of uterus (diagnosis)
C2018702|spindle cell type neoplasm of uterus
C2075662|clear cell type neoplasm of uterus
C2075662|clear cell type neoplasm of uterus (diagnosis)
C2075662|uterine neoplasm malignant clear cell type
C0848454|Uterine carcinoma
C0848454|carcinoma of uterus (diagnosis)
C0848454|carcinoma of uterus
C0848454|Carcinoma;uterus
C0848454|carcinoma of the uterus
C2211972|myosarcoma of uterus (diagnosis)
C2211972|myosarcoma of uterus
C2211981|fibrosarcoma of uterus (diagnosis)
C2211981|fibrosarcoma of uterus
C2211991|malignant mesenchymoma of uterus (diagnosis)
C2211991|malignant mesenchymoma of uterus
C2211992|malignant mesonephroma of uterus (diagnosis)
C2211992|malignant mesonephroma of uterus
C2211993|Mullerian mixed tumor of uterus
C2211993|Mullerian mixed tumor of uterus (diagnosis)
C1704376|Uterine Corpus Carcinosarcoma
C1704376|malignant mesodermal mixed tumor of uterus
C1704376|malignant mesodermal mixed tumor of uterus (diagnosis)
C1704376|Mixed Müllerian Sarcoma of the Uterus
C1704376|Mixed Müllerian Sarcoma of Uterus
C1704376|Uterine Corpus Malignant Mixed Mesodermal (Müllerian) Tumor
C1704376|Uterine Corpus Malignant Mixed Müllerian Neoplasm
C1704376|Uterine Mixed Müllerian Sarcoma
C1704376|Uterine Corpus Malignant Mixed Müllerian Tumor
C1704376|Corpus Uteri Malignant Mixed Mesodermal Tumor
C1704376|Malignant Mixed Mesodermal Neoplasm of Uterine Body
C1704376|Malignant Mixed Mesodermal Neoplasm of Uterine Corpus
C1704376|Malignant Mixed Mesodermal Neoplasm of Uterus
C1704376|Malignant Mixed Mesodermal Neoplasm of the Uterine Body
C1704376|Malignant Mixed Mesodermal Neoplasm of the Uterine Corpus
C1704376|Malignant Mixed Mesodermal Neoplasm of the Uterus
C1704376|Malignant Mixed Mesodermal Tumor of Uterine Body
C1704376|Malignant Mixed Mesodermal Tumor of Uterine Corpus
C1704376|Malignant Mixed Mesodermal Tumor of Uterus
C1704376|Malignant Mixed Mesodermal Tumor of the Uterine Body
C1704376|Malignant Mixed Mesodermal Tumor of the Uterine Corpus
C1704376|Malignant Mixed Mesodermal Tumor of the Uterus
C1704376|Uterine Body Carcinosarcoma
C1704376|Uterine Body Malignant Mixed Mesodermal Neoplasm
C1704376|Uterine Body Malignant Mixed Mesodermal Tumor
C1704376|Uterine Carcinosarcoma
C1704376|Uterine Corpus Malignant Mixed Mesodermal Neoplasm
C1704376|Uterine Corpus Malignant Mixed Mesodermal Tumor
C1704376|Uterine Malignant Mixed Mesodermal Neoplasm
C1704376|Uterine Malignant Mixed Mesodermal Tumor
C1704376|Carcinosarcoma of Corpus Uteri
C1704376|Carcinosarcoma of Uterine Body
C1704376|Carcinosarcoma of Uterine Corpus
C1704376|Carcinosarcoma of Uterus
C1704376|Carcinosarcoma of the Corpus Uteri
C1704376|Carcinosarcoma of the Uterine Body
C1704376|Carcinosarcoma of the Uterine Corpus
C1704376|Carcinosarcoma of the Uterus
C2211995|malignant lymphoma of uterus
C2211995|malignant lymphoma of uterus (diagnosis)
C2211998|malignant plasmacytoma of uterus (diagnosis)
C2211998|malignant plasmacytoma of uterus
C2212000|malignant mastocytosis of uterus
C2212000|malignant mastocytosis of uterus (diagnosis)
C2217776|malignant neoplasm of uterus staging (diagnosis)
C2217776|malignant neoplasm of uterus staging
C2217776|uterine cancer staging
C2217776|malignant tumor of uterus staging
C0496821|Fundus uteri
C0496821|Malignant neoplasm of fundus uteri
C0496821|Malignant neoplasm of the fundus uteri
C0496821|malignant neoplasm of fundus of uterus
C0496821|malignant neoplasm of fundus of uterus (diagnosis)
C0496821|malignant tumor of fundus of uterus
C0496821|Malignant neoplasm of fundus of corpus uteri
C0496821|Malignant neoplasm of fundus of corpus uteri (disorder)
C0496818|Isthmus uteri
C0496818|Malignant neoplasm of isthmus uteri
C0496818|Malignant neoplasm of isthmus of uterus
C0496818|malignant neoplasm of isthmus of uterus (diagnosis)
C0496818|malignant tumor of isthmus of uterus
C0496818|Malignant neoplasm of isthmus of uterine body NOS (disorder)
C0496818|Malignant neoplasm of isthmus of uterine body NOS
C0496818|Malignant neoplasm of isthmus of uterine body
C0496818|Malignant neoplasm of isthmus of uterine body (disorder)
C2103110|adenosarcoma of uterus (diagnosis)
C2103110|adenosarcoma of uterus
C2103110|uterine adenosarcoma
C2103110|Mullerian adenosarcoma of the uterus
C2103110|Adenosarcoma of the uterus
C2103110|Adenosarcoma of uterus (disorder)
C2006983|carcinofibroma of uterus
C2006983|carcinofibroma of uterus (diagnosis)
C0280630|Uterine Carcinosarcoma
C0280630|Carcinosarcoma of the Uterus
C0280630|Uterine Malignant Mixed Mesodermal (Mullerian) Tumor
C0280630|Malignant Mixed Mesodermal (Mullerian) Tumor of the Uterus
C0280630|carcinosarcoma of uterus (diagnosis)
C0280630|carcinosarcoma of uterus
C0280630|Carcinosarcoma of uterus (disorder)
C0280630|Carcinosarcoma uterus
C0280630|Carcino-sarcoma uterus
C0280630|carcinosarcoma, uterine
C0280630|mixed Mullerian sarcoma, uterine
C0280630|uterine mixed Mullerian sarcoma
C0280630|Mullerian sarcoma, uterine mixed
C0280630|Mullerian tumor, uterine mixed
C0153584|Malignant neoplasm of uterine adnexa
C0153584|Malignant neoplasm of uterine adnexa, unspecified
C0153584|Uterine adnexa, unspecified
C0153584|Malignant neoplasm of uterine adnexa (disorder)
C0153584|malignant neoplasm of uterine adnexa (diagnosis)
C0153584|malignant tumor of uterine adnexa
C0153584|Mal neo adnexa NOS
C0153584|Malignant neoplasm of uterine adnexa, unspecified site
C0153584|[X]Malignant neoplasm of uterine adnexa, unspecified (disorder)
C0153584|Malignant neoplasm of uterine adnexa NOS (disorder)
C0153584|Malignant neoplasm of uterine adnexa NOS
C0153584|[X]Malignant neoplasm of uterine adnexa, unspecified
C0153584|Malignant neoplasm of uterine adnexa, NOS
C2960452|Malignant epithelial neoplasm of uterus (disorder)
C2960452|Malignant epithelial neoplasm of uterus
C2960452|Carcinoma of uterus
C0280631|Uterine leiomyosarcoma
C0280631|leiomyosarcoma of uterus
C0280631|leiomyosarcoma of uterus (diagnosis)
C0280631|Leiomyosarcoma of uterus (disorder)
C0280631|Leiomyosarcoma of the uterus
C0280631|Leiomyosarcoma - uterus
C0280631|leiomyosarcoma, uterine
C0280631|Corpus Uteri Leiomyosarcoma
C0280631|Leiomyosarcoma of Body of Uterus
C0280631|Leiomyosarcoma of Corpus Uteri
C0280631|Leiomyosarcoma of Uterine Body
C0280631|Leiomyosarcoma of Uterine Corpus
C0280631|Leiomyosarcoma of the Body of Uterus
C0280631|Leiomyosarcoma of the Corpus Uteri
C0280631|Leiomyosarcoma of the Uterine Body
C0280631|Leiomyosarcoma of the Uterine Corpus
C0280631|Uterine Body Leiomyosarcoma
C0280631|Uterine Corpus Leiomyosarcoma
C0280631|Body of Uterus Leiomyosarcoma
C3164916|Malignant mixed Mullerian tumor of uterus
C3164916|Malignant mixed Mullerian tumour of uterus
C3164916|Malignant mixed Mullerian tumor of uterus (disorder)
C0153572|Malignant neoplasm of placenta
C0153572|malignant neoplasm of placenta (diagnosis)
C0153572|malignant tumor of placenta
C0153572|Malignant neopl placenta
C0153572|placental cancer
C0153572|Malignant neoplasm of placenta (disorder)
C0153572|Cancer of placenta
C0153572|DECIDUOMA, MALIGNANT
C0153572|Malignant Placental Neoplasm
C0153572|Malignant Tumor of the Placenta
C0153572|Malignant Neoplasm of the Placenta
C0153572|Malignant Placental Tumor
C0153572|Malignant Placenta Neoplasm
C0153572|Malignant Placenta Tumor
C0153572|Neoplasm malig;placenta
C0153572|malignant neosplasm of the placenta
C2211985|adult type pleomorphic rhabdomyosarcoma of uterus (diagnosis)
C2211985|uterine rhabdomyosarcoma pleomorphic, adult type
C2211985|adult type pleomorphic rhabdomyosarcoma of uterus
C3468483|endometrial cancer susceptibility (diagnosis)
C3468483|endometrial cancer susceptibility
C0007103|Endometrium
C0007103|Malignant neoplasm of endometrium
C0007103|Endometrial neoplasms malignant
C0007103|malignant neoplasm of endometrium (diagnosis)
C0007103|uterine neoplasm, malignant - of the endometrium
C0007103|Endometrial Cancer
C0007103|Endometrial neoplasm malignant
C0007103|Malignant Endometrial Neoplasm
C0007103|malignant neoplasm of the endometrium
C0007103|Neoplasm malig;endometrial
C1879358|Primary malignant neoplasm of endometrium
C1879358|Malignant neoplasm of endometrium
C1879358|Primary malignant neoplasm of endometrium (diagnosis)
C1879358|uterine neoplasm, malignant - of the endometrium primary
C1879358|Cancer of endometrium
C1879358|Primary malignant neoplasm of endometrium (disorder)
C0008493|Malignant hydatidiform mole
C0008493|Chorioadenomas
C0008493|Hydatidiform Mole, Invasive
C0008493|Hydatidiform Moles, Invasive
C0008493|Invasive Hydatidiform Moles
C0008493|Invasive Moles
C0008493|Moles, Invasive
C0008493|Moles, Invasive Hydatidiform
C0008493|Invasive Hydatidiform Mole
C0008493|Mole, Invasive
C0008493|Mole, Invasive Hydatidiform
C0008493|invasive hydatidiform mole (diagnosis)
C0008493|molar pregnancy, invasive (non-metastatic GTD)
C0008493|Chorioadenoma destruens
C0008493|Chorioadenoma
C0008493|Hydatidiform Mole, Invasive [Disease/Finding]
C0008493|Invasive Mole
C0008493|Mole;malignant
C0008493|Molar pregnancy with invasive hydatidiform mole
C0008493|Malignant hydatidiform mole (disorder)
C0008493|Molar pregnancy with malignant hydatidiform mole
C0008493|Molar pregnancy with chorioadenoma destruens
C0008493|Invasive mole - placenta
C0008493|Molar pregnancy with chorioadenoma
C0008493|IM - Invasive mole
C0008493|Choriadenoma (destruens)
C0008493|Molar pregnancy with invasive mole
C0008493|Molar pregnancy with invasive hydatidiform mole (disorder)
C0008493|[M]Chorioadenoma destruens
C0008493|[M]Invasive hydatidiform mole
C0008493|[M]Chorioadenoma
C0008493|Hydatidiform mole malignant
C0008493|Invasive hydatidiform mole (morphologic abnormality)
C0008493|GTT, invasive mole
C0008493|gestational trophoblastic tumor, invasive mole
C0008493|destructive; mole
C0008493|hydatidiform mole; invasive
C0008493|hydatidiform mole; malignant
C0008493|invasive; hydatidiform mole
C0008493|invasive; mole
C0008493|malignant; hydatidiform mole
C0008493|malignant; mole, hydatidiform
C0008493|mole; destructive
C0008493|mole; hydatidiform, invasive
C0008493|mole; hydatidiform, malignant
C0008493|mole; invasive
C0008493|mole; malignant, hydatidiform mole
C0008493|Invasive mole, NOS
C0008493|Invasive Gestational Trophoblastic Neoplasm
C0008493|Malignant hydatid mole
C0008493|Invasive hydatidiform mole (disorder)
C0008493|malignant mole
C1299275|Primary malignant neoplasm of body of uterus
C1299275|Primary malignant neoplasm of body of uterus (disorder)
C1299275|primary malignant neoplasm of corpus uteri
C1299275|primary malignant neoplasm of corpus uteri (diagnosis)
C1299275|uterine neoplasm, malignant - corpus uteri primary
C2703078|Malignant neoplasm of placenta
C2703078|Primary malignant neoplasm of placenta
C2703078|placental neoplasm malignant primary
C2703078|Primary malignant neoplasm of placenta (diagnosis)
C2703078|Primary malignant neoplasm of placenta (disorder)
C1263776|Overlapping malignant neoplasm of body of uterus (disorder)
C1263776|Overlapping malignant neoplasm of body of uterus
C1263776|Overlapping malignant neoplasm of corpus uteri
C1306053|Primary malignant neoplasm of isthmus of uterus (disorder)
C1306053|Primary malignant neoplasm of isthmus of uterus
C1314886|Primary malignant neoplasm of parametrium (disorder)
C1314886|Primary malignant neoplasm of parametrium
C0007847|Malignant neoplasm of cervix uteri
C0007847|Malignant neoplasm of cervix uteri, unspecified
C0007847|Cervix uteri, unspecified
C0007847|Malignant neoplasm of uterine cervix
C0007847|cancer of cervix
C0007847|malignant neoplasm of cervix
C0007847|cervical cancer
C0007847|malignant neoplasm of cervix (diagnosis)
C0007847|malignant cervical neoplasm
C0007847|Malignant tumor of cervix
C0007847|Mal neo cervix uteri NOS
C0007847|Cervix neoplasms malignant
C0007847|Malignant neoplasm of cervix uteri, unspecified site
C0007847|malignant neoplasm of cervix uteri (diagnosis)
C0007847|cervical neoplasm malignant cervix uteri
C0007847|Malignant tumour of cervix (disorder)
C0007847|Malignant neoplasm of cervix uteri NOS (disorder)
C0007847|Malignant tumour of cervix
C0007847|Malignant neoplasm of cervix uteri NOS
C0007847|Cancer of the uterine cervix
C0007847|Malignant tumor of cervix (disorder)
C0007847|Malignant Cervical Tumor
C0007847|Malignant Cervix Neoplasm
C0007847|Malignant Cervix Tumor
C0007847|Malignant Cervix Uteri Neoplasm
C0007847|Malignant Cervix Uteri Tumor
C0007847|Malignant Neoplasm of the Cervix Uteri
C0007847|Malignant Neoplasm of the Cervix
C0007847|Malignant Neoplasm of the Uterine Cervix
C0007847|Malignant Tumor of Cervix Uteri
C0007847|Malignant Tumor of Uterine Cervix
C0007847|Malignant Tumor of the Cervix Uteri
C0007847|Malignant Tumor of the Cervix
C0007847|Malignant Tumor of the Uterine Cervix
C0007847|Malignant Uterine Cervix Neoplasm
C0007847|Malignant Uterine Cervix Tumor
C0007847|Neoplasm malig;cervix
C0007847|malignant neosplasm of the cervix
C0346995|metastasis of malignant neoplasm to the uterus
C0346995|metastasis of malignant neoplasm to uterus (diagnosis)
C0346995|metastasis of malignant neoplasm to uterus
C0346995|Metastases to uterus
C0346995|uterine neoplasm malignant secondary
C0346995|Secondary malignant neoplasm of uterus
C0346995|Secondary malignant neoplasm of uterus (diagnosis)
C0346995|Cancer metastatic to uterus
C0346995|Metastasis to uterus
C0346995|Metastatic malignant neoplasm to uterus
C0346995|Secondary malignant neoplasm of uterus (disorder)
C0346995|Metastatic malignant neoplasm to uterus, NOS
C0346995|Secondary malignant neoplasm of uterus, NOS
C1282495|metastasis from malignant neoplasm of uterus
C1282495|metastasis from malignant neoplasm of uterus (diagnosis)
C1282495|Metastasis from malignant tumor of uterus (disorder)
C1282495|Metastasis from malignant tumor of uterus
C1282495|Metastasis from malignant tumour of uterus
C3838720|Primary malignant neoplasm of uterus (disorder)
C3838720|Primary malignant neoplasm of uterus
C1336899|Hemangiosarcoma of Uterus
C1336899|Hemangiosarcoma of the Uterus
C1336899|Angiosarcoma of Uterus
C1336899|Angiosarcoma of the Uterus
C1336899|Uterine Angiosarcoma
C1336899|Uterine Hemangiosarcoma
C2217769|malignant neoplasm of uterus stage IIa
C2217769|malignant neoplasm of uterus stage IIa (diagnosis)
C2217769|malignant tumor of uterus stage IIa
C2217769|uterine cancer stage IIa
C2111694|large cell carcinoma of uterus with rhabdoid phenotype
C2111694|large cell carcinoma of uterus with rhabdoid phenotype (diagnosis)
C2111694|uterine malignant carcinoma large cell with rhabdoid phenotype
C2018413|spindle cell carcinoma of uterus
C2018413|spindle cell carcinoma of uterus (diagnosis)
C2033322|papillary squamous cell carcinoma of uterus
C2033322|papillary squamous cell carcinoma of uterus (diagnosis)
C2211953|nonkeratinizing squamous cell carcinoma of uterus
C2211953|nonkeratinizing squamous cell carcinoma of uterus (diagnosis)
C2211953|uterine malignant carcinoma squamous cell small cell nonkeratinizing
C2211954|adenoid squamous cell carcinoma of uterus
C2211954|adenoid squamous cell carcinoma of uterus (diagnosis)
C2211956|basaloid squamous cell carcinoma of uterus (diagnosis)
C2211956|basaloid squamous cell carcinoma of uterus
C2075854|cloacogenic carcinoma of uterus
C2075854|cloacogenic carcinoma of uterus (diagnosis)
C2211979|mast cell sarcoma of uterus
C2211979|mast cell sarcoma of uterus (diagnosis)
C2188881|lymphocyte-rich nodular Hodgkin's lymphoma of uterus (diagnosis)
C2188881|lymphocyte-rich nodular Hodgkin's lymphoma of uterus
C2188883|nodular sclerosing Hodgkin's lymphoma in cellular phase of uterus (diagnosis)
C2188883|nodular sclerosing Hodgkin's lymphoma in cellular phase of uterus
C2188885|grade 2 nodular sclerosing Hodgkin's lymphoma of uterus
C2188885|grade 2 nodular sclerosing Hodgkin's lymphoma of uterus (diagnosis)
C2188897|lymphoplasmacytic lymphoma of uterus (diagnosis)
C2188897|lymphoplasmacytic lymphoma of uterus
C2188899|marginal zone B-cell lymphoma of uterus
C2188899|marginal zone B-cell lymphoma of uterus (diagnosis)
C2188900|mature T-cell lymphoma of uterus (diagnosis)
C2188900|mature T-cell lymphoma of uterus
C2188903|NK/T-cell lymphoma of uterus
C2188903|NK/T-cell lymphoma of uterus (diagnosis)
C2212001|Sezary syndrome of uterus
C2212001|Sezary syndrome of uterus (diagnosis)
C2111693|large cell carcinoma of uterus (diagnosis)
C2111693|large cell carcinoma of uterus
C2012125|glassy cell carcinoma of uterus (diagnosis)
C2012125|glassy cell carcinoma of uterus
C2033341|papillary transitional cell carcinoma of uterus (diagnosis)
C2033341|papillary transitional cell carcinoma of uterus
C2011238|giant cell and spindle cell carcinoma of uterus
C2011238|giant cell and spindle cell carcinoma of uterus (diagnosis)
C2007043|carcinoma of uterus with osteoclast-like giant cells
C2007043|carcinoma of uterus with osteoclast-like giant cells (diagnosis)
C2007043|uterine carcinoma with osteoclast-like giant cells
C0279764|papillary carcinoma of uterus
C0279764|papillary carcinoma of uterus (diagnosis)
C0279764|endometrial papillary carcinoma
C0279764|carcinoma of the uterus, papillary
C0279764|carcinoma, papillary, endometrial
C0279764|papillary carcinoma of the uterus
C0279764|uterine cancer, papillary carcinoma
C0279764|uterine corpus cancer, papillary carcinoma
C0279764|uterus cancer, papillary carcinoma
C2019462|uterine malignant carcinoma squamous cell with horn formation
C2019462|squamous cell carcinoma of uterus with horn formation (diagnosis)
C2019462|squamous cell carcinoma of uterus with horn formation
C2019462|squamous cell carcinoma with horn formation of uterus
C2075582|clear cell squamous cell carcinoma of uterus
C2075582|clear cell squamous cell carcinoma of uterus (diagnosis)
C2211957|Schneiderian carcinoma of uterus
C2211957|Schneiderian carcinoma of uterus (diagnosis)
C2211957|uterine malignant carcinoma Schneiderian
C2211958|basaloid carcinoma of uterus
C2211958|basaloid carcinoma of uterus (diagnosis)
C2188891|grade 1 follicular lymphoma of uterus (diagnosis)
C2188891|grade 1 follicular lymphoma of uterus
C2188892|grade 2 follicular lymphoma of uterus
C2188892|grade 2 follicular lymphoma of uterus (diagnosis)
C2217767|malignant neoplasm of uterus stage Ib
C2217767|malignant neoplasm of uterus stage Ib (diagnosis)
C2217767|malignant tumor of uterus stage Ib
C2217767|uterine cancer stage Ib
C2217775|malignant neoplasm of uterus stage IVb
C2217775|malignant neoplasm of uterus stage IVb (diagnosis)
C2217775|malignant tumor of uterus stage IVb
C2217775|uterine cancer stage IVb
C2111825|polygonal cell carcinoma of uterus (diagnosis)
C2111825|polygonal cell carcinoma of uterus
C2018579|spindle cell squamous cell carcinoma of uterus (diagnosis)
C2018579|spindle cell squamous cell carcinoma of uterus
C2211960|mucoepidermoid carcinoma of uterus
C2211960|mucoepidermoid carcinoma of uterus (diagnosis)
C2017462|solid carcinoma of uterus (diagnosis)
C2017462|solid carcinoma of uterus
C2211984|malignant solitary fibrous tumor of uterus (diagnosis)
C2211984|malignant solitary fibrous tumor of uterus
C2188898|mantle cell lymphoma of uterus (diagnosis)
C2188898|mantle cell lymphoma of uterus
C2188895|large B-cell diffuse lymphoma of uterus
C2188895|large B-cell diffuse lymphoma of uterus (diagnosis)
C2113667|precursor B-cell lymphoblastic lymphoma of uterus (diagnosis)
C2113667|precursor B-cell lymphoblastic lymphoma of uterus
C2113807|precursor T-cell lymphoblastic lymphoma of uterus (diagnosis)
C2113807|precursor T-cell lymphoblastic lymphoma of uterus
C2103109|undifferentiated carcinoma of uterus (diagnosis)
C2103109|undifferentiated carcinoma of uterus
C2217766|malignant neoplasm of uterus stage Ia
C2217766|malignant neoplasm of uterus stage Ia (diagnosis)
C2217766|malignant tumor of uterus stage Ia
C2217766|uterine cancer stage Ia
C2111760|large cell neuroendocrine carcinoma of uterus
C2111760|large cell neuroendocrine carcinoma of uterus (diagnosis)
C2211950|anaplastic carcinoma of uterus
C2211950|anaplastic carcinoma of uterus (diagnosis)
C2211952|micropapillary transitional cell carcinoma of uterus
C2211952|micropapillary transitional cell carcinoma of uterus (diagnosis)
C2018619|spindle cell transitional cell carcinoma of uterus (diagnosis)
C2018619|spindle cell transitional cell carcinoma of uterus
C2211963|medullary carcinoma of uterus (diagnosis)
C2211963|medullary carcinoma of uterus
C2188880|mixed cellularity Hodgkin's lymphoma of uterus
C2188880|mixed cellularity Hodgkin's lymphoma of uterus (diagnosis)
C2188878|Hodgkin's disease, lymphocytic depletion of uterus
C2188878|Hodgkin's disease, lymphocytic depletion of uterus (diagnosis)
C2188896|immunoblastic large B-cell diffuse lymphoma of uterus (diagnosis)
C2188896|immunoblastic large B-cell diffuse lymphoma of uterus
C2188894|malignant histiocytosis of uterus (diagnosis)
C2188894|malignant histiocytosis of uterus
C2217773|malignant neoplasm of uterus stage IIIc (diagnosis)
C2217773|malignant neoplasm of uterus stage IIIc
C2217773|uterine cancer stage IIIc
C2217773|malignant tumor of uterus stage IIIc
C2109332|keratinizing squamous cell carcinoma of uterus (diagnosis)
C2109332|keratinizing squamous cell carcinoma of uterus
C2138886|large cell nonkeratinizing squamous cell carcinoma of uterus (diagnosis)
C2138886|uterine malignant carcinoma squamous cell large cell nonkeratinizing
C2138886|large cell nonkeratinizing squamous cell carcinoma of uterus
C2211955|microinvasive squamous cell carcinoma of uterus (diagnosis)
C2211955|microinvasive squamous cell carcinoma of uterus
C2188884|grade 1 nodular sclerosing Hodgkin's lymphoma of uterus (diagnosis)
C2188884|grade 1 nodular sclerosing Hodgkin's lymphoma of uterus
C2046746|Hodgkin's sarcoma of uterus
C2046746|Hodgkin's sarcoma of uterus (diagnosis)
C2188902|mixed small and large cell diffuse lymphoma of uterus
C2188902|mixed small and large cell diffuse lymphoma of uterus (diagnosis)
C2113738|precursor cell lymphoblastic lymphoma of uterus (diagnosis)
C2113738|precursor cell lymphoblastic lymphoma of uterus
C2009896|fusiform type small cell carcinoma of uterus
C2009896|fusiform type small cell carcinoma of uterus (diagnosis)
C2189372|verrucous carcinoma of uterus
C2189372|verrucous carcinoma of uterus (diagnosis)
C2145473|transitional cell carcinoma of uterus (diagnosis)
C2145473|transitional cell carcinoma of uterus
C2138465|cribriform carcinoma of uterus (diagnosis)
C2138465|cribriform carcinoma of uterus
C2211961|adenosquamous carcinoma of uterus (diagnosis)
C2211961|adenosquamous carcinoma of uterus
C2007053|carcinoma simplex of uterus
C2007053|carcinoma simplex of uterus (diagnosis)
C2007053|carcinoma simplex of urethra (diagnosis)
C2007053|carcinoma simplex of urethra
C2012551|granular cell carcinoma of uterus (diagnosis)
C2012551|granular cell carcinoma of uterus
C2182940|desmoplastic small round cell tumor of uterus (diagnosis)
C2182940|desmoplastic small round cell tumor of uterus
C2046534|uterine malignant lymphoma Hodgkin's and non-Hodgkin's
C2046534|composite Hodgkin's and non-Hodgkin's lymphoma of uterus (diagnosis)
C2046534|composite Hodgkin's and non-Hodgkin's lymphoma of uterus
C2188904|small B-cell lymphocytic lymphoma of uterus (diagnosis)
C2188904|small B-cell lymphocytic lymphoma of uterus
C2217770|malignant neoplasm of uterus stage IIb
C2217770|malignant neoplasm of uterus stage IIb (diagnosis)
C2217770|uterine cancer stage IIb
C2217770|malignant tumor of uterus stage IIb
C2217771|malignant neoplasm of uterus stage IIIa (diagnosis)
C2217771|malignant neoplasm of uterus stage IIIa
C2217771|uterine cancer stage IIIa
C2217771|malignant tumor of uterus stage IIIa
C2217772|malignant neoplasm of uterus stage IIIb (diagnosis)
C2217772|malignant neoplasm of uterus stage IIIb
C2217772|malignant tumor of uterus stage IIIb
C2217772|uterine cancer stage IIIb
C2211949|malignant epithelioma of uterus (diagnosis)
C2211949|malignant epithelioma of uterus
C2211951|small cell carcinoma of uterus (diagnosis)
C2211951|small cell carcinoma of uterus
C2211962|epithelial-myoepithelial carcinoma of uterus (diagnosis)
C2211962|epithelial-myoepithelial carcinoma of uterus
C2046606|Hodgkin's granuloma of uterus
C2046606|Hodgkin's granuloma of uterus (diagnosis)
C2188890|follicular lymphoma of uterus
C2188890|follicular lymphoma of uterus (diagnosis)
C2188901|angioimmunoblastic T-cell lymphoma of uterus (diagnosis)
C2188901|angioimmunoblastic T-cell lymphoma of uterus
C2188901|angioimmunoblastic lymphadenopathy with dysproteinemia (AILD) of uterus
C2019461|squamous cell carcinoma of uterus (diagnosis)
C2019461|squamous cell carcinoma of uterus
C2217768|malignant neoplasm of uterus stage Ic
C2217768|malignant neoplasm of uterus stage Ic (diagnosis)
C2217768|malignant tumor of uterus stage Ic
C2217768|uterine cancer stage Ic
C2217774|malignant neoplasm of uterus stage IVa (diagnosis)
C2217774|malignant neoplasm of uterus stage IVa
C2217774|malignant tumor of uterus stage IVa
C2217774|uterine cancer stage IVa
C2082473|pleomorphic carcinoma of uterus (diagnosis)
C2082473|pleomorphic carcinoma of uterus
C2011273|giant cell carcinoma of uterus (diagnosis)
C2011273|giant cell carcinoma of uterus
C2142943|pseudosarcomatous carcinoma of uterus
C2142943|pseudosarcomatous carcinoma of uterus (diagnosis)
C2200280|lymphoepithelial squamous cell carcinoma of uterus (diagnosis)
C2200280|lymphoepithelial squamous cell carcinoma of uterus
C2211959|adenoid cystic carcinoma of uterus (diagnosis)
C2211959|adenoid cystic carcinoma of uterus
C2188877|lymphocyte-rich Hodgkin's lymphoma of uterus (diagnosis)
C2188877|lymphocyte-rich Hodgkin's lymphoma of uterus
C2188876|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of uterus
C2188876|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of uterus (diagnosis)
C2188882|nodular sclerosing Hodgkin's lymphoma of uterus (diagnosis)
C2188882|nodular sclerosing Hodgkin's lymphoma of uterus
C2188893|grade 3 follicular lymphoma of uterus (diagnosis)
C2188893|grade 3 follicular lymphoma of uterus
C2188879|Hodgkin's disease, lymphocytic depletion, reticular of uterus (diagnosis)
C2188879|Hodgkin's disease, lymphocytic depletion, reticular of uterus
C0153595|Undescended testis
C0153595|Malignant neoplasm of undescended testis
C0153595|Malignant tumor of undescended testis
C0153595|malignant neoplasm of undescended testis (diagnosis)
C0153595|malignant neoplasm of retained testis
C0153595|malignant neoplasm of retained testis (diagnosis)
C0153595|malignant tumor of retained testis
C0153595|Mal neo undescend testis
C0153595|Malignant tumor of retained testis (disorder)
C0153595|Malignant tumour of retained testis
C0153595|Malignant neoplasm of undescended testis NOS (disorder)
C0153595|Cancer of intra-abdominal testis
C0153595|Malignant neoplasm of undescended testis NOS
C0153595|Malignant neoplasm of testis, undescended
C0153595|Cancer of undescended testis
C0153595|Malignant tumour of undescended testis
C0153595|Malignant tumor of undescended testis (disorder)
C0348906|Malignant neoplasm of descended testis
C0348906|Descended testis
C0348906|testicular neoplasm malignant descended testis
C0348906|Malignant neoplasm of descended testis (diagnosis)
C0348906|Malignant neoplasm of descended testis (disorder)
C0348906|Primary malignant neoplasm of descended testis (diagnosis)
C0348906|Primary malignant neoplasm of descended testis
C0348906|testicular neoplasm malignant descended testis primary
C0348906|Primary malignant neoplasm of descended testis (disorder)
C0348906|Malignant neoplasm of testis, descended
C0153594|Malignant neoplasm of testis
C0153594|testicular cancer
C0153594|Malignant neoplasm of testis, unspecified
C0153594|Testis, unspecified
C0153594|testicular cancer (diagnosis)
C0153594|malignant neoplasm of testis (diagnosis)
C0153594|Cancers, Testis
C0153594|Testis Cancers
C0153594|Cancer, Testicular
C0153594|Cancers, Testicular
C0153594|Testicular Cancers
C0153594|malignant tumor of testis
C0153594|Cancer of testis
C0153594|Malignant neoplasm of testis NOS
C0153594|Malignant neoplasm of testis, unspecified whether descended or undescended
C0153594|Cancer, Testis
C0153594|Malignant neoplasm of testis NOS (disorder)
C0153594|Testis cancer
C0153594|Testis--Cancer
C0153594|Testis neoplasm malignant
C0153594|Testicular neoplasms malignant
C0153594|Cancer of the Testis
C0153594|Cancer of the Testes
C0153594|Malignant tumour of testis
C0153594|Malignant tumor of testis (disorder)
C0153594|testicle cancer
C0153594|Malignant neoplasm of testis, NOS
C0153594|Malignant Neoplasm of the Testis
C0153594|Malignant Testicular Neoplasm
C0153594|Malignant Testicular Tumor
C0153594|Malignant Tumor of the Testis
C0153594|Neoplasm malig;testis
C0153594|malignant neosplasm of the testis
C0036631|Seminoma
C0036631|Seminomas
C0036631|Testicular seminoma
C0036631|seminoma of testis (diagnosis)
C0036631|seminoma of testis
C0036631|Seminoma (disorder)
C0036631|Seminoma (morphologic abnormality)
C0036631|Seminoma, no ICD-O subtype
C0036631|Seminoma [Disease/Finding]
C0036631|[M]Seminomas
C0036631|Seminoma testis
C0036631|[M]Seminomas (morphologic abnormality)
C0036631|[M]Seminoma NOS
C0036631|[M]Seminoma NOS (morphologic abnormality)
C0036631|malignant neoplasm seminoma
C0036631|seminoma (diagnosis)
C0036631|Seminoma, no ICD-O subtype (morphologic abnormality)
C0036631|Seminoma, no International Classification of Diseases for Oncology subtype
C0036631|Seminoma, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0036631|SEMINOMA, MALIGNANT
C0036631|Seminoma, Pure
C0036631|Testicular seminoma pure NOS
C0036631|Testicular seminoma (pure)
C0036631|Seminoma of testis (disorder)
C0036631|seminoma of the testis
C0036631|seminoma, testicular
C0036631|testicle cancer, seminoma
C0036631|testicular cancer, seminoma
C0036631|testis cancer, seminoma
C0036631|Seminoma, NOS
C0036631|Testicular Seminoma Pure
C0855193|Testicular choriocarcinoma stage I
C0855193|Stage I Testicular Choriocarcinoma AJCC v7
C0855193|Stage I Testicular Choriocarcinoma AJCC v6
C0855193|Stage I Testicular Choriocarcinoma
C0853869|Testicular choriocarcinoma stage II
C0853869|Stage II Testicular Choriocarcinoma AJCC v6
C0853869|Stage II Testicular Choriocarcinoma AJCC v7
C0853869|Stage II Testicular Choriocarcinoma
C0855184|Testicular choriocarcinoma stage III
C0855184|Stage III Testicular Choriocarcinoma AJCC v6
C0855184|Stage III Testicular Choriocarcinoma AJCC v7
C0855184|Stage III Testicular Choriocarcinoma
C0855194|Testicular embryonal carcinoma stage I
C0855194|Stage I Testicular Embryonal Carcinoma AJCC v6
C0855194|Stage I Testicular Embryonal Carcinoma AJCC v7
C0855194|Stage I Testicular Embryonal Carcinoma
C0855195|Testicular embryonal carcinoma stage II
C0855195|Stage II Testicular Embryonal Carcinoma AJCC v6
C0855195|Stage II Testicular Embryonal Carcinoma AJCC v7
C0855195|Stage II Testicular Embryonal Carcinoma
C0855196|Testicular embryonal carcinoma stage III
C0855196|Stage III Testicular Embryonal Carcinoma AJCC v7
C0855196|Stage III Testicular Embryonal Carcinoma AJCC v6
C0855196|Stage III Testicular Embryonal Carcinoma
C0855203|Testicular germ cell tumour mixed stage I
C0855203|Stage I Testicular Mixed Germ Cell Tumor AJCC v6
C0855203|Stage I Testicular Mixed Germ Cell Tumor AJCC v7
C0855203|Testicular germ cell tumor mixed stage I
C0855203|Stage I Testicular Mixed Germ Cell Tumor
C0855199|Testicular germ cell tumour mixed stage II
C0855199|Stage II Testicular Mixed Germ Cell Tumor AJCC v7
C0855199|Stage II Testicular Mixed Germ Cell Tumor AJCC v6
C0855199|Testicular germ cell tumor mixed stage II
C0855199|Stage II Testicular Mixed Germ Cell Tumor
C0855204|Testicular germ cell tumour mixed stage III
C0855204|Stage III Testicular Mixed Germ Cell Tumor AJCC v6
C0855204|Stage III Testicular Mixed Germ Cell Tumor AJCC v7
C0855204|Testicular germ cell tumor mixed stage III
C0855204|Stage III Testicular Mixed Germ Cell Tumor
C0855205|Testicular malignant teratoma stage I
C0855206|Testicular malignant teratoma stage II
C0855207|Testicular malignant teratoma stage III
C0855208|Testicular seminoma (pure) stage I
C0855209|Testicular seminoma (pure) stage II
C0855210|Testicular seminoma (pure) stage III
C0855213|Testicular yolk sac tumour stage I
C0855213|Stage I Testicular Yolk Sac Tumor AJCC v6
C0855213|Stage I Testicular Yolk Sac Tumor AJCC v7
C0855213|Testicular endodermal sinus tumor stage I
C0855213|Testicular endodermal sinus tumour stage I
C0855213|Testicular yolk sac tumor stage I
C0855213|Stage I Testicular Yolk Sac Tumor
C0855214|Testicular yolk sac tumour stage II
C0855214|Stage II Testicular Yolk Sac Tumor AJCC v6
C0855214|Stage II Testicular Yolk Sac Tumor AJCC v7
C0855214|Testicular endodermal sinus tumour stage II
C0855214|Testicular yolk sac tumor stage II
C0855214|Testicular endodermal sinus tumor stage II
C0855214|Stage II Testicular Yolk Sac Tumor
C0855215|Testicular yolk sac tumour stage III
C0855215|Stage III Testicular Yolk Sac Tumor AJCC v6
C0855215|Stage III Testicular Yolk Sac Tumor AJCC v7
C0855215|Testicular yolk sac tumor stage III
C0855215|Testicular endodermal sinus tumor stage III
C0855215|Testicular endodermal sinus tumour stage III
C0855215|Stage III Testicular Yolk Sac Tumor
C0855197|Testicular cancer (excluding germ cell or trophoblastic cancer)
C0855197|Testicular ca. (no germ/tropho.)
C0855197|testicular cancer
C0855197|Testicular germ cell cancer NOS
C0855197|Testicular malignant germ cell tumor NOS
C0855197|Testicular germ cell cancer
C0855197|Malignant germ cell tumor of testis
C0855197|Malignant germ cell tumour of testis
C0855197|Malignant germ cell tumor of testis (disorder)
C0855197|Testicular malignant germ cell tumor
C0855197|Malignant Germ Cell Neoplasm of Testis
C0855197|Malignant Germ Cell Neoplasm of the Testis
C0855197|Malignant Germ Cell Tumor of the Testis
C0855197|Malignant Testicular Germ Cell Neoplasm
C0855197|Malignant Testicular Germ Cell Tumor
C0238449|choriocarcinoma of testis
C0238449|choriocarcinoma of testis (diagnosis)
C0238449|testicular choriocarcinoma
C0238449|Testicular choriocarcinoma NOS
C0238449|Choriocarcinoma of testis (disorder)
C0238449|choriocarcinoma of the testis
C0238449|choriocarcinoma, testicular
C0238449|testicle cancer, choriocarcinoma
C0238449|testicular cancer, choriocarcinoma
C0238449|testis cancer, choriocarcinoma
C0238448|embryonal carcinoma of testis (diagnosis)
C0238448|embryonal carcinoma of testis
C0238448|Testicular embryonal carcinoma
C0238448|Testicular embryonal carcinoma NOS
C0238448|embryonal carcinoma of the testis
C0238448|embryonal carcinoma, testicular
C0238448|testicle cancer, embryonal
C0238448|testicular cancer, embryonal
C0238448|testis cancer, embryonal
C2363951|Testicular germ cell cancer metastatic
C1096715|Testicular cancer metastatic
C1096715|Metastatic Malignant Testicular Germ Cell Tumor
C1096715|Metastatic Testicular Cancer
C2747856|Testicular choriocarcinoma recurrent
C0278841|Recurrent Malignant Testicular Germ Cell Tumor
C0278841|Recurrent Testicular Cancer
C0278841|Testis cancer recurrent
C0278841|cancer of the testis, recurrent
C0278841|cancer of the testis, relapsed
C0278841|carcinoma of the testis, recurrent
C0278841|carcinoma of the testis, relapsed
C0278841|recurrent cancer of the testis
C0278841|recurrent carcinoma of the testis
C0278841|recurrent or refractory testicular cancer
C0278841|recurrent testis cancer
C0278841|relapsed cancer of the testis
C0278841|relapsed carcinoma of the testis
C0278841|relapsed testicular cancer
C0278841|relapsed testis cancer
C0278841|testicle cancer, recurrent
C0278841|testicle cancer, refractory
C0278841|testicle cancer, relapsed
C0278841|testicular cancer, recurrent
C0278841|testicular cancer, relapsed
C0278841|testis cancer, recurrent
C0278841|testis cancer, relapsed
C0278841|Recurrent Cancer of Testis
C0278841|Relapsed Cancer of Testis
C2845878|Malignant neoplasm of unspecified testis, unspecified whether descended or undescended
C2845878|Malig neoplasm of unsp testis, unsp descended or undescended
C2845879|Malignant neoplasm of right testis, unspecified whether descended or undescended
C2845879|Malig neoplm of right testis, unsp descended or undescended
C2845880|Malignant neoplasm of left testis, unspecified whether descended or undescended
C2845880|Malig neoplasm of left testis, unsp descended or undescended
C2212306|testicular neoplasm malignant small cell type
C2212306|malignant small cell neoplasm of testis (diagnosis)
C2212306|malignant small cell neoplasm of testis
C2011413|giant cell type neoplasm of testis (diagnosis)
C2011413|giant cell type neoplasm of testis
C2011413|testicular neoplasm malignant giant cell type
C2018694|testicular neoplasm malignant spindle cell type
C2018694|spindle cell type neoplasm of testis (diagnosis)
C2018694|spindle cell type neoplasm of testis
C2075654|testicular neoplasm malignant clear cell type
C2075654|clear cell type neoplasm of testis
C2075654|clear cell type neoplasm of testis (diagnosis)
C0677483|carcinoma of testis (diagnosis)
C0677483|carcinoma of testis
C0677483|testicular carcinoma
C0677483|Carcinoma;testis
C0677483|Testicular Ca
C0677483|Carcinoma testis
C0677483|Carcinoma testes
C0677483|carcinoma of the testis
C2212309|adenocarcinoma of testis
C2212309|adenocarcinoma of testis (diagnosis)
C2212309|testicular adenocarcinoma
C2212312|malignant gonadal neoplasm of testis
C2212312|malignant gonadal neoplasm of testis (diagnosis)
C1336727|sarcoma of testis (diagnosis)
C1336727|sarcoma of testis
C1336727|Sarcoma of the Testis
C1336727|Testicular Sarcoma
C1336726|testicular myosarcoma rhabdomyosarcoma
C1336726|rhabdomyosarcoma of testis (diagnosis)
C1336726|rhabdomyosarcoma of testis
C1336726|Rhabdomyosarcoma of the Testis
C1336726|Testicular Rhabdomyosarcoma
C2242809|germinoma of testis
C2242809|germinoma of testis (diagnosis)
C1334154|malignant teratoma of testis
C1334154|malignant teratoma of testis (diagnosis)
C1334154|Testicular malignant teratoma
C1334154|Immature Teratoma of Testis
C1334154|Immature Teratoma of the Testis
C1334154|Immature Testicular Teratoma
C1334154|Malignant Teratoma of the Testis
C1334154|Malignant Testicular Teratoma
C1334154|Testicular Immature Teratoma
C1334154|Malignant teratoma of testis (disorder)
C2057624|malignant epithelioid trophoblastic tumor of testis
C2057624|malignant epithelioid trophoblastic tumor of testis (diagnosis)
C0349644|Primary Testicular Lymphoma
C0349644|malignant lymphoma of testis (diagnosis)
C0349644|malignant lymphoma of testis
C0349644|Malignant lymphoma of testis (disorder)
C0349644|Lymphoma of Testis
C0349644|Lymphoma of the Testis
C0349644|Testicular Lymphoma
C2212324|malignant plasmacytoma of testis (diagnosis)
C2212324|malignant plasmacytoma of testis
C2212326|malignant mastocytosis of testis
C2212326|malignant mastocytosis of testis (diagnosis)
C2217647|malignant neoplasm of testis staging
C2217647|malignant neoplasm of testis staging (diagnosis)
C2217647|malignant testicular neoplasm staging
C2217647|malignant tumor of testis staging
C2217647|testicular cancer staging
C2188087|undifferentiated carcinoma of testis (diagnosis)
C2188087|undifferentiated carcinoma of testis
C2057597|choriocarcinoma of testis with other germ cell elements (diagnosis)
C2057597|choriocarcinoma of testis with other germ cell elements
C2057597|testicular choriocarcinoma combined with other germ cell elements
C2057494|teratocarcinoma of testis (diagnosis)
C2057494|teratocarcinoma of testis
C2057494|testicular teratocarcinoma
C0334517|Spermatocytic Seminoma
C0334517|Spermatocytoma
C0334517|Spermatocytic seminoma (morphologic abnormality)
C0334517|Testicular Spermatocytic Seminoma
C0279708|yolk sac tumor of testis (diagnosis)
C0279708|yolk sac tumor of testis
C0279708|Testicular yolk sac tumour
C0279708|Testicular yolk sac tumor
C0279708|testicle cancer, yolk sac tumor
C0279708|testicular cancer, yolk sac tumor
C0279708|testis cancer, yolk sac tumor
C0279708|yolk sac tumor of the testis
C0279708|yolk sac tumor, testicular
C0279708|Endodermal Sinus Neoplasm of Testis
C0279708|Endodermal Sinus Neoplasm of the Testis
C0279708|Endodermal Sinus Tumor of Testis
C0279708|Endodermal Sinus Tumor of the Testis
C0279708|Testicular Endodermal Sinus Neoplasm
C0279708|Testicular Endodermal Sinus Tumor
C0279708|Testicular Yolk Sac Neoplasm
C0279708|Yolk Sac Neoplasm of Testis
C0279708|Yolk Sac Neoplasm of the Testis
C1336720|malignant mixed germ cell tumor of testis (diagnosis)
C1336720|malignant mixed germ cell tumor of testis
C1336720|Testicular germ cell tumour mixed
C1336720|Testicular germ cell tumor mixed
C1336720|Mixed Germ Cell Neoplasm of Testis
C1336720|Mixed Germ Cell Neoplasm of the Testis
C1336720|Mixed Germ Cell Tumor of Testis
C1336720|Mixed Germ Cell Tumor of the Testis
C1336720|Testicular Germ Cell Tumor (Mixed)
C1336720|Testicular Mixed Germ Cell Neoplasm
C1336720|Testicular Mixed Germ Cell Tumor
C3646009|testicular malignant neoplasm secondary
C3646009|secondary malignant testicular neoplasm (diagnosis)
C3646009|secondary malignant testicular neoplasm
C3646010|primary malignant testicular neoplasm
C3646010|testicular malignant neoplasm primary
C3646010|primary malignant testicular neoplasm (diagnosis)
C2315963|testicular neoplasm malignant non-seminomatous
C2315963|Non-seminomatous malignant neoplasm of testis (diagnosis)
C2315963|Non-seminomatous malignant neoplasm of testis
C2315963|Non-seminomatous malignant neoplasm of testis (disorder)
C0346236|malignant neoplasm of ectopic testis
C0346236|malignant neoplasm of ectopic testis (diagnosis)
C0346236|malignant tumor of ectopic testis
C0346236|Cancer of ectopic testis
C0346236|Malignant tumour of ectopic testis
C0346236|Malignant tumor of ectopic testis (disorder)
C0346241|malignant neoplasm of tunica vaginalis (diagnosis)
C0346241|malignant neoplasm of tunica vaginalis
C0346241|malignant tumor of tunica vaginalis
C0346241|Malignant tumour of tunica vaginalis
C0346241|Malignant tumor of tunica vaginalis (disorder)
C0347003|Metastatic Neoplasm to the Testis
C0347003|Metastases to testicle
C0347003|Metastatic Malignant Neoplasm in the Testis
C0347003|Metastatic Malignant Neoplasm to the Testis
C0347003|Metastasis to testis
C0347003|Metastatic tumor to testis
C0347003|Metastatic tumour to testis
C0347003|Secondary malignant neoplasm of testis
C0347003|Metastatic malignant neoplasm to testis
C0347003|Secondary malignant neoplasm of testis (disorder)
C0347003|Metastatic malignant neoplasm to testis, NOS
C0347003|Secondary malignant neoplasm of testis, NOS
C0347003|Metastatic Tumor to the Testis
C1304869|Primary malignant neoplasm of testis (disorder)
C1304869|Primary malignant neoplasm of testis
C0153596|Malig neo testis NEC
C0153596|Malignant neoplasm of other and unspecified testis
C0153596|Malignant neoplasm of testis, other and unspecified
C0852641|Testis cancer (excl germ cell)
C0852641|Testis cancer (excluding germ cell)
C1387440|seminoma; anaplastic, unspecified site
C1387440|anaplastic; seminoma, unspecified site
C1388417|malignant; androblastoma, unspecified site, male
C1388417|malignant; arrhenoblastoma, unspecified site, male
C1388417|androblastoma; malignant, unspecified site, male
C1388417|arrhenoblastoma; malignant, unspecified site, male
C1391898|carcinoma; chorion, unspecified site, male
C1391898|chorion; carcinoma, unspecified site, male
C1391920|carcinoma; Leydig cell, unspecified site, male
C1391920|Leydig cell; carcinoma, unspecified site, male
C1391943|carcinoma; Sertoli cell, unspecified site
C1391943|Sertoli cell; carcinoma, unspecified site
C1391944|carcinoma; Sertoli cell, unspecified site, male
C1391944|Sertoli cell; carcinoma, unspecified site, male
C1392523|choriocarcinoma; male
C1392523|choriocarcinoma; unspecified site, male
C1395770|tumor; yolk sac, unspecified site, male
C1395770|yolk sac; tumor, unspecified site, male
C1395936|dysgerminoma; unspecified site, male
C1396368|embryoma; malignant, testis
C1396368|malignant; embryoma, testis
C1396371|embryoma; testis
C1396371|testis; embryoma
C1396615|endodermal; sinus, tumor, unspecified site, male
C1396615|tumor; endodermal sinus, unspecified site, male
C1402881|Leydig cell; tumor, malignant, unspecified site, male
C1402881|tumor; Leydig cell, malignant, unspecified site, male
C0334528|Malignant Trophoblastic Teratoma
C0334528|trophoblastic malignant teratoma (diagnosis)
C0334528|trophoblastic malignant teratoma
C0334528|Malignant teratoma, trophoblastic
C0334528|Malignant teratoma, trophoblastic (morphologic abnormality)
C0334528|malignant; teratoma, trophoblastic, unspecified site
C0334528|teratoma; malignant, trophoblastic, unspecified site
C0014145|Endodermal Sinus Tumor
C0014145|Endodermal Sinus Tumors
C0014145|Tumor, Endodermal Sinus
C0014145|Tumor, Yolk Sac
C0014145|Tumors, Endodermal Sinus
C0014145|Tumors, Yolk Sac
C0014145|Yolk Sac Tumors
C0014145|yolk sac tumor (diagnosis)
C0014145|yolk sac tumor
C0014145|Yolk sac tumour site unspecified
C0014145|Endodermal Sinus Tumor [Disease/Finding]
C0014145|YOLK SAC TUMOR, MALIGNANT
C0014145|Yolk Sac Neoplasm
C0014145|Endodermal Sinus Neoplasm
C0014145|Yolk Sac Tumor Site Unspecified
C0014145|Endodermal sinus tumour site unspecified
C0014145|Endodermal sinus tumor site unspecified
C0014145|Polyvesicular vitelline tumor
C0014145|Orchioblastoma
C0014145|Embryonal carcinoma, infantile
C0014145|Endodermal sinus tumour
C0014145|Infantile embryonal carcinoma
C0014145|Polyvesicular vitelline tumour
C0014145|Yolk sac tumour
C0014145|Endodermal sinus tumor (morphologic abnormality)
C0014145|Hepatoid yolk sac tumor
C0014145|Hepatoid yolk sac tumour
C0014145|Yolk sac tumor (disorder)
C1405366|polyvesicular; tumor, unspecified site, male
C1405366|tumor; polyvesicular, unspecified site, male
C1409893|seminoma; unspecified site
C1409893|spermatocytoma; unspecified site
C1409698|seminoma; spermatocytic, unspecified site
C1409698|spermatocytic; seminoma, unspecified site
C0238451|TERATOMA, TESTICULAR
C0238451|testicular teratoma
C0238451|Teratoma of testis
C0238451|Teratoma of testis (disorder)
C0238451|Teratoma of testes
C0238451|teratoma of the testis
C0238451|testicle cancer, teratoma
C0238451|testicular cancer, teratoma
C0238451|testis cancer, teratoma
C0238451|teratoma; testis
C0238451|testis; teratoma
C0280256|stage, testicular cancer
C0280256|testicular cancer stage
C0279869|cellular diagnosis, testicular cancer
C0279869|testicular cancer cellular diagnosis
C1336711|Testicular Leukemia
C1515289|Malignant Testicular Sex Cord-Stromal Tumor
C2212316|mast cell sarcoma of testis (diagnosis)
C2212316|mast cell sarcoma of testis
C2057633|malignant histiocytosis of testis
C2057633|malignant histiocytosis of testis (diagnosis)
C0153597|Malignant neoplasm of penis and other male genital organs
C0153597|Malignant neoplasm of penis and other male genital organs (disorder)
C0153597|Malignant neoplasm of penis and other male genital organ NOS
C0153597|Malignant neoplasm of penis and other male genital organ NOS (disorder)
C0376358|Malignant neoplasm of prostate
C0376358|prostate cancer
C0376358|prostatic cancer
C0376358|Cancer of prostate
C0376358|Cancer, Prostate
C0376358|Cancers, Prostate
C0376358|Prostate Cancers
C0376358|Cancer, Prostatic
C0376358|Cancers, Prostatic
C0376358|Prostatic Cancers
C0376358|prostate cancer (diagnosis)
C0376358|malignant neoplasm of prostate gland (diagnosis)
C0376358|malignant neoplasm of prostate gland
C0376358|Ca prostate
C0376358|malignant tumor of prostate gland
C0376358|Malign neopl prostate
C0376358|Prostatic neoplasms malignant
C0376358|Malignant prostatic tumor
C0376358|Malignant tumour of prostate
C0376358|CA - Cancer of prostate
C0376358|Malignant tumor of prostate
C0376358|Malignant prostatic tumour
C0376358|Malignant tumor of prostate (disorder)
C0376358|Prostate--Cancer
C0376358|-- Prostate Cancer
C0376358|Prostate cancer NOS
C0376358|Cancer of the Prostate
C0376358|Malignant Neoplasm of the Prostate
C0376358|Malignant Prostate Neoplasm
C0376358|Malignant Prostate Tumor
C0376358|Malignant Tumor of the Prostate
C0376358|Neoplasm malig;prostate
C0376358|malignant neosplasm of the prostate
C0497581|Malignant neoplasm of other and unspecified male genital organs
C0497581|Other male genital malignant neoplasm
C0497581|Cancer of other male genital organs
C0497581|Malignant neoplasm of other male genital organ
C0497581|Malignant neoplasm of other male genital organ NOS (disorder)
C0497581|Malignant neoplasm of other male genital organ NOS
C0497581|Malignant neoplasm of other male genital organ (disorder)
C0153601|Malignant neoplasm of penis
C0153601|Malignant neoplasm of penis, unspecified
C0153601|Penis, unspecified
C0153601|malignant neoplasm of penis (diagnosis)
C0153601|malignant penile neoplasm
C0153601|Cancer, Penile
C0153601|Cancers, Penile
C0153601|Penile Cancers
C0153601|Cancers, Penis
C0153601|Penis Cancers
C0153601|malignant tumor of penis
C0153601|penile cancer
C0153601|Malig neo penis NOS
C0153601|Cancer, Penis
C0153601|Penile neoplasms malignant
C0153601|Ca penis (disorder)
C0153601|Malignant neoplasm of penis, part unspecified (disorder)
C0153601|Ca penis
C0153601|Malignant neoplasm of penis, part unspecified
C0153601|Cancer of penis
C0153601|Penile Ca
C0153601|CA - Cancer of penis
C0153601|Malignant tumour of penis
C0153601|Penis--Cancer
C0153601|Penile malignant neoplasm NOS
C0153601|Penile malignant neoplasm
C0153601|Penis Cancer
C0153601|Cancer of the Penis
C0153601|Malignant tumor of penis (disorder)
C0153601|Malignant neoplasm of penis, NOS
C0153601|Malignant Neoplasm of the Penis
C0153601|Malignant Penile Tumor
C0153601|Malignant Tumor of the Penis
C0153606|Malignant neoplasm of male genital organ, unspecified
C0153606|Male genital organ, unspecified
C0153606|malignant tumor of male genital organ
C0153606|Malignant neoplasm of male genital organ
C0153606|male genital cancer
C0153606|male genital cancer (diagnosis)
C0153606|Malignant neoplasms of male genital organs
C0153606|malignant tumor of male genitalia
C0153606|Mal neo male genital NOS
C0153606|Cancer of male genital organs
C0153606|Malignant neoplasms of male genital organs (C60-C63)
C0153606|malignant neoplasm of male genitalia
C0153606|malignant neoplasm of the male genital organs (diagnosis)
C0153606|malignant neoplasm of the male genital organs
C0153606|malignant neoplasm of male genital organs
C0153606|Genital cancer male
C0153606|[X]Malignant neoplasm of male genital organs (disorder)
C0153606|[X]Malignant neoplasm of male genital organ, unspecified (disorder)
C0153606|[X]Malignant neoplasm of male genital organ, unspecified
C0153606|[X]Malignant neoplasm of male genital organs
C0153606|Male reprod. system cancer, NOS
C0153606|Male reproductive system cancer, NOS
C0153606|Malignant neoplasm of male genital organ, site unspecified
C0153606|Malignant tumour of male genital organ
C0153606|Malignant tumor of male genital organ (disorder)
C0153606|Malignant neoplasm of male genital organ, NOS
C0153606|Malignant Male Reproductive System Neoplasm
C0153606|Malignant Male Reproductive System Tumor
C0153606|Malignant Neoplasm of Male Reproductive System
C0153606|Malignant Neoplasm of the Male Reproductive System
C0153606|Malignant Tumor of Male Reproductive System
C0153606|Malignant Tumor of the Male Reproductive System
C0153606|Malignant neoplasm of male genital organ or tract NOS
C0153606|Neoplasm malig;genital sys;M
C0153606|malignant neosplasm of the male genital system
C2217869|male genital neoplasm malignant small cell type
C2217869|malignant small cell neoplasm of male genitalia
C2217869|malignant small cell neoplasm of male genitalia (diagnosis)
C2011384|giant cell type neoplasm of male genitalia (diagnosis)
C2011384|giant cell type neoplasm of male genitalia
C2018667|spindle cell type neoplasm of male genitalia
C2018667|spindle cell type neoplasm of male genitalia (diagnosis)
C2075627|clear cell type neoplasm of male genitalia
C2075627|clear cell type neoplasm of male genitalia (diagnosis)
C2007032|carcinoma of male genitalia
C2007032|carcinoma of male genitalia (diagnosis)
C2215312|adenocarcinoma of male genitalia
C2215312|adenocarcinoma of male genitalia (diagnosis)
C2219527|sarcoma of male genitalia (diagnosis)
C2219527|sarcoma of male genitalia
C2230877|fibrosarcoma of male genitalia (diagnosis)
C2230877|fibrosarcoma of male genitalia
C2184067|liposarcoma of male genitalia (diagnosis)
C2184067|liposarcoma of male genitalia
C2230880|myosarcoma of male genitalia
C2230880|myosarcoma of male genitalia (diagnosis)
C2007077|carcinosarcoma of male genitalia
C2007077|carcinosarcoma of male genitalia (diagnosis)
C2216612|malignant mesenchymoma of male genitalia
C2216612|malignant mesenchymoma of male genitalia (diagnosis)
C2216469|marginal zone B-cell lymphoma of male genitalia
C2216469|marginal zone B-cell lymphoma of male genitalia (diagnosis)
C2216535|malignant fibrous histiocytoma of male genitalia
C2216535|malignant fibrous histiocytoma of male genitalia (diagnosis)
C2230882|Mullerian mixed tumor of male genitalia (diagnosis)
C2230882|Mullerian mixed tumor of male genitalia
C2216616|malignant mesodermal mixed tumor of male genitalia (diagnosis)
C2216616|malignant mesodermal mixed tumor of male genitalia
C2188071|undifferentiated carcinoma of male genitalia (diagnosis)
C2188071|undifferentiated carcinoma of male genitalia
C2230874|basaloid carcinoma of male genitalia
C2230874|basaloid carcinoma of male genitalia (diagnosis)
C2230874|basaloid carcinoma of male genital tract
C2216459|fibroblastic liposarcoma of male genitalia (diagnosis)
C2216459|fibroblastic liposarcoma of male genitalia
C1306367|Primary malignant neoplasm of male genital organ (diagnosis)
C1306367|Primary malignant neoplasm of male genital organ
C1306367|male genital malignant neoplasm primary
C1306367|Primary malignant neoplasm of male genital organ (disorder)
C0348369|Malignant neoplasm overlapping male genital organ site
C0348369|Overlapping lesion of male genital organs
C0348369|Malignant neoplasm of overlapping sites of male genital organs
C0348369|Malignant neoplasm of ovrlp sites of male genital organs
C0348369|malignant neoplasm of overlapping sites of male genital organs (diagnosis)
C0348369|male genital neoplasm malignant overlapping sites
C0348369|Malignant neoplasm, overlapping lesion of male genital organs
C0348369|[X]Malignant neoplasm of overlapping lesion of male genital organs
C0348369|[X]Malignant neoplasm of overlapping lesion of male genital organs (disorder)
C0348369|Malignant neoplasm, overlapping lesion of male genital organs (disorder)
C0348369|Overlapping malignant neoplasm of male genital organs (disorder)
C0348369|Overlapping malignant neoplasm of male genital organs
C0686232|Secondary malignant neoplasm of vas deferens
C0686232|spermatic cord neoplasm malignant vas deferens secondary
C0686232|Secondary malignant neoplasm of vas deferens (diagnosis)
C0686232|Metastatic malignant neoplasm to vas deferens
C0686232|Secondary malignant neoplasm of vas deferens (disorder)
C0864963|Malignant neoplasm of skin of scrotum
C0864963|Cancer of scrotal skin
C0864963|Malignant neoplasm of skin of scrotum (disorder)
C0864963|scrotal neoplasm malignant of skin
C0864963|malignant neoplasm of scrotal skin
C0864963|malignant neoplasm of scrotal skin (diagnosis)
C0346225|Malignant neoplasm of skin of penis NOS
C0346225|malignant neoplasm of skin of penis
C0346225|malignant neoplasm of skin of penis (diagnosis)
C0346225|penile neoplasm malignant of skin
C0346225|Cancer of penile skin
C0346225|Malignant tumor of penile skin
C0346225|Malignant tumor of skin of penis
C0346225|Malignant tumour of penile skin
C0346225|Malignant tumour of skin of penis
C0346225|Malignant tumor of skin of penis (disorder)
C0153602|Epididymis
C0153602|Malignant neoplasm of epididymis
C0153602|Malignant tumor of epididymis
C0153602|malignant neoplasm of epididymis (diagnosis)
C0153602|cancer of epididymis
C0153602|Malig neo epididymis
C0153602|Epididymal cancer
C0153602|Malignant epididymal neoplasm NOS
C0153602|Malignant tumour of epididymis
C0153602|Malignant tumor of epididymis (disorder)
C0153602|Malignant Epididymal Neoplasm
C0153602|Malignant Epididymal Tumor
C0153602|Malignant Neoplasm of the Epididymis
C0153602|Malignant Tumor of the Epididymis
C0346216|malignant neoplasm of seminal vesicle (diagnosis)
C0346216|malignant neoplasm of seminal vesicle
C0346216|malignant tumor of seminal vesicle
C0346216|Malignant tumour of seminal vesicle
C0346216|Malignant tumor of seminal vesicle (disorder)
C0153603|Malignant neoplasm of spermatic cord
C0153603|Spermatic cord
C0153603|malignant neoplasm of spermatic cord (diagnosis)
C0153603|malignant tumor of spermatic cord
C0153603|Mal neo spermatic cord
C0153603|Spermatic cord Ca
C0153603|Malignant tumour of spermatic cord
C0153603|Malignant tumor of spermatic cord (disorder)
C0153603|Malignant Neoplasm of the Spermatic Cord
C0153603|Malignant Spermatic Cord Neoplasm
C0153603|Malignant Spermatic Cord Tumor
C0153603|Malignant Tumor of the Spermatic Cord
C0347000|male genital malignant neoplasm secondary
C0347000|Secondary malignant neoplasm of male genital organ (diagnosis)
C0347000|Secondary malignant neoplasm of male genital organ
C0347000|Cancer metastatic to male genital organ
C0347000|Cancer metastatic to male genitalia
C0347000|Metastasis to male genital organ
C0347000|Metastatic malignant neoplasm to male genital organ
C0347000|Secondary malignant neoplasm of male genital organ (disorder)
C0347000|Metastatic malignant neoplasm to male genital organ, NOS
C0347000|Secondary malignant neoplasm of male genital organ, NOS
C0348368|Malignant neoplasm of other specified male genital organs
C0348368|Other specified male genital organs
C0348368|[X]Malignant neoplasm of other specified male genital organs
C0348368|[X]Malignant neoplasm of other specified male genital organs (disorder)
C1398495|genital organs; melanoma, male (external)
C1398495|melanoma; genital organs, male (external)
C0863024|Adenocarcinoma of the rete testis
C0863024|Adenocarcinoma of Rete Testis
C0863024|Rete Testis Adenocarcinoma
C1519233|Seminal Vesicle Adenocarcinoma
C1335705|Recurrent Male Reproductive System Carcinoma
C1335705|Recurrent Male Reproductive System Cancer
C0746787|Malignant neoplasm of neck
C0746787|neck cancer
C0746787|malignant neoplasm of neck (diagnosis)
C0746787|Malignant neoplasm of neck NOS
C0746787|Malignant neoplasm of neck NOS (disorder)
C0746787|Neck--Cancer
C0746787|Cancer of Neck
C0746787|Cancer of the Neck
C0746787|Malignant tumor of neck
C0746787|Malignant tumour of neck
C0746787|Malignant tumor of neck (disorder)
C0746787|Malignant neoplasm of neck, NOS
C0746787|Malignant Neck Neoplasm
C0746787|Malignant Neck Tumor
C0746787|Malignant Neoplasm of the Neck
C0746787|Malignant Tumor of the Neck
C2711842|Adenocarcinoma of head and neck
C2711842|Adenocarcinoma of head and neck (disorder)
C2711842|Adenocarcinoma of head and neck (diagnosis)
C2711842|malignant neoplasm of ill-defined site head and neck adenocarcinoma
C1263914|Primary malignant neoplasm of peripheral nerves of face (diagnosis)
C1263914|Primary malignant neoplasm of peripheral nerves of face
C1263914|neoplasm - pns malignant face primary
C1263914|Primary malignant neoplasm of peripheral nerves of face (disorder)
C0153744|Hodgkin's sarcoma of lymph nodes of head, face, and neck
C0153744|Hodgkins sarcoma head
C0153744|Hodgkin sarcoma of lymph nodes of head, face and neck
C0153744|Hodgkin sarcoma of lymph nodes of head, face AND/OR neck
C0153744|Hodgkin's sarcoma involving lymph nodes of head, face, and neck
C0153744|Hodgkin's sarcoma, lymph nodes of head, face, and neck
C0153744|Hodgkin sarcoma of lymph nodes of head, face, or neck
C0153744|Hodgkin sarcoma of lymph nodes of head, face, or neck (diagnosis)
C0153744|Hodgkin's sarcoma of lymph nodes of head, face and neck
C0153744|Hodgkin's sarcoma of lymph nodes of head, face AND/OR neck (disorder)
C0153744|Hodgkin's sarcoma of lymph nodes of head, face AND/OR neck
C0153744|Hodgkin's sarcoma of lymph nodes of head, face and neck (disorder)
C0153744|Hodgkin's sarcoma involving lymph nodes of head, face and neck
C0587226|Secondary malignant neoplasm of tongue (disorder)
C0587226|Secondary malignant neoplasm of tongue
C0587226|Tongue cancer metastatic
C0587226|tongue neoplasm malignant secondary
C0587226|Secondary malignant neoplasm of tongue (diagnosis)
C0587226|Metastatic malignant neoplasm to tongue
C0587226|Metastatic malignant neoplasm to tongue, NOS
C0587226|Secondary malignant neoplasm of tongue, NOS
C0346931|malignant neoplasm of nasolacrimal duct
C0346931|malignant neoplasm of nasolacrimal duct (diagnosis)
C0346931|malignant tumor of nasolacrimal duct
C0346931|Malignant neoplasm of nasolacrimal duct (disorder)
C0153379|Malignant neoplasm of retromolar area
C0153379|Retromolar area
C0153379|malignant neoplasm of retromolar area (diagnosis)
C0153379|malignant retromolar area neoplasm
C0153379|malignant tumor of retromolar area
C0153379|Malig neo retromolar
C0153379|Malignant tumour of retromolar area
C0153379|Malignant tumor of retromolar area (disorder)
C0349031|Melanoma in situ of scalp and neck
C0349031|skin neoplasm melanoma in situ of scalp and neck
C0349031|melanoma in situ of scalp and neck (diagnosis)
C0349031|Melanoma in situ of scalp and neck (disorder)
C0220636|Malignant neoplasm of salivary gland
C0220636|Malignant neoplasm of salivary gland duct
C0220636|malignant neoplasm of salivary gland (diagnosis)
C0220636|Cancers, Salivary Gland
C0220636|Salivary Gland Cancers
C0220636|malignant tumor of salivary gland
C0220636|Mal neo salivary NOS
C0220636|Cancer, Salivary Gland
C0220636|Salivary gland neoplasms malignant
C0220636|Salivary Gland Cancer
C0220636|Salivary glands--Cancer
C0220636|Salivary gland cancer NOS
C0220636|Malignant salivary gland cancer
C0220636|Malignant salivary gland neoplasm
C0220636|Malignant neoplasm of salivary gland, unspecified
C0220636|Cancer of the Salivary Gland
C0220636|CA - Cancer of salivary gland
C0220636|Cancer of salivary gland
C0220636|Malignant tumour of salivary gland
C0220636|Malignant tumor of salivary gland (disorder)
C0220636|Malignant Neoplasm of the Salivary Gland
C0220636|Malignant Salivary Gland Tumor
C0220636|Malignant Tumor of the Salivary Gland
C0220636|Malignant neoplasm of salivary gland NOS
C0684535|bone neoplasm, malignant - face secondary
C0684535|Secondary malignant neoplasm of bone of face
C0684535|Secondary malignant neoplasm of bone of face (diagnosis)
C0684535|Metastatic malignant neoplasm to bone of face
C0684535|Secondary malignant neoplasm of bone of face (disorder)
C0684535|Metastatic malignant neoplasm to bone of face, NOS
C0684535|Secondary malignant neoplasm of bone of face, NOS
C0585362|malignant squamous cell neoplasm of oral cavity (diagnosis)
C0585362|malignant squamous cell neoplasm of oral cavity
C0585362|Squamous cell carcinoma of the oral cavity
C0585362|Squamous cell carcinoma of mouth
C0585362|Squamous cell carcinoma of mouth (disorder)
C0585362|Mouth SCC
C0585362|Mouth Squamous Cell Carcinoma
C0585362|Oral Cavity SCC
C0585362|Oral Cavity Squamous Cell Carcinoma
C0585362|SCC of Mouth
C0585362|SCC of Oral Cavity
C0585362|SCC of the Mouth
C0585362|SCC of the Oral Cavity
C0585362|Squamous Cell Carcinoma of Oral Cavity
C0585362|Squamous Cell Carcinoma of the Mouth
C0686635|Secondary and unspecified malignant neoplasm of submental lymph nodes (disorder)
C0686635|Secondary and unspecified malignant neoplasm of submental lymph nodes
C0686635|lymph node neoplasm malignant secondary face submental
C0686635|Secondary malignant neoplasm of submental lymph nodes
C0686635|Secondary malignant neoplasm of submental lymph nodes (diagnosis)
C0686635|Metastatic malignant neoplasm to submental lymph nodes
C0686635|Secondary malignant neoplasm of submental lymph nodes (disorder)
C0153802|Mycosis fungoides of lymph nodes of head, face, and neck
C0153802|mycosis fungoides of head, face, and neck
C0153802|mycosis fungoides of head, face, and neck (diagnosis)
C0153802|Mycosis fungoides head
C0153802|Mycosis fungoides, lymph nodes of head, face, and neck
C0153802|Mycosis fungoides involving lymph nodes of head, face, and neck
C0153802|Mycosis fungoides of the lymph nodes of head, face and neck (disorder)
C0153802|Mycosis fungoides of the lymph nodes of head, face and neck
C0153802|Mycosis fungoides of lymph nodes of head, face AND/OR neck (disorder)
C0153802|Mycosis fungoides of lymph nodes of head, face AND/OR neck
C0153802|Mycosis fungoides involving lymph nodes of head, face and neck
C0684747|malignant neoplasm of muscle of head primary
C0684747|Primary malignant neoplasm of muscle of head (diagnosis)
C0684747|Primary malignant neoplasm of muscle of head
C0684747|Primary malignant neoplasm of muscle of head (disorder)
C0339112|Bowen disease of eyelid
C0339112|Bowen's disease of eyelid
C0339112|Bowen's disease of eyelid (diagnosis)
C0339112|Bowen's disease of eyelid (disorder)
C0686633|Secondary and unspecified malignant neoplasm of submandibular lymph nodes (disorder)
C0686633|Secondary and unspecified malignant neoplasm of submandibular lymph nodes
C0686633|Secondary malignant neoplasm of submandibular lymph nodes
C0686633|Secondary malignant neoplasm of submandibular lymph nodes (diagnosis)
C0686633|lymph node neoplasm malignant secondary neck submandibular
C0686633|Metastatic malignant neoplasm to submandibular lymph nodes
C0686633|Secondary malignant neoplasm of submandibular lymph nodes (disorder)
C0684530|Secondary malignant neoplasm of sphenoid bone
C0684530|Secondary malignant neoplasm of sphenoid bone (diagnosis)
C0684530|bone neoplasm, malignant - skull sphenoid bone secondary
C0684530|Metastatic malignant neoplasm to sphenoid bone
C0684530|Secondary malignant neoplasm of sphenoid bone (disorder)
C0153712|Burkitt's lymphoma of lymph nodes of head, face, and neck (diagnosis)
C0153712|Burkitt's lymphoma of head, face, and neck
C0153712|Burkitt's lymphoma of lymph nodes of head, face, and neck
C0153712|Burkitt's tumor head
C0153712|Burkitt lymphoma of lymph nodes of head, face and neck
C0153712|Burkitt lymphoma, lymph nodes of head, face, and neck
C0153712|Burkitt's tumor or lymphoma, lymph nodes of head, face, and neck
C0153712|Burkitt's tumor or lymphoma involving lymph nodes of head, face, and neck
C0153712|Burkitt's tumour or lymphoma involving lymph nodes of head, face, and neck
C0153712|Burkitt's lymphoma of lymph nodes of head, face and neck
C0153712|Burkitt's lymphoma of lymph nodes of head, face and neck (disorder)
C0153712|Burkitt's tumor or lymphoma involving lymph nodes of head, face and neck
C0686010|secondary malignant neoplasm of oral cavity
C0686010|oral cavity malignant neoplasm secondary
C0686010|secondary malignant neoplasm of oral cavity (diagnosis)
C0686010|Metastatic malignant neoplasm to mouth
C0686010|Secondary malignant neoplasm of mouth (disorder)
C0686010|Secondary malignant neoplasm of mouth
C0686010|Metastatic malignant neoplasm to mouth, NOS
C0686010|Secondary malignant neoplasm of mouth, NOS
C0563210|Squamous cell carcinoma of skin of cheek
C0563210|skin neoplasm face malignant squamous cell carcinoma cheek
C0563210|Squamous cell carcinoma of skin of cheek (diagnosis)
C0563210|Squamous cell carcinoma of skin of cheek (disorder)
C0684922|Secondary malignant neoplasm of upper respiratory tract
C0684922|Secondary malignant neoplasm of upper respiratory tract (diagnosis)
C0684922|malignant neoplasm upper respiratory tract secondary
C0684922|Metastatic malignant neoplasm to upper respiratory tract
C0684922|Secondary malignant neoplasm of upper respiratory tract (disorder)
C0684922|Metastatic malignant neoplasm to upper respiratory tract, NOS
C0684922|Secondary malignant neoplasm of upper respiratory tract, NOS
C1306049|hypopharyngeal neoplasm malignant postcricoid region primary
C1306049|Primary malignant neoplasm of postcricoid region
C1306049|Primary malignant neoplasm of postcricoid region (diagnosis)
C1306049|Primary malignant neoplasm of postcricoid region (disorder)
C0153728|Hodgkin's paragranuloma of lymph nodes of head, face, and neck
C0153728|Hodgkins paragran head
C0153728|Hodgkin paragranuloma of lymph nodes of head, face AND/OR neck
C0153728|Hodgkin's paragranuloma, lymph nodes of head, face, and neck
C0153728|Hodgkin's paragranuloma involving lymph nodes of head, face, and neck
C0153728|Hodgkin's paragranuloma of lymph nodes of head, face, and neck (disorder)
C0153728|Hodgkin disease paragranuloma - head, face, & neck
C0153728|Hodgkin paragranuloma of lymph nodes of head, face, & neck (diagnosis)
C0153728|Hodgkin paragranuloma of lymph nodes of head, face, & neck
C0153728|Hodgkin's paragranuloma of lymph nodes of head, face AND/OR neck (disorder)
C0153728|Hodgkin's paragranuloma of lymph nodes of head, face AND/OR neck
C0153728|Hodgkin's paragranuloma involving lymph nodes of head, face and neck
C0686024|Secondary malignant neoplasm of palate
C0686024|Secondary malignant neoplasm of palate (diagnosis)
C0686024|palate neoplasm malignant secondary
C0686024|Metastatic malignant neoplasm to palate
C0686024|Secondary malignant neoplasm of palate (disorder)
C0686024|Metastatic malignant neoplasm to palate, NOS
C0686024|Secondary malignant neoplasm of palate, NOS
C0686492|Secondary malignant neoplasm of mastoid air cells (diagnosis)
C0686492|Secondary malignant neoplasm of mastoid air cells
C0686492|bone neoplasm, malignant - skull and face, mastoid air cells secondary
C0686492|Metastatic malignant neoplasm to mastoid air cells
C0686492|Secondary malignant neoplasm of mastoid air cells (disorder)
C1304846|malignant neoplasm of neck primary
C1304846|Primary malignant neoplasm of neck
C1304846|Primary malignant neoplasm of neck (diagnosis)
C1304846|Primary malignant neoplasm of neck (disorder)
C0346980|secondary malignant skin neoplasm of head (diagnosis)
C0346980|skin neoplasm head secondary
C0346980|secondary malignant skin neoplasm of head
C0346980|Secondary malignant neoplasm of skin of head
C0346980|Secondary malignant neoplasm of skin of head (disorder)
C0496755|Malignant neoplasm of tip and lateral border of tongue
C0496755|Border of tongue
C0496755|Malignant neoplasm of border of tongue
C0496755|malignant neoplasm of tip and lateral border of tongue (diagnosis)
C0496755|malignant tumor of tip and lateral border of tongue
C0496755|Mal neo tip/lat tongue
C0496755|Malignant neoplasm of tip AND/OR lateral border of tongue
C0496755|tongue neoplasm malignant border
C0496755|malignant neoplasm of border of tongue (diagnosis)
C0496755|Malignant neoplasm of tongue, tip and lateral border
C0496755|Malignant neoplasm of border of tongue (disorder)
C0496755|Malignant neoplasm of tongue, tip and lateral border (disorder)
C0685133|Secondary malignant neoplasm of blood vessel of face
C0685133|Secondary malignant neoplasm of blood vessel of face (diagnosis)
C0685133|neoplasm - soft tissue types blood vessel malignant of face secondary
C0685133|Metastatic malignant neoplasm to blood vessel of face
C0685133|Secondary malignant neoplasm of blood vessel of face (disorder)
C0153644|MALIGNANT CRANIAL NERVE NEOPL
C0153644|CRANIAL NERVE NEOPL MALIGNANT
C0153644|NEOPL CRANIAL NERVE MALIGNANT
C0153644|Malignant neoplasm of cranial nerve
C0153644|malignant neoplasm of cranial nerve (diagnosis)
C0153644|malignant tumor of cranial nerve
C0153644|Mal neo cranial nerves
C0153644|Malignant neoplasm of cranial nerve NOS
C0153644|Malignant neoplasm of cranial nerves NOS
C0153644|Malignant neoplasm of cranial nerves NOS (disorder)
C0153644|Malignant neoplasm of cranial nerves
C0153644|Malignant cranial nerve neoplasm NOS
C0153644|Malignant cranial nerve neoplasm
C0153644|Tumors, Cranial Nerve, Malignant
C0153644|Malignant Cranial Nerve Tumors
C0153644|Malignant Cranial Nerve Neoplasms
C0153644|Neoplasms, Cranial Nerve, Malignant
C0153644|Cranial Nerve Tumors, Malignant
C0153644|Cranial Nerve Neoplasms, Malignant
C0153644|Malignant tumour of cranial nerve
C0153644|Malignant tumor of cranial nerve (disorder)
C0153644|Malignant neoplasm of cranial nerve, NOS
C0153644|Cranial Nerve Neoplasm, Malignant
C0153644|Malignant Cranial Nerve Tumor
C0153644|Malignant Neoplasm of the Cranial Nerve
C0153644|Malignant Tumor of the Cranial Nerve
C0686408|Secondary malignant neoplasm of cranial nerve
C0686408|Secondary malignant neoplasm of cranial nerve (diagnosis)
C0686408|cranial nerve neoplasm malignant secondary
C0686408|Metastatic malignant neoplasm to cranial nerve
C0686408|Secondary malignant neoplasm of cranial nerve (disorder)
C0686408|Metastatic malignant neoplasm to cranial nerve, NOS
C0686408|Secondary malignant neoplasm of cranial nerve, NOS
C0153696|Reticulosarcoma head
C0153696|Reticulosarcoma, lymph nodes of head, face, and neck
C0153696|Reticulosarcoma involving lymph nodes of head, face, and neck
C0153696|Reticulosarcoma of lymph nodes of head, face, and neck (disorder)
C0153696|Reticulosarcoma of lymph nodes of head, face, and neck
C0153696|Reticulosarcoma of lymph nodes of head, face and neck
C0153696|Reticulosarcoma of lymph nodes of head, face and neck (disorder)
C0153696|Reticulosarcoma involving lymph nodes of head, face and neck
C0684941|Secondary malignant neoplasm of accessory sinus (diagnosis)
C0684941|Secondary malignant neoplasm of accessory sinus
C0684941|accessory sinus neoplasm malignant secondary
C0684941|Metastatic malignant neoplasm to accessory sinus
C0684941|Secondary malignant neoplasm of accessory sinus (disorder)
C0684941|Metastatic malignant neoplasm to accessory sinus, NOS
C0684941|Secondary malignant neoplasm of accessory sinus, NOS
C0686623|Secondary malignant neoplasm of lymph nodes of face
C0686623|lymph node neoplasm malignant secondary face
C0686623|Secondary malignant neoplasm of lymph nodes of face (diagnosis)
C0686623|Cancer metastatic to lymph nodes of face
C0686623|Metastatic malignant neoplasm to lymph nodes of face
C0686623|Secondary malignant neoplasm of lymph nodes of face (disorder)
C0686623|Metastatic malignant neoplasm to lymph nodes of face, NOS
C0686623|Secondary malignant neoplasm of lymph nodes of face, NOS
C0685136|Secondary malignant neoplasm of blood vessel of neck
C0685136|neoplasm - soft tissue types blood vessel malignant of neck secondary
C0685136|Secondary malignant neoplasm of blood vessel of neck (diagnosis)
C0685136|Metastatic malignant neoplasm to blood vessel of neck
C0685136|Secondary malignant neoplasm of blood vessel of neck (disorder)
C0345614|Malignant neoplasm of minor salivary gland
C0345614|malignant neoplasm of minor salivary gland (diagnosis)
C0345614|malignant tumor of minor salivary gland
C0345614|malignant salivary gland neoplasm minor (diagnosis)
C0345614|malignant salivary gland neoplasm minor
C0345614|Malignant tumour of minor salivary gland
C0345614|Malignant tumor of minor salivary gland (disorder)
C0345614|Malignant Minor Salivary Gland Neoplasm
C0345614|Malignant Minor Salivary Gland Tumor
C0345614|Malignant Neoplasm of the Minor Salivary Gland
C0345614|Malignant Tumor of the Minor Salivary Gland
C0686608|oropharyngeal neoplasm tonsil malignant secondary
C0686608|secondary malignant neoplasm of of tonsil
C0686608|secondary malignant neoplasm of of tonsil (diagnosis)
C0686608|Metastatic malignant neoplasm to palatine tonsil
C0686608|Metastatic malignant neoplasm to tonsil
C0686608|Secondary malignant neoplasm of palatine tonsil
C0686608|Secondary malignant neoplasm of tonsil
C0686608|Secondary malignant neoplasm of tonsil (disorder)
C0346575|Malignant tumour posterior margin nasal septum and choanae
C0346575|Malignant tumor posterior margin nasal septum and choanae (disorder)
C0346575|Malignant neoplasm of posterior margin of nasal septum and choanae
C0346575|Malignant tumor posterior margin nasal septum and choanae
C0346575|nasal cavity neoplasm malignant of posterior margin of septum and choanae
C0346575|malignant neoplasm of posterior margin of nasal septum and choanae (diagnosis)
C0346575|Malignant tumor of posterior margin of nasal septum and choanae
C0346575|Malignant tumour of posterior margin of nasal septum and choanae
C0346575|Malignant tumor of posterior margin of nasal septum and choanae (disorder)
C0346726|Malignant neoplasm of skin of ear and external auricular canal
C0346726|Skin of ear and external auricular canal
C0346726|Malignant neoplasm of skin of ear and external auditory canal
C0346726|Malignant neoplasm of skin of ear and external auditory canal (disorder)
C0346726|Malignant neoplasm of skin of ear and external auricular canal (disorder)
C0346726|Malignant neoplasm of skin of ear and external auricular canal NOS (disorder)
C0346726|Malignant neoplasm of skin of ear and external auricular canal NOS
C0346726|malignant neoplasm of skin of external ear and auditory canal (diagnosis)
C0346726|malignant neoplasm of skin of external ear and auditory canal
C0346726|skin neoplasm external ear malignant and auditory canal
C0685135|Malignant neoplasm of blood vessel of neck
C0685135|neoplasm - soft tissue types blood vessel malignant of neck primary
C0685135|Primary malignant neoplasm of blood vessel of neck
C0685135|Primary malignant neoplasm of blood vessel of neck (diagnosis)
C0685135|Primary malignant neoplasm of blood vessel of neck (disorder)
C0346323|Optic nerve
C0346323|Malignant neoplasm of optic nerve
C0346323|Malignant tumor of optic nerve
C0346323|MALIGNANT OPTIC NERVE NEOPL
C0346323|Malignant tumour of optic nerve
C0346323|Malignant tumour of optic nerve (disorder)
C0346323|Malignant Optic Nerve Tumor
C0346323|Tumor, Optic Nerve, Malignant
C0346323|Optic Nerve Tumor, Malignant
C0346323|Tumor, Malignant, Optic Nerve
C0346323|Malignant Optic Nerve Neoplasm
C0346323|Malignant tumor of optic nerve (disorder)
C0153654|Malignant neoplasm of pituitary gland and craniopharyngeal duct
C0153654|Malig neo pituitary
C0153654|Malignant neoplasm of pituitary gland or craniopharyngeal duct NOS (disorder)
C0153654|Malignant neoplasm of pituitary gland or craniopharyngeal duct NOS
C0153654|malignant neoplasm of pituitary gland and craniopharyngeal duct (diagnosis)
C0153654|Malignant neoplasm of pituitary gland and craniopharyngeal duct (disorder)
C0685130|Secondary malignant neoplasm of blood vessel of head
C0685130|Secondary malignant neoplasm of blood vessel of head (diagnosis)
C0685130|neoplasm - soft tissue types blood vessel malignant of head secondary
C0685130|Metastatic malignant neoplasm to blood vessel of head
C0685130|Secondary malignant neoplasm of blood vessel of head (disorder)
C0496788|Middle ear
C0496788|Malignant neoplasm of middle ear
C0496788|auditory neoplasm malignant of middle ear
C0496788|malignant neoplasm of middle ear (diagnosis)
C0496788|Malignant middle ear neoplasm NOS
C0496788|Malignant middle ear neoplasm
C0496788|Malignant tumor of middle ear
C0496788|Malignant tumour of middle ear
C0496788|Malignant tumor of middle ear (disorder)
C0496788|Malignant Middle Ear Tumor
C0496788|Malignant Neoplasm of the Middle Ear
C0496788|Malignant Tumor of the Middle Ear
C0684689|soft tissue neoplasm head malignant secondary
C0684689|secondary malignant soft tissue neoplasm of head
C0684689|secondary malignant soft tissue neoplasm of head (diagnosis)
C0684689|Metastatic malignant neoplasm to soft tissues of head
C0684689|Secondary malignant neoplasm of soft tissues of head
C0684689|Secondary malignant neoplasm of soft tissues of head (disorder)
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance of lymph nodes of head, face, and neck
C0153752|Hodg lymph-histio head
C0153752|Hodgkin disease, lymphocytic-histiocytic predominance of lymph nodes of head, face AND/OR neck
C0153752|Hodgkin disease, lymphocytic-histiocytic predominance of lymph nodes of head, face and neck
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance involving lymph nodes of head, face, and neck
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance, lymph nodes of head, face, and neck
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance of lymph nodes of head, face, or neck
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance of lymph nodes of head, face, and neck (diagnosis)
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance of lymph nodes of head, face and neck
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance of lymph nodes of head, face AND/OR neck (disorder)
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance of lymph nodes of head, face AND/OR neck
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance of lymph nodes of head, face and neck (disorder)
C0153752|Hodgkin's disease, lymphocytic-histiocytic predominance involving lymph nodes of head, face and neck
C0153688|Secondary malignant neoplasm of brain and spinal cord
C0153688|Sec mal neo brain/spine
C0153688|secondary malignant neoplasm brain and spinal cord
C0153688|secondary malignant neoplasm brain and spinal cord (diagnosis)
C0153688|Secondary malignant neoplasm of brain or spinal cord NOS (disorder)
C0153688|Secondary malignant neoplasm of brain or spinal cord NOS
C0153688|Secondary malignant neoplasm of brain and spinal cord (disorder)
C0685132|Malignant neoplasm of blood vessel of face
C0685132|Primary malignant neoplasm of blood vessel of face
C0685132|Primary malignant neoplasm of blood vessel of face (diagnosis)
C0685132|neoplasm - soft tissue types blood vessel malignant of face primary
C0685132|Primary malignant neoplasm of blood vessel of face (disorder)
C0684756|Secondary malignant neoplasm of muscle of neck (diagnosis)
C0684756|Secondary malignant neoplasm of muscle of neck
C0684756|malignant neoplasm of muscle of neck secondary
C0684756|Metastatic malignant neoplasm to muscle of neck
C0684756|Secondary malignant neoplasm of muscle of neck (disorder)
C0684692|secondary malignant soft tissue neoplasm of face
C0684692|soft tissue neoplasm face malignant secondary
C0684692|secondary malignant soft tissue neoplasm of face (diagnosis)
C0684692|Metastatic malignant neoplasm to soft tissues of face
C0684692|Secondary malignant neoplasm of soft tissues of face
C0684692|Secondary malignant neoplasm of soft tissues of face (disorder)
C0346124|Malignant neoplasm of soft tissues of head
C0346124|malignant soft tissue neoplasm of head
C0346124|malignant soft tissue neoplasm of head (diagnosis)
C0346124|soft tissue neoplasm head malignant
C0346124|Malignant tumor of soft tissue of head
C0346124|Malignant tumour of soft tissue of head
C0346124|Malignant neoplasm of soft tissue of head
C0346124|Malignant tumor of soft tissue of head (disorder)
C0349038|Malignant neoplasm overlapping nasopharynx site
C0349038|Overlapping lesion of nasopharynx
C0349038|Malignant neoplasm of overlapping sites of nasopharynx
C0349038|Malignant neoplasm, overlapping lesion of nasopharynx (disorder)
C0349038|Malignant neoplasm, overlapping lesion of nasopharynx
C0349038|Overlapping malignant neoplasm of nasopharyngeal wall
C0349038|Overlapping malignant neoplasm of nasopharynx (disorder)
C0349038|Overlapping malignant neoplasm of nasopharynx
C1263917|Primary malignant neoplasm of peripheral nerves of neck
C1263917|neoplasm - pns malignant neck primary
C1263917|Primary malignant neoplasm of peripheral nerves of neck (diagnosis)
C1263917|Primary malignant neoplasm of peripheral nerves of neck (disorder)
C0345628|Malignant neoplasm of mastoid air cells
C0345628|bone neoplasm, malignant - skull and face, mastoid air cells
C0345628|malignant neoplasm of mastoid air cells (diagnosis)
C0345628|Malignant tumor of mastoid air cells
C0345628|Malignant tumour of mastoid air cells
C0345628|Malignant tumor of mastoid air cells (disorder)
C0153704|Lymphosarcoma of lymph nodes of head, face AND/OR neck -RETIRED-
C0153704|Lymphosarcoma head
C0153704|Lymphosarcoma involving lymph nodes of head, face, and neck
C0153704|Lymphosarcoma, lymph nodes of head, face, and neck
C0153704|Lymphosarcoma of lymph nodes of head, face, and neck
C0153704|Lymphosarcoma of lymph nodes of head, face AND/OR neck (disorder)
C0153704|lymphosarcoma of head, face, and neck lymph nodes
C0153704|lymphosarcoma of lymph nodes of head, face, and neck (diagnosis)
C0153704|Lymphosarcoma of lymph nodes of head, face and neck
C0153704|Lymphosarcoma of lymph nodes of head, face and neck (disorder)
C0153704|Lymphosarcoma involving lymph nodes of head, face and neck
C0345586|oral cavity neoplasm malignant labial sulcus, lower
C0345586|malignant neoplasm of lower labial sulcus (diagnosis)
C0345586|malignant neoplasm of lower labial sulcus
C0345586|Malignant tumor of lower labial sulcus
C0345586|Malignant tumour of lower labial sulcus
C0345586|Malignant tumor of lower labial sulcus (disorder)
C0686641|Secondary and unspecified malignant neoplasm of infraclavicular lymph nodes
C0686641|Secondary and unspecified malignant neoplasm of infraclavicular lymph nodes (disorder)
C0686641|lymph node neoplasm malignant secondary neck infraclavicular
C0686641|Secondary malignant neoplasm of infraclavicular lymph nodes (diagnosis)
C0686641|Secondary malignant neoplasm of infraclavicular lymph nodes
C0686641|Metastatic malignant neoplasm to infraclavicular lymph nodes
C0686641|Secondary malignant neoplasm of infraclavicular lymph nodes (disorder)
C0153354|Malignant neoplasm of anterior two-thirds of tongue, part unspecified
C0153354|Anterior two-thirds of tongue, part unspecified
C0153354|Malignant neoplasm of anterior two-thirds of tongue
C0153354|malignant neoplasm of anterior two-thirds of tongue (diagnosis)
C0153354|malignant tumor of anterior two-thirds of tongue
C0153354|Mal neo ant 2/3 tongue
C0153354|Malignant neoplasm of mobile part of tongue NOS
C0153354|Malig neoplasm of anterior two-thirds of tongue, part unsp
C0153354|Malignant neoplasm of anterior 2/3 of tongue unspecified
C0153354|Malignant tumour of mobile part of tongue
C0153354|Malignant tumor of mobile part of tongue
C0153354|Malignant neoplasm of anterior 2/3 of tongue unspecified (disorder)
C0153354|Malignant tumour of anterior two-thirds of tongue
C0153354|Malignant tumor of anterior two-thirds of tongue (disorder)
C0153354|Malignant neoplasm of anterior two-thirds of tongue, NOS
C0153736|Hodgkin's granuloma of lymph nodes of head, face, and neck
C0153736|Hodgkins granulom head
C0153736|Hodgkin granuloma of lymph nodes of head, face and neck
C0153736|Hodgkin granuloma of lymph nodes of head, face AND/OR neck
C0153736|Hodgkin's granuloma, lymph nodes of head, face, and neck
C0153736|Hodgkin's granuloma involving lymph nodes of head, face, and neck
C0153736|Hodgkin disease granuloma - head, face, & neck
C0153736|Hodgkin granuloma of lymph nodes of head, face, & neck (diagnosis)
C0153736|Hodgkin granuloma of lymph nodes of head, face, & neck
C0153736|Hodgkin's granuloma of lymph nodes of head, face and neck
C0153736|Hodgkin's granuloma of lymph nodes of head, face AND/OR neck (disorder)
C0153736|Hodgkin's granuloma of lymph nodes of head, face AND/OR neck
C0153736|Hodgkin's granuloma of lymph nodes of head, face and neck (disorder)
C0153736|Hodgkin's granuloma involving lymph nodes of head, face and neck
C0684554|secondary malignant neoplasm of cervical vertebral column (diagnosis)
C0684554|secondary malignant neoplasm of cervical vertebral column
C0684554|bone neoplasm, malignant - vertebral column cervical secondary
C0684554|Metastatic malignant neoplasm to cervical vertebral column
C0684554|Secondary malignant neoplasm of cervical vertebral column (disorder)
C0347957|Connective and soft tissue of head, face and neck
C0347957|Malignant neoplasm of connective and soft tissue of head, face and neck
C0347957|Malig neoplm of conn and soft tissue of head, face and neck
C0347957|Malignant neoplasm of connective and soft tissue of head, face, and neck (disorder)
C0347957|Malignant neoplasm of connective and soft tissue of head, face, and neck
C0347957|Malignant neoplasm of connective and soft tissue of head, face and neck (disorder)
C0153768|Hodgkin's disease, mixed cellularity of lymph nodes of head, face, and neck
C0153768|Hodgkin's disease, mixed cellularity, involving lymph nodes of head, face, and neck.
C0153768|Hodgkins mix cell head
C0153768|Hodgkin disease, mixed cellularity of lymph nodes of head, face AND/OR neck
C0153768|Hodgkin disease, mixed cellularity of lymph nodes of head, face and neck
C0153768|Hodgkin's disease, mixed cellularity, lymph nodes of head, face, and neck
C0153768|Hodgkin's disease, mixed cellularity, involving lymph nodes of head, face, and neck
C0153768|mixed cellularity Hodgkin's lymphoma of lymph nodes of head, face, and neck
C0153768|Hodgkin's lymphoma mixed cellularity of head, face, and neck
C0153768|mixed cellularity Hodgkin's lymphoma of lymph nodes of head, face, and neck (diagnosis)
C0153768|Hodgkin's disease, mixed cellularity of lymph nodes of head, face and neck
C0153768|Hodgkin's disease, mixed cellularity of lymph nodes of head, face AND/OR neck (disorder)
C0153768|Hodgkin's disease, mixed cellularity of lymph nodes of head, face AND/OR neck
C0153768|Hodgkin's disease, mixed cellularity of lymph nodes of head, face and neck (disorder)
C0153768|Hodgkin's disease, mixed cellularity, involving lymph nodes of head, face and neck
C1263911|Primary malignant neoplasm of peripheral nerves of head
C1263911|Primary malignant neoplasm of peripheral nerves of head (diagnosis)
C1263911|neoplasm - pns malignant head primary
C1263911|Primary malignant neoplasm of peripheral nerves of head (disorder)
C0346322|MALIGNANT OPTIC NERVE SHEATH NEOPL
C0346322|OPTIC NERVE SHEATH NEOPL MALIGNANT
C0346322|malignant neoplasm of optic nerve (II) and sheath
C0346322|malignant neoplasm of optic nerve (II) and sheath (diagnosis)
C0346322|malignant neoplasm of optic nerve sheath (diagnosis)
C0346322|neoplasm - malignant of optic nerve (ii) and sheath
C0346322|malignant neoplasm of optic nerve sheath
C0346322|Malignant Optic Nerve Sheath Tumors
C0346322|Optic Nerve Sheath Neoplasms, Malignant
C0346322|Optic Nerve Sheath Tumors, Malignant
C0346322|Malignant Optic Nerve Sheath Neoplasms
C0346322|Malignant tumor of optic nerve and sheath
C0346322|Malignant tumor of optic nerve sheath
C0346322|Malignant tumour of optic nerve and sheath
C0346322|Malignant tumour of optic nerve sheath
C0346322|Malignant tumor of optic nerve and sheath (disorder)
C0346322|Malignant tumor of optic nerve sheath (disorder)
C0684520|bone neoplasm, malignant - skull secondary
C0684520|secondary malignant neoplasm of skull
C0684520|secondary malignant neoplasm of skull (diagnosis)
C0684520|Metastatic malignant neoplasm to bone of skull
C0684520|Secondary malignant neoplasm of bone of skull (disorder)
C0684520|Secondary malignant neoplasm of bone of skull
C0684520|Metastatic malignant neoplasm to bone of skull, NOS
C0684520|Secondary malignant neoplasm of bone of skull, NOS
C0206115|WAGR Syndrome
C0206115|Syndrome, WAGR
C0206115|WAGR Syndromes
C0206115|WAGR
C0206115|WILMS TUMOR, ANIRIDIA, GENITOURINARY ANOMALIES, AND MENTAL RETARDATION SYNDROME
C0206115|Complex, WAGR
C0206115|Contiguous Gene Syndrome, WAGR
C0206115|WAGR Complex
C0206115|Wilms Tumor-Aniridia-Genitourinary Anomalies-MR Syndrome
C0206115|WAGR Contiguous Gene Syndrome
C0206115|WAGR Syndrome [Disease/Finding]
C0206115|Wilms Tumor, Aniridia, Genitourinary Anomalies, Mental Retardation Syndrome
C0206115|Wilms Tumor-Aniridia-Gonadoblastoma-Mental Retardation Syndrome
C0206115|WAGR Complices
C0206115|Chromosome 11p13 Deletion Syndrome
C0206115|11p partial monosomy syndrome
C0206115|anomaly of chromosome pair 11p partial monosomy syndrome
C0206115|11p partial monosomy syndrome (diagnosis)
C0206115|Wilms Tumor-Aniridia-Genital Anomalies-Retardation Syndrome
C0206115|Wilms tumor-aniridia-genitourinary anomalies-mental retardation syndrome
C0206115|Aniridia-Wilms tumor association
C0206115|Aniridia-Wilms tumour association
C0206115|11p partial monosomy syndrome (disorder)
C0496763|Malignant neoplasm of major salivary glands
C0496763|Major salivary gland, unspecified
C0496763|Malignant neoplasm of major salivary gland
C0496763|Malignant neoplasm of major salivary gland, unspecified
C0496763|Malignant neoplasm of salivary gland (major) NOS
C0496763|Malignant neoplasm of major salivary gland NOS
C0496763|Malignant neoplasm of major salivary gland NOS (disorder)
C0496763|malignant salivary gland neoplasm major
C0496763|malignant neoplasm of major salivary gland (diagnosis)
C0496763|Malignant tumor of major salivary gland
C0496763|Malignant tumour of major salivary gland
C0496763|Malignant tumor of major salivary gland (disorder)
C0496763|Malignant neoplasm of major salivary gland, NOS
C0496763|Malignant Major Salivary Gland Neoplasm
C0496763|Malignant Major Salivary Gland Tumor
C0496763|Malignant Neoplasm of the Major Salivary Gland
C0496763|Malignant Tumor of the Major Salivary Gland
C0684967|secondary malignant neoplasm of postcricoid region (diagnosis)
C0684967|hypopharyngeal neoplasm malignant postcricoid region secondary
C0684967|secondary malignant neoplasm of postcricoid region
C0684967|Metastatic malignant neoplasm to postcricoid region
C0684967|Secondary malignant neoplasm of postcricoid region (disorder)
C1305982|cranial nerve neoplasm malignant primary
C1305982|Primary malignant neoplasm of cranial nerve (diagnosis)
C1305982|Primary malignant neoplasm of cranial nerve
C1305982|Primary malignant neoplasm of cranial nerve (disorder)
C1304838|Primary malignant neoplasm of upper respiratory tract
C1304838|malignant neoplasm upper respiratory tract primary
C1304838|Primary malignant neoplasm of upper respiratory tract (diagnosis)
C1304838|Primary malignant neoplasm of upper respiratory tract (disorder)
C0346776|malignant melanoma of the chin (diagnosis)
C0346776|malignant melanoma of the chin
C0346776|Malignant melanoma of chin
C0346776|Malignant melanoma of skin of chin
C0346776|Malignant melanoma of chin (disorder)
C0346776|Malignant melanoma of skin of chin (disorder)
C0347013|Metastasis to nervous system and eye (diagnosis)
C0347013|malignant neoplasm metastatic cancer to nervous system and eye
C0347013|Metastasis to nervous system and eye
C0347013|Metastasis to nervous system and eye (disorder)
C0153810|Sézary's disease of lymph nodes of head, face and neck
C0153810|Sézary's disease of lymph nodes of head, face and neck (disorder)
C0153810|Sézary's disease of lymph nodes of head, face, and neck
C0153810|Sezary syndrome of head, face, and neck (diagnosis)
C0153810|Sezary syndrome of head, face, and neck
C0153810|Sezary's disease of lymph nodes of head, face AND/OR neck
C0153810|Sezary's disease head
C0153810|Sézary disease of lymph nodes of head, face and neck
C0153810|Sézary disease of lymph nodes of head, face AND/OR neck
C0153810|Sézary disease, lymph nodes of head, face, and neck
C0153810|Sezary's disease, lymph nodes of head, face, and neck
C0153810|Sezary's disease involving lymph nodes of head, face, and neck
C0153810|Sézary's disease of lymph nodes of head, face AND/OR neck (disorder)
C0153810|Sezary's disease involving lymph nodes of head, face and neck
C0685010|Secondary malignant neoplasm of laryngeal aspect of aryepiglottic fold
C0685010|Secondary malignant neoplasm of laryngeal aspect of aryepiglottic fold (diagnosis)
C0685010|malignant neoplasm supraglottis laryngeal aspect of aryepiglottic fold secondary
C0685010|Metastatic malignant neoplasm to laryngeal aspect of aryepiglottic fold
C0685010|Secondary malignant neoplasm of laryngeal aspect of aryepiglottic fold (disorder)
C3647449|Malignant neoplasm of anterior wall of nasopharynx
C3647449|Primary malignant neoplasm of anterior wall of nasopharynx (disorder)
C3647449|primary malignant nasopharyngeal neoplasm of anterior wall
C3647449|primary malignant nasopharyngeal neoplasm of anterior wall (diagnosis)
C3647449|nasopharyngeal neoplasm anterior wall, malignant primary
C3647449|Primary malignant neoplasm of anterior wall of nasopharynx
C0686627|Secondary and unspecified malignant neoplasm of occipital lymph nodes (disorder)
C0686627|Secondary and unspecified malignant neoplasm of occipital lymph nodes
C0686627|Secondary malignant neoplasm of occipital lymph nodes
C0686627|Secondary malignant neoplasm of occipital lymph nodes (diagnosis)
C0686627|lymph node neoplasm malignant secondary head occipital
C0686627|Metastatic malignant neoplasm to occipital lymph nodes
C0686627|Secondary malignant neoplasm of occipital lymph nodes (disorder)
C0018197|Granuloma, Lethal Midline
C0018197|Granulomas, Lethal Midline
C0018197|Lethal Midline Granulomas
C0018197|Midline Granuloma, Lethal
C0018197|Midline Granulomas, Lethal
C0018197|Lethal midline granuloma
C0018197|lethal midline granuloma (diagnosis)
C0018197|Midline Lethal Granuloma of Nasal Cavity and Paranasal Sinus
C0018197|Midline Lethal Granuloma of the Nasal Cavity and Paranasal Sinus
C0018197|Nasal Cavity and Paranasal Sinus Lethal Midline Granuloma
C0018197|Granuloma, Lethal Midline [Disease/Finding]
C0018197|Idiopathic midline granuloma
C0018197|Lethal midline granuloma of face
C0018197|Malignant granuloma of face
C0018197|Lethal midline granuloma (disorder)
C0018197|paranasal sinus and nasal cavity midline lethal granuloma
C0018197|lethal midline reticulosis
C0018197|midline lethal granuloma, paranasal sinus and nasal cavity
C0018197|nasal cavity and paranasal sinus midline lethal granuloma
C0018197|granuloma; midline
C0018197|midline; granuloma
C0018197|Midfacial Necrotising Lesion
C0153381|Malignant neoplasm of mouth
C0153381|Malignant neoplasm of mouth, unspecified
C0153381|Mouth, unspecified
C0153381|malignant neoplasm of oral cavity (diagnosis)
C0153381|malignant neoplasm of oral cavity
C0153381|Malignant oral cavity neoplasms
C0153381|Cancers, Mouth
C0153381|Mouth Cancers
C0153381|Cancer, Oral
C0153381|Cancers, Oral
C0153381|Oral Cancers
C0153381|malignant tumor of oral cavity
C0153381|Malig neoplasm mouth NOS
C0153381|Malignant neoplasm of oral cavity NOS
C0153381|Cancer, Mouth
C0153381|Mouth Cancer
C0153381|Malignant tumour of mouth
C0153381|Cancer of oral cavity
C0153381|CA - Mouth cancer
C0153381|Malignant neoplasm of mouth NOS (disorder)
C0153381|Malignant tumor of mouth
C0153381|Malignant neoplasm of mouth NOS
C0153381|Malignant tumour of oral cavity
C0153381|Mouth--Cancer
C0153381|Oral neoplasm malignant
C0153381|Oral Cancer
C0153381|Cancer of the Mouth
C0153381|Malignant tumor of oral cavity (disorder)
C0153381|Malignant neoplasm of mouth, NOS
C0153381|Malignant Mouth Neoplasm
C0153381|Malignant Mouth Tumor
C0153381|Malignant Neoplasm of the Mouth
C0153381|Malignant Oral Cavity Neoplasm
C0153381|Malignant Oral Cavity Tumor
C0153381|Malignant Oral Neoplasm
C0153381|Malignant Tumor of the Mouth
C0153381|Cancer of Mouth
C0684992|Secondary malignant neoplasm of vocal cord
C0684992|Secondary malignant neoplasm of vocal cord (diagnosis)
C0684992|laryngeal neoplasm vocal cord malignant secondary
C0684992|Metastatic malignant neoplasm to vocal cord
C0684992|Secondary malignant neoplasm of vocal cord (disorder)
C0684748|Secondary malignant neoplasm of muscle of head
C0684748|Secondary malignant neoplasm of muscle of head (diagnosis)
C0684748|malignant neoplasm of muscle of head secondary
C0684748|Metastatic malignant neoplasm to muscle of head
C0684748|Secondary malignant neoplasm of muscle of head (disorder)
C0240803|Primary Cerebral Lymphoma
C0240803|Primary Lymphoma of Cerebrum
C0240803|Primary Lymphoma of the Cerebrum
C0240803|Primary Lymphoma, Brain
C0240803|malignant lymphoma of brain (diagnosis)
C0240803|malignant lymphoma of brain
C0240803|neoplasm - brain cerebrum, malignant primary lymphoma
C0240803|Primary cerebral lymphoma (diagnosis)
C0240803|primary malignant lymphoma of brain (diagnosis)
C0240803|primary malignant lymphoma of brain
C0240803|malignant neoplasm lymphoma of brain primary
C0240803|Brain lymphoma
C0240803|Cerebral lymphoma
C0240803|Primary cerebral lymphoma (disorder)
C0686612|Secondary malignant neoplasm of adenoid (diagnosis)
C0686612|Secondary malignant neoplasm of adenoid
C0686612|Metastatic malignant neoplasm to adenoid
C0686612|Secondary malignant neoplasm of adenoid (disorder)
C0686507|Metastatic Neoplasm to the Parathyroid
C0686507|Metastatic Parathyroid Neoplasm
C0686507|Metastatic Malignant Parathyroid Gland Neoplasm
C0686507|Secondary malignant neoplasm of parathyroid gland (diagnosis)
C0686507|Secondary malignant neoplasm of parathyroid gland
C0686507|parathyroid neoplasm malignant secondary
C0686507|Metastatic Malignant Neoplasm in the Parathyroid Glands
C0686507|Metastatic Malignant Neoplasm to the Parathyroid Glands
C0686507|Metastatic malignant neoplasm to parathyroid gland
C0686507|Secondary malignant neoplasm of parathyroid gland (disorder)
C0686507|Metastasis to the Parathyroid Gland
C0686507|Metastatic Neoplasm of Parathyroid Gland
C0686507|Metastatic Neoplasm of Parathyroid
C0686507|Metastatic Neoplasm of the Parathyroid Gland
C0686507|Metastatic Neoplasm of the Parathyroid
C0686507|Metastatic Neoplasm to the Parathyroid Gland
C0686507|Metastatic Parathyroid Gland Neoplasm
C0686507|Metastatic Parathyroid Gland Tumor
C0686507|Metastatic Parathyroid Tumor
C0686507|Metastatic Tumor of Parathyroid Gland
C0686507|Metastatic Tumor of Parathyroid
C0686507|Metastatic Tumor of the Parathyroid Gland
C0686507|Metastatic Tumor of the Parathyroid
C0686507|Metastatic Tumor to the Parathyroid Gland
C0686507|Metastatic Tumor to the Parathyroid
C0153776|Hodgkin's disease, lymphocytic depletion of lymph nodes of head, face, and neck
C0153776|lymphocyte depletion Hodgkin's disease of lymph nodes of head, face, or neck
C0153776|lymphocyte depletion Hodgkin's disease of lymph nodes of head, face, or neck (diagnosis)
C0153776|Hodgkin's disease, lymphocytic depletion, involving lymph nodes of head, face, and neck.
C0153776|Hodg lymph deplet head
C0153776|Hodgkin disease, lymphocytic depletion of lymph nodes of head, face AND/OR neck
C0153776|Hodgkin disease, lymphocytic depletion of lymph nodes of head, face and neck
C0153776|Hodgkin's disease, lymphocytic depletion, lymph nodes of head, face, and neck
C0153776|Hodgkin's disease, lymphocytic depletion, involving lymph nodes of head, face, and neck
C0153776|Hodgkin's disease, lymphocytic depletion of lymph nodes of head, face and neck
C0153776|Hodgkin's disease, lymphocytic depletion of lymph nodes of head, face AND/OR neck (disorder)
C0153776|Hodgkin's disease, lymphocytic depletion of lymph nodes of head, face AND/OR neck
C0153776|Hodgkin's disease, lymphocytic depletion of lymph nodes of head, face and neck (disorder)
C0153776|Hodgkin's disease, lymphocytic depletion, involving lymph nodes of head, face and neck
C0685991|Metastatic malignant neoplasm to submaxillary gland
C0685991|Secondary malignant neoplasm of submaxillary gland
C0685991|Secondary malignant neoplasm of submaxillary gland (disorder)
C1304847|jaw neoplasm malignant primary
C1304847|Primary malignant neoplasm of jaw (diagnosis)
C1304847|Primary malignant neoplasm of jaw
C1304847|Primary malignant neoplasm of jaw (disorder)
C0153350|Malignant neoplasm of base of tongue
C0153350|malignant neoplasm of base of tongue (diagnosis)
C0153350|malignant tumor of base of tongue
C0153350|Mal neo tongue base
C0153350|Malignant neoplasm of posterior third of tongue
C0153350|Malignant neoplasm of fixed part of tongue NOS
C0153350|Malignant neoplasm of fixed part of tongue NOS (disorder)
C0153350|Malignant tumor of fixed part of tongue
C0153350|Malignant tumor of posterior third of tongue
C0153350|Malignant tumor of tongue posterior to vallate papillae
C0153350|Malignant tumour of base of tongue
C0153350|Malignant tumour of fixed part of tongue
C0153350|Malignant tumour of posterior third of tongue
C0153350|Malignant tumour of tongue posterior to vallate papillae
C0153350|Malignant tumor of base of tongue (disorder)
C0153350|Malignant Base of Tongue Neoplasm
C0153350|Malignant Base of Tongue Tumor
C0153350|Malignant Base of the Tongue Neoplasm
C0153350|Malignant Base of the Tongue Tumor
C0153350|Malignant Neoplasm of Posterior Tongue
C0153350|Malignant Neoplasm of the Base of the Tongue
C0153350|Malignant Neoplasm of the Posterior Tongue
C0153350|Malignant Posterior Tongue Neoplasm
C0153350|Malignant Posterior Tongue Tumor
C0153350|Malignant Tumor of Posterior Tongue
C0153350|Malignant Tumor of the Base of the Tongue
C0153350|Malignant Tumor of the Posterior Tongue
C0345741|Malignant neoplasm of false vocal cord
C0345741|Malignant neoplasm of ventricular bands of larynx
C0345741|laryngeal neoplasm false vocal cord malignant
C0345741|malignant neoplasm of false vocal cord (diagnosis)
C0345741|Malignant tumor of false cord
C0345741|Malignant tumor of ventricular band
C0345741|Malignant tumor of vestibular fold
C0345741|Malignant tumour of false cord
C0345741|Malignant tumour of ventricular band
C0345741|Malignant tumour of vestibular fold
C0345741|Malignant tumor of false cord (disorder)
C0345741|Malignant neoplasm of false vocal cords
C0686013|Secondary malignant neoplasm of floor of mouth
C0686013|floor of mouth malignant neoplasm secondary
C0686013|Secondary malignant neoplasm of floor of mouth (diagnosis)
C0686013|Secondary malignant neoplasm of floor of mouth (disorder)
C0686013|Metastatic malignant neoplasm to floor of mouth
C0686013|Metastatic malignant neoplasm to floor of mouth, NOS
C0686013|Secondary malignant neoplasm of floor of mouth, NOS
C0345756|pharyngeal neoplasm malignant parapharynegal space
C0345756|malignant neoplasm of parapharyngeal space
C0345756|malignant neoplasm of parapharyngeal space (diagnosis)
C0345756|Malignant tumor of parapharyngeal space
C0345756|Malignant tumour of parapharyngeal space
C0345756|Malignant tumor of parapharyngeal space (disorder)
C0685129|Malignant neoplasm of blood vessel of head
C0685129|Primary malignant neoplasm of blood vessel of head (diagnosis)
C0685129|Primary malignant neoplasm of blood vessel of head
C0685129|neoplasm - soft tissue types blood vessel malignant of head primary
C0685129|Primary malignant neoplasm of blood vessel of head (disorder)
C0153405|Malignant neoplasm of pharynx
C0153405|Malignant neoplasm of pharynx, unspecified
C0153405|Pharynx, unspecified
C0153405|malignant neoplasm of pharynx (diagnosis)
C0153405|malignant pharyngeal neoplasm
C0153405|Cancer, Pharnyx
C0153405|Cancers, Pharnyx
C0153405|Pharnyx Cancers
C0153405|Cancer, Pharyngeal
C0153405|Cancers, Pharyngeal
C0153405|Pharyngeal Cancers
C0153405|Pharynx Cancer
C0153405|Pharynx Cancers
C0153405|Pharyngeal cancer
C0153405|malignant tumor of pharynx
C0153405|Mal neo pharynx NOS
C0153405|Malignant neoplasm of pharynx unspecified (disorder)
C0153405|Malignant neoplasm of pharynx unspecified
C0153405|Pharynx--Cancer
C0153405|Pharyngeal cancer stage unspecified
C0153405|Pharynx neoplasm malignant
C0153405|Cancer of the Pharynx
C0153405|Pharnyx Cancer
C0153405|Malignant tumour of pharynx
C0153405|CA - Cancer of pharynx
C0153405|Cancer of pharynx
C0153405|Malignant tumor of pharynx (disorder)
C0153405|Malignant neoplasm of pharynx, NOS
C0153405|Malignant Pharyngeal Tumor
C0153405|Malignant Pharynx Neoplasm
C0153405|Malignant Pharynx Tumor
C0153405|Malignant Tumor of the Pharynx
C0346825|Malignant tumor of soft tissue of head, face and neck
C0346825|Malignant tumour of soft tissue of head, face and neck
C0346825|Malignant tumor of soft tissue of head, face and neck (disorder)
C0153760|Hodgkin's disease, nodular sclerosis of lymph nodes of head, face, and neck
C0153760|Hodgkin's disease, nodular sclerosis, involving lymph nodes of head, face, and neck.
C0153760|Hodg nodul sclero head
C0153760|Hodgkin disease, nodular sclerosis of lymph nodes of head, face and neck
C0153760|Hodgkin disease, nodular sclerosis of lymph nodes of head, face AND/OR neck
C0153760|Hodgkin's disease, nodular sclerosis, lymph nodes of head, face, and neck
C0153760|Hodgkin's disease, nodular sclerosis, involving lymph nodes of head, face, and neck
C0153760|nodular sclerosing Hodgkin's disease of lymph nodes of head, face, and neck
C0153760|nodular sclerosis Hodgkin's lymphoma of lymph nodes of head, face, and neck
C0153760|nodular sclerosing Hodgkin's disease of lymph nodes of head, face, and neck (diagnosis)
C0153760|Hodgkin's disease, nodular sclerosis of lymph nodes of head, face and neck
C0153760|Hodgkin's disease, nodular sclerosis of lymph nodes of head, face AND/OR neck (disorder)
C0153760|Hodgkin's disease, nodular sclerosis of lymph nodes of head, face AND/OR neck
C0153760|Hodgkin's disease, nodular sclerosis of lymph nodes of head, face and neck (disorder)
C0153760|Hodgkin's disease, nodular sclerosis, involving lymph nodes of head, face and neck
C0153794|Nodular lymphoma head
C0153794|Nodular lymphoma, lymph nodes of head, face, and neck
C0153794|Nodular lymphoma involving lymph nodes of head, face, and neck
C0153794|Nodular lymphoma of lymph nodes of head, face, and neck (disorder)
C0153794|Nodular lymphoma of lymph nodes of head, face, and neck
C0153794|nodular lymphoma of lymph nodes of head, face, and neck (diagnosis)
C0153794|Nodular lymphoma of lymph nodes of head, face and neck
C0153794|Nodular lymphoma of lymph nodes of head, face and neck (disorder)
C0153794|Nodular lymphoma involving lymph nodes of head, face and neck
C1290119|Melanoma in situ of face (disorder)
C1290119|Melanoma in situ of face
C1290119|face; melanoma in situ
C1290119|melanoma in situ; face
C0751255|Malignant neoplasm of jaw
C0751255|malignant neoplasm of jaw (diagnosis)
C0751255|Cancers, Jaw
C0751255|Jaw Cancers
C0751255|malignant tumor of jaw
C0751255|Cancer, Jaw
C0751255|Malignant neoplasm of jaw NOS
C0751255|Malignant neoplasm of jaw NOS (disorder)
C0751255|Jaws--Cancer
C0751255|Jaw Cancer
C0751255|Cancer of the Jaw
C0751255|Malignant neoplasm of jaw, NOS
C0751255|Cancer of Jaw
C0346944|Malignant neoplasm of supraclavicular fossa NOS
C0346944|Malignant neoplasm of supraclavicular fossa NOS (disorder)
C1299284|Primary malignant neoplasm of false vocal cord
C1299284|Primary malignant neoplasm of false vocal cord (disorder)
C1299284|laryngeal neoplasm false vocal cord malignant primary
C1299284|Primary malignant neoplasm of false vocal cord (diagnosis)
C0751177|Malignant neoplasm of head
C0751177|head cancer
C0751177|Malignant neoplasm of head NOS
C0751177|Malignant neoplasm of head NOS (disorder)
C0751177|malignant neoplasm of ill-defined site head
C0751177|malignant neoplasm of head (diagnosis)
C0751177|Head--Cancer
C0751177|Cancer of Head
C0751177|Cancer of the Head
C0751177|Malignant neoplasm of head, NOS
C0349019|Malignant neoplasm of peripheral nerves of head, face and neck
C0349019|Peripheral nerves of head, face and neck
C0349019|Malignant neoplasm of prph nerves of head, face and neck
C0349019|malignant neoplasm of peripheral nerves of head, face, and neck (diagnosis)
C0349019|malignant neoplasm of peripheral nerves of head, face, and neck
C0349019|neoplasm - pns peripheral malignant head face and neck
C0349019|Malignant neoplasm of peripheral nerves of head, face and neck (disorder)
C0587060|Malignant melanoma of head and neck
C0587060|Malignant melanoma of head and neck (disorder)
C0587060|malignant melanoma of head and neck (diagnosis)
C0587060|malignant neoplasm of ill-defined site head and neck melanoma
C0346568|malignant neoplasm of ear, nose, and throat (diagnosis)
C0346568|malignant neoplasm of ill-defined site ear, nose, and throat
C0346568|malignant neoplasm of ear, nose, and throat
C0346568|Malignant tumor of ear, nose and throat
C0346568|Malignant tumour of ear, nose and throat
C0346568|Malignant tumor of ear, nose and throat (disorder)
C0496836|Eye, unspecified
C0496836|Malignant neoplasm of eye, unspecified
C0496836|Malignant tumor of eye
C0496836|malignant neoplasm of eye
C0496836|malignant neoplasm of eye (diagnosis)
C0496836|eye cancer (diagnosis)
C0496836|eye cancer
C0496836|malignant eye neoplasm
C0496836|Cancers, Eye
C0496836|Eye Cancers
C0496836|Malign neopl eye NOS
C0496836|Malignant neoplasm of unspecified site of eye
C0496836|Cancer, Eye
C0496836|Malignant tumour of eye
C0496836|Malignant neoplasm of eye NOS
C0496836|Ca eye
C0496836|Malignant neoplasm of eye NOS (disorder)
C0496836|Eye--Cancer
C0496836|Malignant eye cancer, NOS
C0496836|Malignant neoplasm of eye, part unspecified
C0496836|Malignant eye neoplasm NOS
C0496836|Cancer of the Eye
C0496836|Malignant tumor of eye (disorder)
C0496836|ocular cancer
C0496836|Malignant neoplasm of eye, NOS
C0496836|Cancer of Eye
C0496836|Eye Neoplasm, Malignant
C0496836|Malignant Eye Tumor
C0496836|Malignant Neoplasm of the Eye
C0496836|Malignant Ocular Neoplasm
C0496836|Malignant Ocular Tumor
C0496836|Malignant Tumor of the Eye
C0496836|Neoplasm malig;eye
C0496836|malignant neosplasm of the eye
C0153645|Malignant neoplasm of cerebral meninges
C0153645|Cerebral meninges
C0153645|malignant neoplasm of cerebral meninges (diagnosis)
C0153645|malignant tumor of cerebral meninges
C0153645|Mal neo cerebral mening
C0153645|Malignant neoplasm of cerebral meninges NOS (disorder)
C0153645|Malignant neoplasm of cerebral meninges NOS
C0153645|Cancer of the cerebral meninges
C0153645|Malignant neoplasm of cerebral meninges (disorder)
C0346653|Malignant neoplasm of bones of skull and face
C0346653|Bones of skull and face
C0346653|Malignant neoplasm of bones of skull and face NOS (disorder)
C0346653|Malignant neoplasm of bones of skull and face NOS
C0346653|bone neoplasm, malignant - skull and face
C0346653|malignant neoplasm of bones of skull and face (diagnosis)
C0346653|Malignant neoplasm of bones of skull and face (disorder)
C0178247|Malignant neoplasm of lip, oral cavity and pharynx (disorder)
C0178247|Malignant neoplasm of lip, oral cavity and/or pharynx (disorder)
C0178247|Malignant neoplasms of lip, oral cavity and pharynx
C0178247|Malignant neoplasms of lip, oral cavity and pharynx (C00-C14)
C0178247|Malignant neoplasm of lip, oral cavity and pharynx
C0178247|Malignant neoplasm of lip, oral cavity and pharynx NOS
C0178247|Ca lip, oral, pharynx NOS
C0178247|Malignant neoplasm: [lip] or [oral cavity] or [pharynx] (disorder)
C0178247|Ca lip, oral, pharynx
C0178247|Malignant neoplasm: [lip] or [oral cavity] or [pharynx]
C0178247|Ca lip, oral, pharynx NOS (disorder)
C0178247|Malignant neoplasm of lip, oral cavity and pharynx NOS (disorder)
C0178247|malignant neoplasm of lip, oral cavity, and/or pharynx (diagnosis)
C0178247|malignant neoplasm of lip, oral cavity, and/or pharynx
C0178247|MALIGNANT NEOPLASM OF LIP, ORAL CAVITY, AND PHARYNX
C1828015|Malignant tumor of eyelid (disorder)
C1828015|Malignant neoplasm of eyelid (disorder)
C1828015|Malignant neoplasm of skin of eyelid (disorder)
C1828015|Malignant neoplasm of skin of eyelid
C1828015|Malignant neoplasm of eyelid
C1828015|skin neoplasm eyelid malignant
C1828015|malignant neoplasm of skin of eyelid (diagnosis)
C1828015|malignant neoplasm of eyelid (diagnosis)
C1828015|neoplasm of ocular adnexa eyelid malignant
C1828015|Malignant tumor of eyelid
C1828015|Malignant tumour of eyelid
C1828015|Malignant Eyelid Neoplasm
C1828015|Malignant Eyelid Tumor
C1828015|Malignant Neoplasm of the Eyelid
C1828015|Malignant Tumor of the Eyelid
C0684808|Malignant neoplasm of face
C0684808|malignant neoplasm of face (diagnosis)
C0684808|Malignant tumor of face
C0684808|Malignant tumour of face
C0684808|Malignant tumor of face (disorder)
C0684808|Malignant neoplasm of face, NOS
C0153627|Malignant neoplasm of lacrimal gland
C0153627|malignant neoplasm of lacrimal gland (diagnosis)
C0153627|lacrimal gland neoplasm malignant
C0153627|Mal neo lacrimal gland
C0153627|Malignant tumour of lacrimal gland
C0153627|Malignant tumour of lacrimal gland (disorder)
C0153627|Malignant tumor of lacrimal gland
C0153627|Malignant tumor of lacrimal gland (disorder)
C0153627|Malignant Lacrimal Gland Neoplasm
C0153627|Malignant Lacrimal Gland Tumor
C0153627|Malignant Neoplasm of the Lacrimal Gland
C0153627|Malignant Tumor of the Lacrimal Gland
C0153626|Orbit
C0153626|Malignant neoplasm of orbit
C0153626|Malignant tumor of orbit
C0153626|malignant neoplasm of orbit (diagnosis)
C0153626|Malign neopl orbit
C0153626|Malignant neoplasm of orbit NOS
C0153626|Malignant neoplasm of orbit NOS (disorder)
C0153626|Malignant orbital tumor
C0153626|Malignant orbital tumour
C0153626|Malignant tumour of orbit
C0153626|Malignant tumor of orbit (disorder)
C0153626|Malignant Neoplasm of the Orbit
C0153626|Malignant Orbit Neoplasm
C0153626|Malignant Orbit Tumor
C0153626|Malignant Orbital Neoplasm
C0153626|Malignant Tumor of the Orbit
C0686574|Malignant mast cell tumors involving lymph nodes of head, face, and neck
C0686574|Malignant mast cell tumor of lymph nodes of head, face, and neck
C0686574|malignant mastocytosis of head, face, and neck (diagnosis)
C0686574|malignant mastocytosis of head, face, and neck
C0686574|Mal mastocytosis head
C0686574|Malignant mast cell tumors, lymph nodes of head, face, and neck
C0686574|mast cell malignancy of lymph nodes of head, face, and neck
C0686574|Mast cell malignancy of lymph nodes of head, face and neck
C0686574|mast cell malignancy of lymph nodes of head, face, and neck (diagnosis)
C0686574|Malignant mast cell tumor of lymph nodes of head, face AND/OR neck (disorder)
C0686574|Malignant mast cell tumor of lymph nodes of head, face AND/OR neck
C0686574|Malignant mast cell tumour of lymph nodes of head, face AND/OR neck
C0686574|Mast cell malignancy of lymph nodes of head, face and neck (disorder)
C0686574|Malignant mast cell tumors involving lymph nodes of head, face and neck
C0346903|Malignant neoplasm of cerebrum
C0346903|Malignant neoplasm of cerebrum (disorder)
C0346903|malignant neoplasm of cerebral hemisphere (diagnosis)
C0346903|malignant neoplasm of cerebral hemisphere
C0346903|malignant tumor of cerebral hemisphere
C0346903|Cerebral tumor (malignant)
C0346903|Cerebral tumor - malignant (disorder)
C0346903|Cerebrum Ca (disorder)
C0346903|Malignant cerebral tumor
C0346903|Malignant neoplasm of cerebrum NOS
C0346903|Cerebrum Ca
C0346903|Cerebral tumour (malignant)
C0346903|Cerebral tumour - malignant
C0346903|Malignant neoplasm of cerebrum NOS (disorder)
C0346903|Cerebral tumor - malignant
C0346903|Malignant cerebral tumour
C0346903|malignant neoplasm of cerebrum (diagnosis)
C0346903|brain tumor malignant of cerebrum
C0346903|Malignant neoplasm of cerebrum, NOS
C0346903|Malignant Cerebral Hemispheric Neoplasm
C0346903|Malignant Cerebral Hemispheric Tumor
C0346903|Malignant Cerebral Neoplasm
C0346903|Malignant Neoplasm of Cerebral Hemispheres
C0346903|Malignant Neoplasm of the Cerebral Hemispheres
C0346903|Malignant Neoplasm of the Cerebrum
C0346903|Malignant Tumor of Cerebral Hemispheres
C0346903|Malignant Tumor of Cerebrum
C0346903|Malignant Tumor of the Cerebral Hemispheres
C0346903|Malignant Tumor of the Cerebrum
C0346903|Cerebral Cancer
C0580284|Metastasis to head and neck lymph node
C0580284|Metastasis to head and neck lymph node (disorder)
C0580284|Metastasis to head and neck lymph node (diagnosis)
C0580284|metastatic cancer to head and neck lymph node
C1306467|Primary malignant neoplasm of head (diagnosis)
C1306467|malignant neoplasm of ill-defined site head primary
C1306467|Primary malignant neoplasm of head
C1306467|Primary malignant neoplasm of head (disorder)
C0349750|eye neoplasm malignant lacrimal drainage structure
C0349750|malignant neoplasm of lacrimal drainage structure (diagnosis)
C0349750|malignant neoplasm of lacrimal drainage structure
C0349750|Malignant tumor of lacrimal drainage structure
C0349750|Malignant tumour of lacrimal drainage structure
C0349750|Malignant tumor of lacrimal drainage structure (disorder)
C0684805|Secondary malignant neoplasm of head
C0684805|Secondary malignant neoplasm of head (diagnosis)
C0684805|malignant neoplasm of ill-defined site head secondary
C0684805|Metastatic malignant neoplasm to head
C0684805|Secondary malignant neoplasm of head (disorder)
C0684805|Metastatic malignant neoplasm to head, NOS
C0684805|Secondary malignant neoplasm of head, NOS
C0432547|Letterer-Siwe disease of lymph nodes of head, face, and neck
C0432547|Letterer-Siwe disease of head, face, or neck
C0432547|Letterer-Siwe disease of head, face, or neck (diagnosis)
C0432547|Letterer-siwe dis head
C0432547|Letterer-siwe disease, lymph nodes of head, face, and neck
C0432547|Letterer-Siwe disease involving lymph nodes of head, face, and neck
C0432547|Letterer-Siwe disease of lymph nodes of head, face and neck
C0432547|Letterer-Siwe disease of lymph nodes of head, face and neck (disorder)
C0432547|Letterer-Siwe disease of lymph nodes of head, face AND/OR neck (disorder)
C0432547|Letterer-Siwe disease of lymph nodes of head, face AND/OR neck
C0432547|Letterer-Siwe disease involving lymph nodes of head, face and neck
C0432538|Malignant histiocytosis of lymph nodes of head, face, and neck
C0432538|Mal histiocytosis head
C0432538|Malignant histiocytosis, lymph nodes of head, face, and neck
C0432538|Malignant histiocytosis involving lymph nodes of head, face, and neck
C0432538|malignant histiocytosis of lymph nodes of head, face, and neck (diagnosis)
C0432538|reticuloendothelial system malignant histiocytosis lymph node head, face, neck
C0432538|Malignant histiocytosis of lymph nodes of head, face and neck
C0432538|Malignant histiocytosis of lymph nodes of head, face AND/OR neck (disorder)
C0432538|Malignant histiocytosis of lymph nodes of head, face AND/OR neck
C0432538|Malignant histiocytosis of lymph nodes of head, face and neck (disorder)
C0432538|Malignant histiocytosis involving lymph nodes of head, face and neck
C0432556|lymphoma of head, face, and neck
C0432556|lymphoma of head, face, and neck (diagnosis)
C0432556|Malignant lymphoma NOS of lymph nodes of head, face and neck (disorder)
C0432556|Malignant lymphoma NOS of lymph nodes of head, face and neck
C0432556|Malignant lymphoma of lymph nodes of head, face AND/OR neck (disorder)
C0432556|Malignant lymphoma of lymph nodes of head, face AND/OR neck
C0432556|Malignant lymphoma, NOS of lymph nodes of head, face, and neck
C1719786|Malignant lymphoma of the eye region (disorder)
C1719786|Malignant lymphoma of the eye region
C1827431|Sarcoma of head and neck (disorder)
C1827431|Sarcoma of head and neck
C1827431|malignant neoplasm sarcoma of head and neck (diagnosis)
C1827431|malignant neoplasm sarcoma of head and neck
C0007107|Malignant neoplasm of larynx
C0007107|laryngeal cancer
C0007107|Malignant neoplasm of larynx, unspecified
C0007107|Larynx, unspecified
C0007107|malignant neoplasm of larynx (diagnosis)
C0007107|malignant laryngeal neoplasm
C0007107|Cancer, Laryngeal
C0007107|Cancers, Laryngeal
C0007107|Laryngeal Cancers
C0007107|Cancers, Larynx
C0007107|Larynx Cancers
C0007107|malignant tumor of larynx
C0007107|cancer of larynx
C0007107|Malignant neo larynx NOS
C0007107|Cancer, Larynx
C0007107|Laryngeal neoplasms malignant
C0007107|laryngeal cancer (diagnosis)
C0007107|Malignant neoplasm of larynx NOS (disorder)
C0007107|Ca larynx - NOS
C0007107|Malignant neoplasm of larynx NOS
C0007107|Ca larynx - NOS (disorder)
C0007107|Malignant tumour of larynx
C0007107|CA - Cancer of larynx
C0007107|Larynx--Cancer
C0007107|Laryngeal cancer NOS
C0007107|Larynx cancer
C0007107|Larynx neoplasm malignant
C0007107|Cancer of the Larynx
C0007107|Malignant tumor of larynx (disorder)
C0007107|Malignant neoplasm of larynx, NOS
C0007107|Malignant Laryngeal Tumor
C0007107|Malignant Larynx Neoplasm
C0007107|Malignant Larynx Tumor
C0007107|Malignant Neoplasm of the Larynx
C0007107|Malignant Tumor of the Larynx
C0007107|Neoplasm malig;larynx
C0007107|malignant neosplasm of the larynx
C0220635|Squamous Cell Carcinoma Metastatic in the Neck with Occult Primary
C0220635|Squamous Cell Carcinoma Metastatic to the Neck with Occult Primary
C0220635|Epidermoid Carcinoma Metastatic to the Neck with Occult Primary
C0220635|metastatic squamous neck cancer with occult primary
C0220635|neck cancer, metastatic squamous with occult primary
C0220635|occult primary cancer metastatic squamous to the neck
C0238301|Cancer, Nasopharyngeal
C0238301|Cancers, Nasopharyngeal
C0238301|Nasopharyngeal Cancers
C0238301|Cancers, Nasopharynx
C0238301|Nasopharynx Cancers
C0238301|Cancer, Nasopharynx
C0238301|Cancer of Nasopharynx
C0238301|Nasopharyngeal cancer
C0238301|Nasopharynx--Cancer
C0238301|Cancer of the Nasopharynx
C0238301|Nasopharynx Cancer
C0238301|CA - Cancer of nasopharynx
C1710095|Sinonasal Carcinoma
C1710095|Nasal Cavity and Paranasal Sinus Carcinoma
C1710095|paranasal sinus and nasal cavity cancer
C1710095|nasal cavity and paranasal sinus cancer
C0153398|Malignant neoplasm of hypopharynx
C0153398|Malignant neoplasm of hypopharynx, unspecified
C0153398|Hypopharynx, unspecified
C0153398|malignant neoplasm of hypopharynx (diagnosis)
C0153398|malignant hypopharyngeal neoplasm
C0153398|Cancer, Hypopharyngeal
C0153398|Cancers, Hypopharyngeal
C0153398|Hypopharyngeal Cancers
C0153398|malignant tumor of hypopharynx
C0153398|Mal neo hypopharynx NOS
C0153398|Malignant neoplasm of hypopharynx, unspecified site
C0153398|Hypopharyngeal Cancer
C0153398|Malignant neoplasm of hypopharynx NOS (disorder)
C0153398|Malignant tumour of hypopharynx
C0153398|Malignant neoplasm of hypopharynx NOS
C0153398|Malignant tumour of hypopharynx (disorder)
C0153398|Hypopharynx--Cancer
C0153398|Malignant neoplasm of laryngopharynx
C0153398|Malignant tumor of laryngopharynx
C0153398|Malignant tumour of laryngopharynx
C0153398|Malignant tumor of hypopharynx (disorder)
C0153398|hypopharynx cancer
C0153398|Malignant neoplasm of hypopharynx, NOS
C0153398|Malignant Hypopharyngeal Tumor
C0153398|Malignant Neoplasm of the Hypopharynx
C0153398|Malignant Tumor of the Hypopharynx
C0687150|Parathyroid Carcinoma
C0687150|Parathyroid Gland Carcinoma
C0687150|Parathyroid carcinomas
C0687150|carcinoma of parathyroid gland (diagnosis)
C0687150|adenocarcinoma of parathyroid gland
C0687150|adenocarcinoma of parathyroid gland (diagnosis)
C0687150|carcinoma of parathyroid gland
C0687150|Cancers, Parathyroid
C0687150|Parathyroid Cancers
C0687150|parathyroid adenocarcinoma
C0687150|Parathyroid Gland Cancer
C0687150|Cancer, Parathyroid
C0687150|parathyroid cancer
C0687150|Parathyroid cancer, NOS
C0687150|PRTC
C0687150|Cancer of Parathyroid
C0687150|Cancer of the Parathyroid
C0687150|Parathyroid carcinoma (disorder)
C0687150|carcinoma of the parathyroid
C0687150|Parathyroid Gland Adenocarcinoma
C0687150|Adenocarcinoma of Parathyroid
C0687150|Adenocarcinoma of the Parathyroid Gland
C0687150|Adenocarcinoma of the Parathyroid
C0687150|Cancer of Parathyroid Gland
C0687150|Cancer of the Parathyroid Gland
C0687150|Carcinoma of Parathyroid
C0687150|Carcinoma of the Parathyroid Gland
C0687150|Carcinoma, Parathyroid
C0687150|Carcinomas, Parathyroid
C2349952|carcinoma of oropharynx (diagnosis)
C2349952|carcinoma of oropharynx
C2349952|Oropharyngeal Carcinoma
C2349952|Oropharnyx Cancer
C2349952|Oropharnyx Cancers
C2349952|Cancer, Oropharyngeal
C2349952|Cancers, Oropharyngeal
C2349952|Oropharyngeal Cancers
C2349952|Cancer, Oropharynx
C2349952|Cancers, Oropharynx
C2349952|Oropharynx Cancers
C2349952|Oropharyngeal cancer
C2349952|Cancer of the Oropharynx
C2349952|Oropharynx Cancer
C2349952|Oropharynx Carcinoma
C2349952|Cancer of Oropharynx
C2349952|Carcinoma of the Oropharynx
C2349952|Cancer of Oropharnyx
C0220641|Oral Cancer
C0220641|Oral Carcinoma
C0220641|Lip and Oral Cavity Carcinoma
C0220641|lip and oral cavity cancer
C0220641|oral cavity and lip cancer
C0496842|Pituitary gland
C0496842|Malignant neoplasm of pituitary gland
C0496842|malignant neoplasm of pituitary gland (diagnosis)
C0496842|malignant pituitary neoplasm
C0496842|malignant tumor of pituitary gland
C0496842|Pituitary cancer
C0496842|Malignant pituitary tumour
C0496842|Pituitary tumor malignant
C0496842|Malignant pituitary tumor
C0496842|Pituitary tumour malignant NOS
C0496842|Pituitary tumour malignant
C0496842|Pituitary tumor malignant NOS
C0496842|Malignant tumour of pituitary gland
C0496842|CA - Cancer of pituitary gland
C0496842|Cancer of pituitary gland
C0496842|Malignant tumor of pituitary gland (disorder)
C0496842|Malignant Neoplasm of Pituitary
C0496842|Malignant Neoplasm of the Pituitary Gland
C0496842|Malignant Neoplasm of the Pituitary
C0496842|Malignant Pituitary Gland Neoplasm
C0496842|Malignant Pituitary Gland Tumor
C0496842|Malignant Tumor of Pituitary
C0496842|Malignant Tumor of the Pituitary Gland
C0496842|Malignant Tumor of the Pituitary
C0496842|Pituitary Neoplasms, Malignant
C0496842|Pituitary Tumor, Malignant
C0153656|Malignant neoplasm of carotid body
C0153656|Carotid body
C0153656|carotid body tumor malignant
C0153656|malignant neoplasm of carotid body (diagnosis)
C0153656|Mal neo carotid body
C0153656|Malignant neoplasm of carotid body (disorder)
C0153656|Cancer of carotid body
C0153656|CHEMODECTOMA, MALIGNANT
C0153656|Malignant Carotid Body Neoplasm
C0153656|Malignant Tumor of Carotid Body
C0153656|Malignant Tumor of the Carotid Body
C0153656|Malignant Carotid Body Tumor
C0153656|Malignant Neoplasm of the Carotid Body
C0153656|Malignant carotid body tumour
C0153656|Malignant carotid body tumor (morphologic abnormality)
C0153656|Malignant Carotid Body Paraganglioma
C0153474|Malignant neoplasm of accessory sinus, unspecified
C0153474|Malignant tumor of nasal sinuses
C0153474|Accessory sinus, unspecified
C0153474|Malignant neoplasm of accessory sinuses
C0153474|Malignant neoplasm of accessory sinus
C0153474|malignant neoplasm of accessory sinus (diagnosis)
C0153474|Nasal sinus cancer
C0153474|malignant tumor of accessory sinus
C0153474|Mal neo access sinus NOS
C0153474|Malignant neoplasm of accessory sinus NOS (disorder)
C0153474|Malignant neoplasm of accessory sinus NOS
C0153474|Malignant tumour of nasal sinuses
C0153474|Malignant tumor of nasal sinuses (disorder)
C0153474|Malignant neoplasm of accessory sinus, NOS
C0153474|Malignant Accessory Sinus Neoplasm
C0153474|Malignant Accessory Sinus Tumor
C0153474|Malignant Neoplasm of Paranasal Sinus
C0153474|Malignant Neoplasm of the Accessory Sinus
C0153474|Malignant Neoplasm of the Paranasal Sinus
C0153474|Malignant Paranasal Sinus Neoplasm
C0153474|Malignant Paranasal Sinus Tumor
C0153474|Malignant Tumor of Paranasal Sinus
C0153474|Malignant Tumor of the Accessory Sinus
C0153474|Malignant Tumor of the Paranasal Sinus
C0728864|Nasal cavity
C0728864|Malignant neoplasm of nasal cavity
C0728864|malignant neoplasm of nasal cavity (diagnosis)
C0728864|nasal cavity cancer (diagnosis)
C0728864|nasal cavity cancer
C0728864|malignant nasal cavity neoplasm
C0728864|malignant tumor of nasal cavity
C0728864|Mal neo nasal cavities
C0728864|Cancer of the nasal cavity
C0728864|Malignant neoplasm of nasal cavities NOS (disorder)
C0728864|Malignant neoplasm of nasal cavities NOS
C0728864|Malignant neoplasm of nasal cavities
C0728864|Malignant tumour of nasal cavity
C0728864|Malignant tumor of nasal cavity (disorder)
C0728864|Malignant neoplasm of nasal cavity, NOS
C0728864|Malignant Nasal Cavity Tumor
C0728864|Malignant Neoplasm of the Nasal Cavity
C0728864|Malignant Tumor of the Nasal Cavity
C3887461|Head and Neck Carcinoma
C3887461|Carcinoma of Head and Neck
C3887461|Carcinoma of the Head and Neck
C0347856|Malignant neoplasm of glomus jugulare
C0347856|malignant neoplasm of glomus jugulare (diagnosis)
C0347856|malignant tumor of glomus jugulare
C0347856|Malignant neoplasm of glomus jugulare (disorder)
C0347856|glomus jugulare neoplasm malignant primary
C0347856|Primary malignant neoplasm of glomus jugulare (diagnosis)
C0347856|Primary malignant neoplasm of glomus jugulare
C0347856|Primary malignant neoplasm of glomus jugulare (disorder)
C0347856|Malignant Glomus Jugulare Neoplasm
C0347856|Malignant Glomus Jugulare Tumor
C0347856|Malignant Jugulotympanic Paraganglioma
C0347856|Malignant Neoplasm of the Glomus Jugulare
C0347856|Malignant Tumor of the Glomus Jugulare
C2350059|Cancer of Ear
C2350059|Malignant neoplasm of ear (disorder)
C2350059|Malignant neoplasm of ear
C2350059|Ear neoplasm malignant
C2350059|Malignant neoplasm of ear (diagnosis)
C2350059|neoplasm of ear malignant
C2350059|Ear Cancer
C2350059|Cancer of the Ear
C2350059|Malignant Ear Neoplasm
C2350059|Malignant Ear Tumor
C2350059|Malignant Neoplasm of the Ear
C2350059|Malignant Tumor of Ear
C2350059|Malignant Tumor of the Ear
C2350059|Neoplasm malig;ear
C2350059|malignant neosplasm of the ear
C1335975|Chordoma of Skull Base
C1335975|Chordoma of the Skull Base
C1335975|Skull Base Chordoma
C0153633|Malignant neoplasm of brain
C0153633|Malignant Brain Neoplasm
C0153633|Malignant neoplasm of brain, unspecified
C0153633|Brain, unspecified
C0153633|MALIGNANT NEOPL BRAIN
C0153633|NEOPL BRAIN MALIGNANT
C0153633|BRAIN NEOPL MALIGNANT
C0153633|Malignant neoplasm of brain (disorder)
C0153633|malignant neoplasm of brain (diagnosis)
C0153633|brain cancer (diagnosis)
C0153633|brain cancer
C0153633|malignant brain tumor
C0153633|Brain Cancers
C0153633|Cancers, Brain
C0153633|Brain Malignant Neoplasm
C0153633|Brain Malignant Neoplasms
C0153633|Brain Neoplasm, Malignant
C0153633|Malignant Brain Neoplasms
C0153633|Malignant Neoplasm, Brain
C0153633|cancer of brain
C0153633|malignant tumor of brain
C0153633|Malig neo brain NOS
C0153633|Cancer, Brain
C0153633|Brain Ca
C0153633|Malignant neoplasm of brain NOS (disorder)
C0153633|Malignant brain tumour (disorder)
C0153633|Malignant brain tumour
C0153633|Malignant neoplasm of brain NOS
C0153633|Brain--Cancer
C0153633|Malignant brain neoplasm NOS
C0153633|Brain neoplasm malignant
C0153633|Brain Neoplasms, Malignant
C0153633|Malignant Neoplasms, Brain
C0153633|Cancer of the Brain
C0153633|Neoplasms, Brain, Malignant
C0153633|Malignant neoplasm of brain, NOS
C0153633|Malignant Neoplasm of the Brain
C0153633|Malignant Tumor of the Brain
C0153633|Neoplasm malig;brain
C0153633|malignant neosplasm of the brain
C0518967|Carcinoma of head of pancreas
C0518967|Carcinoma of head of pancreas (disorder)
C0518967|pancreatic neoplasm malignant head, carcinoma
C0518967|Carcinoma of head of pancreas (diagnosis)
C0153459|Malignant neoplasm of body of pancreas
C0153459|Body of pancreas
C0153459|Mal neo pancreas body
C0153459|Ca body of pancreas
C0153459|Ca body of pancreas (disorder)
C0153459|pancreatic neoplasm malignant body
C0153459|malignant neoplasm of body of pancreas (diagnosis)
C0153459|Malignant tumor of body of pancreas
C0153459|Malignant tumour of body of pancreas
C0153459|Malignant tumor of body of pancreas (disorder)
C0153460|Malignant neoplasm of tail of pancreas
C0153460|Tail of pancreas
C0153460|Mal neo pancreas tail
C0153460|Malignant neoplasm of pancreatic tail
C0153460|Ca tail of pancreas (disorder)
C0153460|Ca tail of pancreas
C0153460|malignant neoplasm of tail of pancreas (diagnosis)
C0153460|pancreatic neoplasm malignant tail
C0153460|Malignant tumor of tail of pancreas
C0153460|Malignant tumour of tail of pancreas
C0153460|Malignant tumor of tail of pancreas (disorder)
C0153458|Malignant neoplasm of head of pancreas
C0153458|Head of pancreas
C0153458|Mal neo pancreas head
C0153458|malignant neoplasm of head of pancreas (diagnosis)
C0153458|pancreatic neoplasm malignant head
C0153458|Ca head of pancreas (disorder)
C0153458|Malignant tumour of head of pancreas
C0153458|Ca head of pancreas
C0153458|Malignant tumor of head of pancreas
C0153458|Cancer of head of pancreas
C0153458|Malignant tumor of head of pancreas (disorder)
C1328479|Carcinoma, Islet Cell
C1328479|Carcinomas, Islet Cell
C1328479|Islet Cell Carcinomas
C1328479|Islet Cell Carcinoma
C1328479|Malignant neoplasm of islets of Langerhans
C1328479|islet cell carcinoma of pancreas
C1328479|islet cell carcinoma of pancreas (diagnosis)
C1328479|islet cell carcinoma (diagnosis)
C1328479|Mal neo islet langerhans
C1328479|Carcinoma, Islet Cell [Disease/Finding]
C1328479|Islet Cell Tumor, Malignant
C1328479|High Grade Pancreatic Neuroendocrine Carcinoma
C1328479|Poorly Differentiated Pancreatic Endocrine Carcinoma
C1328479|Pancreatic NEC G3
C1328479|High-Grade Pancreatic Neuroendocrine Carcinoma
C1328479|Pancreatic Endocrine Carcinoma
C1328479|Pancreatic Neuroendocrine Carcinoma
C1328479|Pancreatic NEC
C1328479|islet cell cancer
C1328479|CARCINOMA, ISLET CELL, MALIGNANT
C1328479|pancreatic endocrine cancer
C1328479|pancreatic neoplasm malignant carcinoma endocrine pancreas
C1328479|Carcinoma of endocrine pancreas
C1328479|Carcinoma of endocrine pancreas (diagnosis)
C1328479|malignant neoplasm endocrine glands islets of langerhans
C1328479|malignant neoplasm of Islets of Langerhans (diagnosis)
C1328479|Pancreatic endocrine tumor, malignant
C1328479|Pancreatic endocrine tumour, malignant
C1328479|Malignant Islet Cell Tumor
C1328479|Malignant Pancreatic Endocrine Tumor
C1328479|Pancreatic islet cell neoplasm malignant NOS
C1328479|Malignant pancreatic islet neoplasm
C1328479|Pancreatic islet cell carcinoma
C1328479|Islet cell adenocarcinoma
C1328479|Endocrine pancreatic carcinoma
C1328479|Malignant Islet cell tumour
C1328479|Malignant tumor of Islets of Langerhans
C1328479|Malignant tumour of Islets of Langerhans
C1328479|Carcinoma of endocrine pancreas (disorder)
C1328479|Islet cell carcinoma (morphologic abnormality)
C1328479|Malignant tumor of Islets of Langerhans (disorder)
C1328479|cancer of the endocrine pancreas
C1328479|carcinoma of the endocrine pancreas
C1328479|endocrine pancreatic cancer
C1328479|carcinoma; islet cell, pancreas
C1328479|carcinoma; islet cell, unspecified site
C1328479|islet cell; carcinoma, pancreas
C1328479|islet cell; carcinoma, unspecified site
C1328479|pancreas; carcinoma, islet cell
C1328479|pancreas; islet cell carcinoma
C1328479|Malignant neoplasm of Islets of Langerhans, any part of pancreas
C0496785|Malignant neoplasm of other parts of pancreas
C0496785|Other parts of pancreas
C0496785|Primary malignant neoplasm of other parts of pancreas (disorder)
C0496785|Primary malignant neoplasm of other parts of pancreas
C0153463|Malignant neoplasm of other specified sites of pancreas
C0153463|Malig neo pancreas NEC
C0153463|Malignant neoplasm of other specified sites of pancreas (disorder)
C0153461|Pancreatic duct
C0153461|Malignant neoplasm of pancreatic duct
C0153461|Mal neo pancreatic duct
C0153461|pancreatic neoplasm malignant pancreatic duct
C0153461|malignant neoplasm of pancreatic duct (diagnosis)
C0153461|Malignant tumor of pancreatic duct
C0153461|Malignant tumour of pancreatic duct
C0153461|Malignant tumor of pancreatic duct (disorder)
C0153461|Malignant neoplasm of duct of Wirsung
C0496784|Endocrine pancreas
C0496784|Malignant neoplasm of endocrine pancreas
C0496784|malignant neoplasm of endocrine pancreas (diagnosis)
C0496784|pancreatic neoplasm malignant endocrine pancreas
C0496784|Malignant tumor of endocrine pancreas
C0496784|Malignant tumour of endocrine pancreas
C0496784|Malignant tumor of endocrine pancreas (disorder)
C0349053|Malignant neoplasm overlapping pancreas site
C0349053|Overlapping lesion of pancreas
C0349053|Malignant neoplasm of overlapping sites of pancreas
C0349053|malignant neoplasm of overlapping sites of pancreas (diagnosis)
C0349053|pancreatic neoplasm malignant overlapping sites
C0349053|Malignant neoplasm, overlapping lesion of pancreas
C0349053|Malignant neoplasm, overlapping lesion of pancreas (disorder)
C0349053|Cancer of the pancreas, overlapping sites
C0349053|Overlapping malignant neoplasm of pancreas (disorder)
C0349053|Overlapping malignant neoplasm of pancreas
C0346647|Malignant neoplasm of pancreas
C0346647|pancreatic cancer
C0346647|Malignant neoplasm of pancreas, unspecified
C0346647|Pancreas, unspecified
C0346647|malignant neoplasm of pancreas (diagnosis)
C0346647|malignant pancreatic neoplasm
C0346647|Cancers, Pancreas
C0346647|Pancreas Cancers
C0346647|Cancer, Pancreatic
C0346647|Cancers, Pancreatic
C0346647|Pancreatic Cancers
C0346647|malignant tumor of pancreas
C0346647|Malig neo pancreas NOS
C0346647|Cancer of pancreas
C0346647|Cancer, Pancreas
C0346647|Ca pancreas NOS (disorder)
C0346647|Ca pancreas NOS
C0346647|CA - Cancer of pancreas
C0346647|CA - Pancreatic cancer
C0346647|Malignant tumour of pancreas
C0346647|Malignant neoplasm of pancreas NOS
C0346647|Malignant neoplasm of pancreas NOS (disorder)
C0346647|Pancreas--Cancer
C0346647|Pancreas cancer
C0346647|Neoplasm of the pancreas
C0346647|Cancer of the pancreas
C0346647|Neoplasia of the pancreas
C0346647|Pancreas neoplasm malignant
C0346647|Malignant neoplasm of pancreas, part unspecified
C0346647|Malignant tumor of pancreas (disorder)
C0346647|Malignant neoplasm of pancreas, NOS
C0346647|Malignant Neoplasm of the Pancreas
C0346647|Neoplasm malig;pancreas
C0346647|malignant neosplasm of the pancreas
C2007079|carcinosarcoma of pancreas (diagnosis)
C2007079|carcinosarcoma of pancreas
C0235974|Pancreatic carcinoma
C0235974|carcinoma of pancreas (diagnosis)
C0235974|carcinoma of pancreas
C0235974|Carcinoma;pancreas
C0235974|PANCREATIC CANCER
C0235974|Pancreatic Acinar Carcinoma
C0235974|Carcinoma of pancreas (disorder)
C0235974|exocrine cancer
C0235974|Pancreatic cancer (not Islets)
C0235974|Pancreatic cancer (excluding Islets), NOS
C0235974|Pancreatic carcinoma NOS
C0235974|Pancreas carcinoma
C0235974|Cancer of Pancreas
C0235974|Cancer of the Pancreas
C0235974|Pancreas Cancer
C0235974|Exocrine Pancreas Carcinoma
C0235974|Carcinoma of the Pancreas
C2205484|malignant small cell neoplasm of pancreas (diagnosis)
C2205484|pancreatic neoplasm malignant small cell type
C2205484|malignant small cell neoplasm of pancreas
C2011344|giant cell type neoplasm of pancreas
C2011344|giant cell type neoplasm of pancreas (diagnosis)
C2018676|spindle cell type neoplasm of pancreas (diagnosis)
C2018676|spindle cell type neoplasm of pancreas
C2018676|pancreatic neoplasm malignant spindle cell type
C2075636|clear cell type neoplasm of pancreas
C2075636|pancreatic neoplasm malignant clear cell type
C2075636|clear cell type neoplasm of pancreas (diagnosis)
C3536762|malignant carcinoid tumor of pancreas
C3536762|malignant carcinoid tumor of pancreas (diagnosis)
C3536762|Malignant carcinoid tumor of pancreas (disorder)
C3536762|Malignant carcinoid tumour of pancreas
C1096346|sarcoma of pancreas (diagnosis)
C1096346|sarcoma of pancreas
C1096346|Pancreatic sarcoma
C1096346|Sarcoma of the Pancreas
C2205511|myosarcoma of pancreas (diagnosis)
C2205511|myosarcoma of pancreas
C2205516|malignant lymphoma of pancreas (diagnosis)
C2205516|malignant lymphoma of pancreas
C2205519|malignant plasmacytoma of pancreas
C2205519|malignant plasmacytoma of pancreas (diagnosis)
C2205521|malignant mastocytosis of pancreas (diagnosis)
C2205521|malignant mastocytosis of pancreas
C0281361|Pancreatic adenocarcinoma
C0281361|adenocarcinoma of pancreas
C0281361|adenocarcinoma of pancreas (diagnosis)
C0281361|Adenocarcinoma pancreas
C0281361|Adenocarcinoma of pancreas (disorder)
C0281361|Adenocarcinoma - pancreas
C0281361|Adenocarcinoma of the pancreas
C0281361|Pancreas Adenocarcinoma
C2062546|microadenomatosis of pancreas (diagnosis)
C2062546|microadenomatosis of pancreas
C2062546|pancreatic microadenomatosis
C0086768|Cholera, Pancreatic
C0086768|Verner Morrison Syndrome
C0086768|Syndrome, Verner-Morrison
C0086768|Verner-Morrison syndrome due to pancreatic neoplasm
C0086768|Verner-Morrison syndrome due to pancreatic neoplasm (diagnosis)
C0086768|pancreatic cholera (WDHA syndrome)
C0086768|WDHA Syndromes
C0086768|Excessive vasoactive intestinal peptide secretion (disorder)
C0086768|Excessive vasoactive intestinal peptide secretion
C0086768|Verner-Morrison syndrome
C0086768|Vipoma Syndrome
C0086768|Watery Diarrhea Syndrome
C0086768|WDHH
C0086768|Watery Diarrhea, Hypokalemia, and Achlorhydria Syndrome
C0086768|Watery Diarrhea with Hypokalemic Alkalosis
C0086768|WDHA
C0086768|WDHA Syndrome
C0086768|Syndrome, Vipoma
C0086768|Pseudopancreatic cholera syndrome
C0086768|Pancreatic cholera
C0086768|Werner Morrison syndrome
C0086768|Pseudopancreatic cholera syndrome (disorder)
C0086768|Verner-Morrison syndrome (disorder)
C0086768|islet cell WDHA syndrome
C0086768|pancreatic WDHA syndrome
C0086768|Excessive vasoactive intestinal peptide secretion [Ambiguous]
C1389637|malignant beta cell tumor of pancreas (diagnosis)
C1389637|malignant beta cell tumor of pancreas
C1389637|malignant insulinoma of pancreas
C1389637|malignant pancreatic beta cell tumor
C1389637|malignant insulinoma of pancreas (diagnosis)
C1389637|beta-cell; tumor, malignant, pancreas
C1389637|insulinoma; malignant, pancreas
C1389637|malignant; insulinoma, pancreas
C1389637|pancreas; beta-cell tumor, malignant
C1389637|pancreas; insulinoma, malignant
C1389637|pancreas; malignant insulinoma
C1389637|pancreas; tumor, beta-cell, malignant
C1389637|tumor; beta-cell, malignant, pancreas
C1335315|serous cystadenocarcinoma of pancreas
C1335315|serous cystadenocarcinoma of pancreas (diagnosis)
C1335315|Pancreatic Serous Cystadenocarcinoma
C1335315|Serous Cystadenocarcinoma of the Pancreas
C2063876|invasive mucinous cystadenocarcinoma of pancreas (diagnosis)
C2063876|invasive mucinous cystadenocarcinoma of pancreas
C1335304|intraductal papillary-mucinous carcinoma of pancreas (diagnosis)
C1335304|intraductal papillary-mucinous carcinoma of pancreas
C1335304|Pancreatic Intraductal Papillary-Colloid Carcinoma
C1335304|Pancreatic Intraductal Papillary-Colloidal Carcinoma
C1335304|Intraductal Papillary-Colloidal Carcinoma of the Pancreas
C1335304|Intraductal Papillary-Mucinous Carcinoma of the Pancreas
C1335304|Intraductal Papillary-Colloid Carcinoma of Pancreas
C1335304|Intraductal Papillary-Colloid Carcinoma of the Pancreas
C1335304|Intraductal Papillary-Colloidal Carcinoma of Pancreas
C1335304|Pancreatic Intraductal Papillary-Mucinous Carcinoma
C2063878|mixed acinar-endocrine carcinoma of pancreas (diagnosis)
C2063878|mixed acinar-endocrine carcinoma of pancreas
C2063878|Mucinous Carcinoid Tumor of the Pancreas
C2063878|Mixed Carcinoid-Adenocarcinoma of the Pancreas
C2063878|Mixed Acinar-Endocrine Carcinoma of the Pancreas
C2063878|Mixed Acinar-Neuroendocrine Carcinoma of the Pancreas
C2063878|ACINAR-ISLET CELL TUMOR, MALIGNANT
C0334489|pancreatoblastoma (diagnosis)
C0334489|pancreatoblastoma
C0334489|Pancreatoblastoma (disorder)
C0334489|[M]Pancreatoblastoma
C0334489|[M] Pancreatoblastoma
C0334489|Pancreatoblastoma (morphologic abnormality)
C2205494|scirrhous adenocarcinoma of pancreas (diagnosis)
C2205494|scirrhous adenocarcinoma of pancreas
C2205494|pancreatic neoplasm adenocarcinoma scirrhous
C2037343|pancreatic neoplasm adenocarcinoma superficial spreading
C2037343|superficial spreading adenocarcinoma of pancreas (diagnosis)
C2037343|superficial spreading adenocarcinoma of pancreas
C2205495|basal cell adenocarcinoma of pancreas (diagnosis)
C2205495|basal cell adenocarcinoma of pancreas
C2033127|papillary adenocarcinoma of pancreas (diagnosis)
C2033127|papillary adenocarcinoma of pancreas
C2189643|villous adenocarcinoma of pancreas (diagnosis)
C2189643|villous adenocarcinoma of pancreas
C2205497|adenocarcinoma in tubulovillous adenoma of pancreas
C2205497|adenocarcinoma in tubulovillous adenoma of pancreas (diagnosis)
C2205498|adenocarcinoma in adenomatous polyp of pancreas (diagnosis)
C2205498|adenocarcinoma in adenomatous polyp of pancreas
C2205499|mucin-producing adenocarcinoma of pancreas (diagnosis)
C2205499|mucin-producing adenocarcinoma of pancreas
C2033012|intraductal papillary adenocarcinoma of pancreas with invasion
C2033012|intraductal papillary adenocarcinoma of pancreas with invasion (diagnosis)
C2205500|adenocarcinoma of pancreas with metaplasia (diagnosis)
C2205500|pancreatic adenocarcinoma with metaplasia
C2205500|adenocarcinoma of pancreas with metaplasia
C2205501|adenocarcinoma of pancreas with squamous metaplasia (diagnosis)
C2205501|adenocarcinoma of pancreas with squamous metaplasia
C2205501|pancreatic adenocarcinoma with squamous metaplasia
C2033013|adenocarcinoma with cartilaginous or osseous metaplasia of pancreas
C2033013|adenocarcinoma of pancreas with cartilaginous and osseous metaplasia
C2033013|adenocarcinoma of pancreas with cartilaginous and osseous metaplasia (diagnosis)
C2033013|pancreatic adenocarcinoma with cartilaginous or osseous metaplasia
C2033013|pancreatic adenocarcinoma with cartilaginous and osseous metaplasia
C2205502|pancreatic adenocarcinoma metaplastic spindle cell
C2205502|pancreatic adenocarcinoma with spindle cell metaplasia
C2205502|adenocarcinoma of pancreas with spindle cell metaplasia (diagnosis)
C2205502|adenocarcinoma of pancreas with spindle cell metaplasia
C2205503|pancreatic adenocarcinoma with apocrine metaplasia
C2205503|adenocarcinoma of pancreas with apocrine metaplasia (diagnosis)
C2205503|adenocarcinoma of pancreas with apocrine metaplasia
C2033014|adenocarcinoma of pancreas with neuroendocrine differentiation (diagnosis)
C2033014|adenocarcinoma of pancreas with neuroendocrine differentiation
C2033014|pancreatic adenocarcinoma with neuroendocrine differentiation
C2030694|hepatoid adenocarcinoma of pancreas
C2030694|hepatoid adenocarcinoma of pancreas (diagnosis)
C2170821|tubular adenocarcinoma of pancreas (diagnosis)
C2170821|tubular adenocarcinoma of pancreas
C2075534|clear cell adenocarcinoma of pancreas
C2075534|clear cell adenocarcinoma of pancreas (diagnosis)
C2063871|mucinous adenocarcinoma of pancreas
C2063871|mucinous adenocarcinoma of pancreas (diagnosis)
C2033034|noninvasive intraductal papillary-mucinous carcinoma of pancreas (diagnosis)
C2033034|noninvasive intraductal papillary-mucinous carcinoma of pancreas
C1518871|intraductal papillary-mucinous carcinoma of the pancreas invasive
C1518871|invasive intraductal papillary-mucinous carcinoma of pancreas
C1518871|intraductal papillary-mucinous carcinoma of the pancreas invasive (diagnosis)
C1518871|Pancreatic Intraductal Papillary-Mucinous Neoplasm with an Associated Invasive Carcinoma
C1518871|Pancreatic Invasive Intraductal Papillary-Mucinous Carcinoma
C1518871|Pancreatic Intraductal Papillary Mucinous Neoplasm with an Associated Invasive Carcinoma
C1336861|undifferentiated carcinoma of pancreas (diagnosis)
C1336861|undifferentiated carcinoma of pancreas
C1336861|Pancreatic Carcinosarcoma
C1336861|Pleomorphic Large Cell Pancreatic Carcinoma
C1336861|Sarcomatoid Pancreatic Carcinoma
C1336861|Undifferentiated (Anaplastic) Pancreatic Carcinoma
C1336861|Spindle Cell Pancreatic Carcinoma
C1336861|Undifferentiated Pancreatic Carcinoma
C1336861|Undifferentiated Carcinoma of the Pancreas
C2033249|papillary cystadenocarcinoma of pancreas (diagnosis)
C2033249|papillary cystadenocarcinoma of pancreas
C2033261|papillary mucinous cystadenocarcinoma of pancreas (diagnosis)
C2033261|papillary mucinous cystadenocarcinoma of pancreas
C2106547|comedocarcinoma of pancreas
C2106547|comedocarcinoma of pancreas (diagnosis)
C2205496|adenocarcinoma in villous adenoma of pancreas
C2205496|adenocarcinoma in villous adenoma of pancreas (diagnosis)
C2018503|spindle cell sarcoma of pancreas
C2018503|spindle cell sarcoma of pancreas (diagnosis)
C2011317|giant cell sarcoma of pancreas
C2011317|giant cell sarcoma of pancreas (diagnosis)
C2205507|small cell sarcoma of pancreas (diagnosis)
C2205507|small cell sarcoma of pancreas
C2205508|epithelioid sarcoma of pancreas (diagnosis)
C2205508|epithelioid sarcoma of pancreas
C2188140|undifferentiated sarcoma of pancreas
C2188140|undifferentiated sarcoma of pancreas (diagnosis)
C2182952|desmoplastic small round cell sarcoma of pancreas
C2182952|desmoplastic small round cell sarcoma of pancreas (diagnosis)
C2046335|histiocytic sarcoma of pancreas
C2046335|histiocytic sarcoma of pancreas (diagnosis)
C2111172|Langerhans cell sarcoma of pancreas (diagnosis)
C2111172|Langerhans cell sarcoma of pancreas
C2077758|interdigitating dendritic cell sarcoma of pancreas
C2077758|interdigitating dendritic cell sarcoma of pancreas (diagnosis)
C2205510|follicular dendritic cell sarcoma of pancreas
C2205510|follicular dendritic cell sarcoma of pancreas (diagnosis)
C2205513|angiomyosarcoma of pancreas (diagnosis)
C2205513|angiomyosarcoma of pancreas
C1409081|mixed islet cell and exocrine adenocarcinoma of pancreas (diagnosis)
C1409081|mixed islet cell and exocrine adenocarcinoma of pancreas
C1409081|pancreas; adenocarcinoma islet cell, with exocrine mixed
C2033018|noninfiltrating intraductal carcinoma of pancreas (diagnosis)
C2033018|noninfiltrating intraductal carcinoma of pancreas
C2033017|noninfiltrating intracystic carcinoma of pancreas (diagnosis)
C2033017|noninfiltrating intracystic carcinoma of pancreas
C2033016|intraductal micropapillary carcinoma of pancreas (diagnosis)
C2033016|intraductal micropapillary carcinoma of pancreas
C2205485|malignant epithelioma of pancreas (diagnosis)
C2205485|malignant epithelioma of pancreas
C2111650|large cell carcinoma of pancreas
C2111650|large cell carcinoma of pancreas (diagnosis)
C2111737|large cell neuroendocrine carcinoma of pancreas (diagnosis)
C2111737|large cell neuroendocrine carcinoma of pancreas
C2111651|pancreatic neoplasm carcinoma large cell with rhabdoid phenotype
C2111651|large cell carcinoma of pancreas with rhabdoid phenotype (diagnosis)
C2111651|large cell carcinoma of pancreas with rhabdoid phenotype
C2012101|glassy cell carcinoma of pancreas
C2012101|glassy cell carcinoma of pancreas (diagnosis)
C2082450|pleomorphic carcinoma of pancreas (diagnosis)
C2082450|pleomorphic carcinoma of pancreas
C2011260|giant cell carcinoma of pancreas
C2011260|giant cell carcinoma of pancreas (diagnosis)
C2018400|spindle cell carcinoma of pancreas
C2018400|spindle cell carcinoma of pancreas (diagnosis)
C2011225|giant cell and spindle cell carcinoma of pancreas
C2011225|giant cell and spindle cell carcinoma of pancreas (diagnosis)
C2142930|pseudosarcomatous carcinoma of pancreas
C2142930|pseudosarcomatous carcinoma of pancreas (diagnosis)
C2111812|polygonal cell carcinoma of pancreas
C2111812|polygonal cell carcinoma of pancreas (diagnosis)
C2205486|small cell carcinoma of pancreas
C2205486|small cell carcinoma of pancreas (diagnosis)
C2009884|fusiform type small cell carcinoma of pancreas (diagnosis)
C2009884|fusiform type small cell carcinoma of pancreas
C2033227|papillary carcinoma of pancreas
C2033227|papillary carcinoma of pancreas (diagnosis)
C2033304|papillary squamous cell carcinoma of pancreas
C2033304|papillary squamous cell carcinoma of pancreas (diagnosis)
C2189356|verrucous carcinoma of pancreas
C2189356|verrucous carcinoma of pancreas (diagnosis)
C2675993|squamous cell carcinoma of pancreas (diagnosis)
C2675993|squamous cell carcinoma of pancreas
C2675993|Pancreatic squamous cell carcinoma
C2675993|Squamous cell carcinoma of the pancreas
C2109314|keratinizing squamous cell carcinoma of pancreas
C2109314|keratinizing squamous cell carcinoma of pancreas (diagnosis)
C2205487|pancreatic carcinoma squamous cell large cell nonkeratinizing
C2205487|nonkeratinizing large cell squamous carcinoma cell of pancreas
C2205487|nonkeratinizing large cell squamous carcinoma cell of pancreas (diagnosis)
C2205488|nonkeratinizing small cell squamous cell carcinoma of pancreas (diagnosis)
C2205488|nonkeratinizing small cell squamous cell carcinoma of pancreas
C2018561|spindle cell squamous cell carcinoma of pancreas (diagnosis)
C2018561|spindle cell squamous cell carcinoma of pancreas
C2205489|adenoid squamous cell carcinoma of pancreas (diagnosis)
C2205489|adenoid squamous cell carcinoma of pancreas
C2205490|microinvasive squamous cell carcinoma of pancreas
C2205490|microinvasive squamous cell carcinoma of pancreas (diagnosis)
C2019489|pancreatic neoplasm carcinoma squamous cell with horn formation
C2019489|squamous cell carcinoma of pancreas with horn formation
C2019489|squamous cell carcinoma with horn formation of pancreas
C2019489|squamous cell carcinoma of pancreas with horn formation (diagnosis)
C2017452|solid carcinoma of pancreas
C2017452|solid carcinoma of pancreas (diagnosis)
C2007049|carcinoma simplex of pancreas (diagnosis)
C2007049|carcinoma simplex of pancreas
C2205491|mucoepidermoid carcinoma of pancreas (diagnosis)
C2205491|mucoepidermoid carcinoma of pancreas
C2076527|infiltrating ductal carcinoma of pancreas
C2076527|infiltrating ductal carcinoma of pancreas (diagnosis)
C2078054|intracystic carcinoma of pancreas
C2078054|intracystic carcinoma of pancreas (diagnosis)
C2047536|hypersecretory cystic carcinoma of pancreas
C2047536|hypersecretory cystic carcinoma of pancreas (diagnosis)
C2205492|medullary carcinoma of pancreas (diagnosis)
C2205492|medullary carcinoma of pancreas
C2182972|duct carcinoma, desmoplastic type, of pancreas
C2182972|duct carcinoma, desmoplastic type, of pancreas (diagnosis)
C2076531|infiltrating ductular carcinoma of pancreas (diagnosis)
C2076531|infiltrating ductular carcinoma of pancreas
C2205493|epithelial-myoepithelial carcinoma of pancreas (diagnosis)
C2205493|epithelial-myoepithelial carcinoma of pancreas
C2205506|neuroendocrine carcinoma of pancreas
C2205506|neuroendocrine carcinoma of pancreas (diagnosis)
C2205514|embryonal carcinosarcoma of pancreas (diagnosis)
C2205514|embryonal carcinosarcoma of pancreas
C3469525|pancreatic cancer susceptibility
C3469525|pancreatic cancer susceptibility (diagnosis)
C3469525|PANCREATIC CANCER, SUSCEPTIBILITY TO
C1335317|signet ring cell carcinoma of pancreas
C1335317|signet ring cell carcinoma of pancreas (diagnosis)
C1335317|Pancreatic Signet Ring Cell Carcinoma
C1335317|Signet Ring Cell Carcinoma of the Pancreas
C1335299|adenosquamous carcinoma of pancreas
C1335299|adenosquamous carcinoma of pancreas (diagnosis)
C1335299|Pancreatic Adenoacanthoma
C1335299|Pancreatic Mucoepidermoid Carcinoma
C1335299|Pancreatic Mixed Squamous and Adenocarcinoma
C1335299|Adenosquamous Carcinoma of the Pancreas
C1335299|Pancreatic Adenosquamous Carcinoma
C2063872|anaplastic carcinoma of pancreas
C2063872|anaplastic carcinoma of pancreas (diagnosis)
C2007059|carcinoma of pancreas with osteoclast-like giant cells
C2007059|carcinoma of pancreas with osteoclast-like giant cells (diagnosis)
C2007059|pancreatic carcinoma with osteoclast-like giant cells
C2007059|Pancreatic Osteoclast-Like Giant Cell Carcinoma
C2007059|Undifferentiated Pancreatic Carcinoma with Osteoclast-Like Giant Cells
C2007059|Osteoclast-like Giant Cell Neoplasm of Pancreas
C2007059|Osteoclast-like Giant Cell Neoplasm of the Pancreas
C0279661|acinar cell carcinoma of pancreas
C0279661|acinar cell carcinoma of pancreas (diagnosis)
C0279661|acinar cell adenocarcinoma of the pancreas
C0279661|adenocarcinoma, acinar cell, pancreatic
C0279661|pancreas cancer, acinar cell adenocarcinoma
C0279661|pancreatic cancer, acinar cell adenocarcinoma
C0279661|Acinar Cell Adenocarcinoma of Pancreas
C0279661|Acinar Cell Carcinoma of the Pancreas
C0279661|Pancreas Acinar Cell Adenocarcinoma
C0279661|Pancreatic Acinar Cell Adenocarcinoma
C0279661|Pancreatic Acinar Cell Carcinoma
C1336029|solid pseudopapillary carcinoma of pancreas (diagnosis)
C1336029|solid pseudopapillary carcinoma of pancreas
C1336029|Pancreatic Solid Pseudopapillary Carcinoma
C1336029|Solid Pseudopapillary Carcinoma of the Pancreas
C3472164|Primary adenocarcinoma of pancreas (disorder)
C3472164|Primary adenocarcinoma of pancreas
C3532881|Intraductal papillary mucinous carcinoma in situ of pancreas (disorder)
C3532881|Intraductal papillary mucinous neoplasm with high grade dysplasia
C3532881|Intraductal papillary mucinous carcinoma in situ of pancreas
C0153454|Ampulla of Vater
C0153454|Malignant neoplasm of ampulla of Vater
C0153454|Mal neo ampulla of vater
C0153454|malignant neoplasm ampulla of vater
C0153454|malignant neoplasm ampulla of vater (diagnosis)
C0153454|Malignant tumour of ampulla of Vater
C0153454|Malignant tumor of ampulla of Vater
C0153454|Malignant tumor of ampulla of Vater (disorder)
C0153454|Malignant Ampulla of Vater Neoplasm
C0153454|Malignant Ampulla of Vater Tumor
C0153454|Malignant Neoplasm of the Ampulla of Vater
C0153454|Malignant Tumor of the Ampulla of Vater
C1282477|pancreatic malignant neoplasm, local recurrence
C1282477|local recurrence of malignant neoplasm of pancreas
C1282477|local recurrence of malignant neoplasm of pancreas (diagnosis)
C1282477|Local recurrence of malignant tumor of pancreas (disorder)
C1282477|Local recurrence of malignant tumor of pancreas
C1282477|Local recurrence of malignant tumour of pancreas
C0346976|Metastatic Neoplasm to the Pancreas
C0346976|Metastases to pancreas
C0346976|Secondary malignant neoplasm of pancreas
C0346976|pancreatic malignant neoplasm secondary
C0346976|Secondary malignant neoplasm of pancreas (diagnosis)
C0346976|Metastatic Malignant Neoplasm to the Pancreas
C0346976|Metastatic Malignant Neoplasm in the Pancreas
C0346976|Cancer metastatic to pancreas
C0346976|Malignant neoplasm of pancreas metastatic
C0346976|Pancreas neoplasm malignant metastatic
C0346976|Pancreatic cancer metastatic
C0346976|Metastasis to pancreas
C0346976|Pancreatic metastasis
C0346976|Secondary malignant deposit in pancreas
C0346976|Metastatic malignant neoplasm to pancreas
C0346976|Secondary malignant neoplasm of pancreas (disorder)
C0346976|metastatic pancreas cancer
C0346976|metastatic pancreatic cancer
C0346976|pancreas cancer, metastatic
C0346976|pancreatic cancer, metastatic
C0346976|Metastatic malignant neoplasm to pancreas, NOS
C0346976|Secondary malignant neoplasm of pancreas, NOS
C0346976|Metastatic Cancer to the Pancreas
C0346976|Metastatic Tumor to the Pancreas
C0346976|Secondary Cancer to the Pancreas
C0346976|Secondary Malignant Neoplasm to the Pancreas
C0346976|Secondary Malignant Tumor to the Pancreas
C0346648|malignant neoplasm of exocrine pancreas
C0346648|malignant neoplasm of exocrine pancreas (diagnosis)
C0346648|pancreatic neoplasm malignant exocrine
C0346648|Malignant tumor of exocrine pancreas
C0346648|Malignant tumour of exocrine pancreas
C0346648|Pancreatic exocrine cancer
C0346648|Malignant tumor of exocrine pancreas (disorder)
C0346648|Malignant Exocrine Pancreas Neoplasm
C0346648|Malignant Exocrine Pancreas Tumor
C0346648|Malignant Neoplasm of the Exocrine Pancreas
C0346648|Malignant Tumor of the Exocrine Pancreas
C0346650|malignant neoplasm of ectopic tissue of pancreas
C0346650|pancreatic neoplasm malignant of ectopic tissue
C0346650|malignant neoplasm of ectopic tissue of pancreas (diagnosis)
C0346650|Malignant neoplasm of ectopic pancreatic tissue
C0346650|Malignant neoplasm of ectopic pancreatic tissue (disorder)
C0346651|Malignant neoplasm of specified site of pancreas NOS (disorder)
C0346651|Malignant neoplasm of specified site of pancreas NOS
C1299297|Primary malignant neoplasm of pancreas
C1299297|Primary malignant neoplasm of pancreas (disorder)
C1299297|pancreatic malignant neoplasm primary
C1299297|Primary malignant neoplasm of pancreas (diagnosis)
C2205515|malignant myoepithelioma of pancreas
C2205515|malignant myoepithelioma of pancreas (diagnosis)
C2205515|myoepithelioma of pancreas
C3836561|pancreatic cancer, somatic
C3836561|pancreatic cancer, somatic (diagnosis)
C1851697|Pancreatic islet cell adenoma
C4030391|biopsy of pancreas showed villous adenocarcinoma (procedure)
C4030391|biopsy of pancreas showed villous adenocarcinoma
C4030391|biopsy pancreas malignant neoplasm adenocarcinoma villous
C4030470|biopsy of pancreas showed malignant insulinoma (procedure)
C4030470|biopsy pancreas malignant neoplasm carcinoma islet cell insulinoma
C4030470|biopsy of pancreas showed malignant insulinoma
C4030411|biopsy of pancreas showed small cell sarcoma (procedure)
C4030411|biopsy of pancreas showed small cell sarcoma
C4030411|biopsy pancreas malignant neoplasm sarcoma small cell
C4030557|biopsy of pancreas showed adenoid squamous cell carcinoma (procedure)
C4030557|biopsy of pancreas showed adenoid squamous cell carcinoma
C4030557|biopsy pancreas malignant neoplasm carcinoma squamous cell adenoid
C4030400|biopsy of pancreas showed squamous cell carcinoma (procedure)
C4030400|biopsy of pancreas showed squamous cell carcinoma
C4030400|biopsy pancreas malignant neoplasm carcinoma squamous cell
C4030506|biopsy pancreas malignant neoplasm lymphoma hodgkin's
C4030506|biopsy of pancreas showed Hodgkin's lymphoma
C4030506|biopsy of pancreas showed Hodgkin's lymphoma (procedure)
C4030416|biopsy pancreas malignant neoplasm adenocarcinoma scirrhous
C4030416|biopsy of pancreas showed scirrhous adenocarcinoma (procedure)
C4030416|biopsy of pancreas showed scirrhous adenocarcinoma
C4030419|biopsy pancreas malig lymphoma precursor cell lymphoblastic t-cell
C4030419|biopsy of pancreas showed precursor T-cell lymphoblastic lymphoma (procedure)
C4030419|biopsy of pancreas showed precursor T-cell lymphoblastic lymphoma
C4030510|biopsy of pancreas showed grade 3 follicular lymphoma
C4030510|biopsy of pancreas showed grade 3 follicular lymphoma (procedure)
C4030510|biopsy pancreas malignant neoplasm lymphoma follicular grade 3
C4030482|biopsy of pancreas showed leiomyosarcoma (procedure)
C4030482|biopsy pancreas malignant neoplasm myosarcoma leiomyosarcoma
C4030482|biopsy of pancreas showed leiomyosarcoma
C4030533|biopsy of pancreas showed carcinosarcoma (procedure)
C4030533|biopsy of pancreas showed carcinosarcoma
C4030533|biopsy pancreas malignant neoplasm carcinosarcoma
C4030481|biopsy of pancreas showed lymphocyte-rich Hodgkin's lymphoma
C4030481|biopsy pancreas malig neoplasm lymphoma hodgkin's lymphocyte-rich
C4030481|biopsy of pancreas showed lymphocyte-rich Hodgkin's lymphoma (procedure)
C4030452|biopsy pancreas malig neoplasm lymphoma hodgkin's mixed cellularity
C4030452|biopsy of pancreas showed mixed cellularity Hodgkin's lymphoma
C4030452|biopsy of pancreas showed mixed cellularity Hodgkin's lymphoma (procedure)
C4030505|biopsy pancreas malig lymphoma hodgkin's nodular sclerosis grade 1
C4030505|biopsy of pancreas showed Hodgkin's lymphoma with grade 1 nodular sclerosis (procedure)
C4030505|biopsy of pancreas showed Hodgkin's lymphoma with grade 1 nodular sclerosis
C4030497|biopsy of pancreas showed infiltrating ductular carcinoma
C4030497|biopsy pancreas malignant neoplasm carcinoma infiltrating ductular
C4030497|biopsy of pancreas showed infiltrating ductular carcinoma (procedure)
C4030565|biopsy of pancreas showed adenocarcinoma in tubulovillous adenoma (procedure)
C4030565|biopsy pancreas malig neoplasm adenocarcinoma in tubulovillous adenoma
C4030565|biopsy of pancreas showed adenocarcinoma in tubulovillous adenoma
C4030562|biopsy of pancreas showed adenocarcinoma with cartilaginous and osseous metaplasia (procedure)
C4030562|biopsy of pancreas showed adenocarcinoma with cartilaginous and osseous metaplasia
C4030562|biopsy pancreas malig adenocarcinoma metaplastic cartilaginous & osseous
C4030479|biopsy pancreas malig neoplasm sarcoma desmoplastic small round cell
C4030479|biopsy of pancreas showed malignant desmoplastic small round cell tumor (procedure)
C4030479|biopsy of pancreas showed malignant desmoplastic small round cell tumor
C4030516|biopsy of pancreas showed giant cell carcinoma
C4030516|biopsy of pancreas showed giant cell carcinoma (procedure)
C4030516|biopsy pancreas malignant neoplasm carcinoma giant cell
C4030473|biopsy of pancreas showed malignant glucagonoma
C4030473|biopsy of pancreas showed malignant glucagonoma (procedure)
C4030473|biopsy pancreas malignant neoplasm carcinoma islet cell glucagonoma
C4030504|biopsy of pancreas showed Hodgkin's lymphoma with grade 2 nodular sclerosis
C4030504|biopsy pancreas malig lymphoma hodgkin's nodular sclerosis grade 2
C4030504|biopsy of pancreas showed Hodgkin's lymphoma with grade 2 nodular sclerosis (procedure)
C4030456|biopsy pancreas malignant neoplasm lymphoma mature t-cell
C4030456|biopsy of pancreas showed mature T-cell lymphoma (procedure)
C4030456|biopsy of pancreas showed mature T-cell lymphoma
C4030487|biopsy of pancreas showed Langerhans cell sarcoma
C4030487|biopsy of pancreas showed Langerhans cell sarcoma (procedure)
C4030487|biopsy pancreas malignant neoplasm sarcoma langerhans cell
C4030498|biopsy of pancreas showed infiltrating duct carcinoma (procedure)
C4030498|biopsy of pancreas showed infiltrating duct carcinoma
C4030498|biopsy pancreas malignant neoplasm carcinoma infiltrating duct
C4030488|biopsy of pancreas showed keratinizing squamous cell carcinoma (procedure)
C4030488|biopsy pancreas malignant neoplasm carcinoma squamous cell keratinizing
C4030488|biopsy of pancreas showed keratinizing squamous cell carcinoma
C4030532|biopsy pancreas malignant neoplasm adenocarcinoma clear cell
C4030532|biopsy of pancreas showed clear cell adenocarcinoma
C4030532|biopsy of pancreas showed clear cell adenocarcinoma (procedure)
C4030417|biopsy of pancreas showed sarcoma (procedure)
C4030417|biopsy pancreas malignant neoplasm sarcoma
C4030417|biopsy of pancreas showed sarcoma
C4030484|biopsy of pancreas showed large cell neuroendocrine carcinoma (procedure)
C4030484|biopsy pancreas malig neoplasm carcinoma large cell neuroendocrine
C4030484|biopsy of pancreas showed large cell neuroendocrine carcinoma
C4030392|biopsy of pancreas showed verrucous carcinoma
C4030392|biopsy of pancreas showed verrucous carcinoma (procedure)
C4030392|biopsy pancreas malignant neoplasm carcinoma verrucous
C4030422|biopsy of pancreas showed polygonal cell carcinoma
C4030422|biopsy of pancreas showed polygonal cell carcinoma (procedure)
C4030422|biopsy pancreas malignant neoplasm carcinoma polygonal cell
C4030527|biopsy pancreas malignant neoplasm carcinoma cystic hypersecretory
C4030527|biopsy of pancreas showed cystic hypersecretory carcinoma (procedure)
C4030527|biopsy of pancreas showed cystic hypersecretory carcinoma
C4030513|biopsy of pancreas showed goblet cell carcinoid tumor (procedure)
C4030513|biopsy of pancreas showed goblet cell carcinoid tumor
C4030513|biopsy pancreas malignant neoplasm carcinoid tumor goblet cell
C4030409|biopsy of pancreas showed solid carcinoma (procedure)
C4030409|biopsy of pancreas showed solid carcinoma
C4030409|biopsy pancreas malignant neoplasm carcinoma solid
C4030450|biopsy pancreas malignant neoplasm adenocarcinoma mucinous
C4030450|biopsy of pancreas showed mucinous adenocarcinoma
C4030450|biopsy of pancreas showed mucinous adenocarcinoma (procedure)
C4030521|biopsy of pancreas showed epithelioid sarcoma
C4030521|biopsy pancreas malignant neoplasm sarcoma epithelioid
C4030521|biopsy of pancreas showed epithelioid sarcoma (procedure)
C4030571|biopsy of pancreas showed adenocarcinoma
C4030571|biopsy of pancreas showed adenocarcinoma (procedure)
C4030571|biopsy pancreas malignant neoplasm adenocarcinoma
C4030425|biopsy of pancreas showed papillary squamous cell carcinoma
C4030425|biopsy of pancreas showed papillary squamous cell carcinoma (procedure)
C4030425|biopsy pancreas malignant neoplasm carcinoma papillary squamous cell
C4030480|biopsy of pancreas showed malignant clear cell type neoplasm
C4030480|biopsy of pancreas showed malignant clear cell type neoplasm (procedure)
C4030480|biopsy pancreas malignant neoplasm clear cell type
C4030426|biopsy of pancreas showed papillary mucinous cystadenocarcinoma (procedure)
C4030426|biopsy of pancreas showed papillary mucinous cystadenocarcinoma
C4030426|biopsy pancreas malignant neoplasm cystadenocarcinoma papillary mucinous
C4030460|biopsy of pancreas showed malignant somatostatinoma (procedure)
C4030460|biopsy pancreas malig neoplasm carcinoma islet cell somatostatinoma
C4030460|biopsy of pancreas showed malignant somatostatinoma
C4030458|biopsy pancreas malignant neoplasm lymphoma marginal zone b-cell
C4030458|biopsy of pancreas showed marginal zone B-cell lymphoma
C4030458|biopsy of pancreas showed marginal zone B-cell lymphoma (procedure)
C4030573|biopsy of pancreas showed acinar cell cystadenocarcinoma
C4030573|biopsy of pancreas showed acinar cell cystadenocarcinoma (procedure)
C4030573|biopsy pancreas malignant neoplasm acinar cell cystadenocarcinoma
C4030441|biopsy of pancreas showed neuroendocrine carcinoma
C4030441|biopsy of pancreas showed neuroendocrine carcinoma (procedure)
C4030441|biopsy pancreas malignant neoplasm carcinoma neuroendocrine
C4030396|biopsy of pancreas showed superficial spreading adenocarcinoma (procedure)
C4030396|biopsy of pancreas showed superficial spreading adenocarcinoma
C4030396|biopsy pancreas malignant neoplasm adenocarcinoma superficial spreading
C4030563|biopsy of pancreas showed adenocarcinoma with apocrine metaplasia
C4030563|biopsy pancreas malignant neoplasm adenocarcinoma metaplastic apocrine
C4030563|biopsy of pancreas showed adenocarcinoma with apocrine metaplasia (procedure)
C4030453|biopsy of pancreas showed microinvasive squamous cell carcinoma
C4030453|biopsy of pancreas showed microinvasive squamous cell carcinoma (procedure)
C4030453|biopsy pancreas malig neoplasm carcinoma squamous cell microinvasive
C4030390|biopsy of pancreas showed vipoma
C4030390|biopsy of pancreas showed vipoma (procedure)
C4030390|biopsy pancreas malignant neoplasm carcinoma islet cell vipoma
C4030486|biopsy pancreas malignant neoplasm carcinoma large cell
C4030486|biopsy of pancreas showed large cell carcinoma (procedure)
C4030486|biopsy of pancreas showed large cell carcinoma
C4030499|biopsy of pancreas showed Hodgkin's sarcoma (procedure)
C4030499|biopsy pancreas malignant neoplasm lymphoma hodgkin's sarcoma
C4030499|biopsy of pancreas showed Hodgkin's sarcoma
C4030431|biopsy pancreas malignant neoplasm pancreatoblastoma
C4030431|biopsy of pancreas showed pancreatoblastoma
C4030431|biopsy of pancreas showed pancreatoblastoma (procedure)
C4030523|biopsy pancreas malignant neoplasm carcinoma epithelial-myoepithelial
C4030523|biopsy of pancreas showed epithelial-myoepithelial carcinoma
C4030523|biopsy of pancreas showed epithelial-myoepithelial carcinoma (procedure)
C4030402|biopsy pancreas malignant neoplasm sarcoma spindle cell
C4030402|biopsy of pancreas showed spindle cell sarcoma (procedure)
C4030402|biopsy of pancreas showed spindle cell sarcoma
C4030412|biopsy pancreas malignant neoplasm carcinoma small cell fusiform cell
C4030412|biopsy of pancreas showed small cell carcinoma, fusiform cell (procedure)
C4030412|biopsy of pancreas showed small cell carcinoma, fusiform cell
C4030507|biopsy of pancreas showed Hodgkin's granuloma
C4030507|biopsy pancreas malignant neoplasm lymphoma hodgkin's granuloma
C4030507|biopsy of pancreas showed Hodgkin's granuloma (procedure)
C4030467|biopsy of pancreas showed malignant lymphoplasmacytic lymphoma
C4030467|biopsy of pancreas showed malignant lymphoplasmacytic lymphoma (procedure)
C4030467|biopsy pancreas malignant neoplasm lymphoma lymphoplasmacytic
C4030405|biopsy pancreas malignant neoplasm carcinoma somatic
C4030405|biopsy of pancreas showed somatic carcinoma
C4030405|biopsy of pancreas showed somatic carcinoma (procedure)
C4030508|biopsy of pancreas showed histiocytic sarcoma
C4030508|biopsy of pancreas showed histiocytic sarcoma (procedure)
C4030508|biopsy pancreas malignant neoplasm sarcoma histiocytic
C4030468|biopsy of pancreas showed malignant lymphoma
C4030468|biopsy pancreas malignant neoplasm lymphoma
C4030468|biopsy of pancreas showed malignant lymphoma (procedure)
C4030414|biopsy of pancreas showed signet ring cell carcinoma
C4030414|biopsy pancreas malignant neoplasm carcinoma signet ring cell
C4030414|biopsy of pancreas showed signet ring cell carcinoma (procedure)
C4030509|biopsy pancreas malignant neoplasm adenocarcinoma hepatoid
C4030509|biopsy of pancreas showed hepatoid adenocarcinoma
C4030509|biopsy of pancreas showed hepatoid adenocarcinoma (procedure)
C4030570|biopsy pancreas malignant neoplasm adenocarcinoma in adenomatous polyp
C4030570|biopsy of pancreas showed adenocarcinoma in adenomatous polyp
C4030570|biopsy of pancreas showed adenocarcinoma in adenomatous polyp (procedure)
C4030524|biopsy of pancreas showed enterochromaffin cell carcinoid tumor (procedure)
C4030524|biopsy pancreas malig neoplasm carcinoid tumor enterochromaffin cell
C4030524|biopsy of pancreas showed enterochromaffin cell carcinoid tumor
C4030530|biopsy of pancreas showed composite carcinoid tumor
C4030530|biopsy pancreas malignant neoplasm carcinoid tumor composite
C4030530|biopsy of pancreas showed composite carcinoid tumor (procedure)
C4030534|biopsy pancreas malig carcinoma with osteoclast-like giant cells
C4030534|biopsy of pancreas showed carcinoma with osteoclast-like giant cells
C4030534|biopsy of pancreas showed carcinoma with osteoclast-like giant cells (procedure)
C4030514|biopsy of pancreas showed glassy cell carcinoma (procedure)
C4030514|biopsy pancreas malignant neoplasm carcinoma glassy cell
C4030514|biopsy of pancreas showed glassy cell carcinoma
C4030401|biopsy of pancreas showed spindle cell squamous cell carcinoma
C4030401|biopsy pancreas malig neoplasm carcinoma squamous cell spindle cell
C4030401|biopsy of pancreas showed spindle cell squamous cell carcinoma (procedure)
C4030418|biopsy pancreas malignant neoplasm carcinoma pseudosarcomatous
C4030418|biopsy of pancreas showed pseudosarcomatous carcinoma
C4030418|biopsy of pancreas showed pseudosarcomatous carcinoma (procedure)
C4030469|biopsy of pancreas showed malignant large B-cell diffuse lymphoma (procedure)
C4030469|biopsy pancreas malignant neoplasm lymphoma large b-cell diffuse
C4030469|biopsy of pancreas showed malignant large B-cell diffuse lymphoma
C4030518|biopsy of pancreas showed follicular lymphoma (procedure)
C4030518|biopsy pancreas malignant neoplasm lymphoma follicular
C4030518|biopsy of pancreas showed follicular lymphoma
C4030465|biopsy pancreas malignant neoplasm mastocytosis
C4030465|biopsy of pancreas showed malignant mastocytosis
C4030465|biopsy of pancreas showed malignant mastocytosis (procedure)
C4030555|biopsy pancreas malignant neoplasm carcinoma adenosquamous
C4030555|biopsy of pancreas showed adenosquamous carcinoma
C4030555|biopsy of pancreas showed adenosquamous carcinoma (procedure)
C4030393|biopsy pancreas malignant neoplasm sarcoma undifferentiated
C4030393|biopsy of pancreas showed undifferentiated sarcoma
C4030393|biopsy of pancreas showed undifferentiated sarcoma (procedure)
C4030449|biopsy of pancreas showed mucinous cystadenocarcinoma (procedure)
C4030449|biopsy pancreas malignant neoplasm cystadenocarcinoma mucinous
C4030449|biopsy of pancreas showed mucinous cystadenocarcinoma
C4030477|biopsy pancreas malig neoplasm carcinoma islet cell enteroglucagonoma
C4030477|biopsy of pancreas showed malignant enteroglucagonoma
C4030477|biopsy of pancreas showed malignant enteroglucagonoma (procedure)
C4030520|biopsy of pancreas showed extramedullary plasmacytoma
C4030520|biopsy pancreas malignant neoplasm plasmacytoma extramedullary
C4030520|biopsy of pancreas showed extramedullary plasmacytoma (procedure)
C4030413|biopsy of pancreas showed small cell carcinoma
C4030413|biopsy of pancreas showed small cell carcinoma (procedure)
C4030413|biopsy pancreas malignant neoplasm carcinoma small cell
C4030525|biopsy pancreas malignant neoplasm carcinosarcoma embryonal
C4030525|biopsy of pancreas showed embryonal carcinosarcoma (procedure)
C4030525|biopsy of pancreas showed embryonal carcinosarcoma
C4030457|biopsy of pancreas showed mast cell sarcoma
C4030457|biopsy pancreas malignant neoplasm sarcoma mast cell
C4030457|biopsy of pancreas showed mast cell sarcoma (procedure)
C4030519|biopsy pancreas malignant neoplasm sarcoma follicular dendritic cell
C4030519|biopsy of pancreas showed follicular dendritic cell sarcoma
C4030519|biopsy of pancreas showed follicular dendritic cell sarcoma (procedure)
C4030443|biopsy pancreas malignant neoplasm myosarcoma leiomyosarcoma myxoid
C4030443|biopsy of pancreas showed myxoid leiomyosarcoma (procedure)
C4030443|biopsy of pancreas showed myxoid leiomyosarcoma
C4030564|biopsy pancreas malignant neoplasm adenocarcinoma in villous adenoma
C4030564|biopsy of pancreas showed adenocarcinoma in villous adenoma
C4030564|biopsy of pancreas showed adenocarcinoma in villous adenoma (procedure)
C4030464|biopsy pancreas malignant neoplasm carcinosarcoma myoepithelioma
C4030464|biopsy of pancreas showed malignant myoepithelioma
C4030464|biopsy of pancreas showed malignant myoepithelioma (procedure)
C4030502|biopsy of pancreas showed Hodgkin's lymphoma with lymphocytic depletion with diffuse fibrosis
C4030502|biopsy pancreas malig lymphoma hodgkin's lymphocyt deplet diffuse fibrosis
C4030502|biopsy of pancreas showed Hodgkin's lymphoma with lymphocytic depletion with diffuse fibrosis (procedure)
C4030500|biopsy of pancreas showed Hodgkin's lymphoma with nodular sclerosis cellular phase (procedure)
C4030500|biopsy of pancreas showed Hodgkin's lymphoma with nodular sclerosis cellular phase
C4030500|biopsy pancreas malig lymphoma hodgkin's nodular sclerosis cellular phase
C4030408|biopsy of pancreas showed solid pseudopapillary carcinoma
C4030408|biopsy pancreas malignant neoplasm carcinoma solid pseudopapillary
C4030408|biopsy of pancreas showed solid pseudopapillary carcinoma (procedure)
C4030495|biopsy of pancreas showed intracystic carcinoma
C4030495|biopsy of pancreas showed intracystic carcinoma (procedure)
C4030495|biopsy pancreas malignant neoplasm carcinoma intracystic
C4030558|biopsy pancreas malig neoplasm adenocarcinoma metaplastic squamous
C4030558|biopsy of pancreas showed adenocarcinoma with squamous metaplasia (procedure)
C4030558|biopsy of pancreas showed adenocarcinoma with squamous metaplasia
C4030560|biopsy of pancreas showed adenocarcinoma with neuroendocrine differentiation
C4030560|biopsy pancreas malig adenocarc metaplastic neuroendocrine differentiation
C4030560|biopsy of pancreas showed adenocarcinoma with neuroendocrine differentiation (procedure)
C4030539|biopsy of pancreas showed carcinoma (procedure)
C4030539|biopsy of pancreas showed carcinoma
C4030539|biopsy pancreas malignant neoplasm carcinoma
C4030403|biopsy of pancreas showed spindle cell carcinoma (procedure)
C4030403|biopsy pancreas malignant neoplasm carcinoma spindle cell
C4030403|biopsy of pancreas showed spindle cell carcinoma
C4030517|biopsy of pancreas showed giant cell and spindle cell carcinoma
C4030517|biopsy of pancreas showed giant cell and spindle cell carcinoma (procedure)
C4030517|biopsy pancreas malig neoplasm carcinoma giant cell and spindle cell
C4030483|biopsy of pancreas showed large cell, nonkeratinizing squamous cell carcinoma
C4030483|biopsy of pancreas showed large cell, nonkeratinizing squamous cell carcinoma (procedure)
C4030483|biopsy pancreas malig carcinoma squamous cell large cell nonkeratinizing
C4030410|biopsy pancreas malig carcinoma squamous cell small cell nonkeratinizing
C4030410|biopsy of pancreas showed small cell, nonkeratinizing squamous cell carcinoma (procedure)
C4030410|biopsy of pancreas showed small cell, nonkeratinizing squamous cell carcinoma
C4030475|biopsy of pancreas showed malignant gastrinoma (procedure)
C4030475|biopsy of pancreas showed malignant gastrinoma
C4030475|biopsy pancreas malignant neoplasm carcinoma islet cell gastrinoma
C4030472|biopsy of pancreas showed malignant histiocytosis (procedure)
C4030472|biopsy of pancreas showed malignant histiocytosis
C4030472|biopsy pancreas malignant neoplasm lymphoma histiocytosis
C4030541|biopsy pancreas malignant neoplasm lymphoma burkitt's
C4030541|biopsy of pancreas showed Burkitt's lymphoma
C4030541|biopsy of pancreas showed Burkitt's lymphoma (procedure)
C4030421|biopsy of pancreas showed precursor B-cell lymphoblastic lymphoma
C4030421|biopsy pancreas malig lymphoma precursor cell lymphoblastic b-cell
C4030421|biopsy of pancreas showed precursor B-cell lymphoblastic lymphoma (procedure)
C4030444|biopsy pancreas malignant neoplasm myosarcoma
C4030444|biopsy of pancreas showed myosarcoma (procedure)
C4030444|biopsy of pancreas showed myosarcoma
C4030446|biopsy pancreas malignant neoplasm adenocarcinoma mucin-producing
C4030446|biopsy of pancreas showed mucin-producing adenocarcinoma
C4030446|biopsy of pancreas showed mucin-producing adenocarcinoma (procedure)
C4030526|biopsy of pancreas showed desmoplastic type duct carcinoma (procedure)
C4030526|biopsy of pancreas showed desmoplastic type duct carcinoma
C4030526|biopsy pancreas malignant neoplasm carcinoma duct, desmoplastic type
C4030429|biopsy pancreas malignant neoplasm carcinoma papillary
C4030429|biopsy of pancreas showed papillary carcinoma (procedure)
C4030429|biopsy of pancreas showed papillary carcinoma
C4030548|biopsy pancreas malignant neoplasm carcinoid tumor atypical
C4030548|biopsy of pancreas showed atypical carcinoid tumor
C4030548|biopsy of pancreas showed atypical carcinoid tumor (procedure)
C4030461|biopsy of pancreas showed malignant small cell type neoplasm
C4030461|biopsy pancreas malignant neoplasm small cell type
C4030461|biopsy of pancreas showed malignant small cell type neoplasm (procedure)
C4030394|biopsy pancreas malignant neoplasm carcinoma undifferentiated
C4030394|biopsy of pancreas showed undifferentiated carcinoma
C4030394|biopsy of pancreas showed undifferentiated carcinoma (procedure)
C4030485|biopsy of pancreas showed large cell carcinoma with rhabdoid phenotype
C4030485|biopsy of pancreas showed large cell carcinoma with rhabdoid phenotype (procedure)
C4030485|biopsy pancreas malig carcinoma large cell with rhabdoid phenotype
C4030529|biopsy of pancreas showed composite Hodgkin's and non-Hodgkin's lymphoma (procedure)
C4030529|biopsy of pancreas showed composite Hodgkin's and non-Hodgkin's lymphoma
C4030529|biopsy pancreas malig lymphoma composite hodgkin's & non-hodgkin's
C4030511|biopsy of pancreas showed grade 2 follicular lymphoma
C4030511|biopsy pancreas malignant neoplasm lymphoma follicular grade 2
C4030511|biopsy of pancreas showed grade 2 follicular lymphoma (procedure)
C4030420|biopsy of pancreas showed precursor cell lymphoblastic lymphoma
C4030420|biopsy of pancreas showed precursor cell lymphoblastic lymphoma (procedure)
C4030420|biopsy pancreas malignant neoplasm lymphoma precursor cell lymphoblastic
C4030424|biopsy of pancreas showed plasmacytoma (procedure)
C4030424|biopsy pancreas malignant neoplasm plasmacytoma
C4030424|biopsy of pancreas showed plasmacytoma
C4030574|biopsy of pancreas showed acinar cell carcinoma
C4030574|biopsy of pancreas showed acinar cell carcinoma (procedure)
C4030574|biopsy pancreas malignant neoplasm carcinoma acinar cell
C4030430|biopsy of pancreas showed papillary adenocarcinoma (procedure)
C4030430|biopsy pancreas malignant neoplasm adenocarcinoma papillary
C4030430|biopsy of pancreas showed papillary adenocarcinoma
C4030478|biopsy of pancreas showed malignant enterochromaffin-like cell carcinoid tumor
C4030478|biopsy pancreas malig carcinoid tumor enterochromaffin-like cell
C4030478|biopsy of pancreas showed malignant enterochromaffin-like cell carcinoid tumor (procedure)
C4030459|biopsy of pancreas showed malignant spindle cell type neoplasm (procedure)
C4030459|biopsy pancreas malignant neoplasm spindle cell type
C4030459|biopsy of pancreas showed malignant spindle cell type neoplasm
C4030423|biopsy of pancreas showed pleomorphic carcinoma (procedure)
C4030423|biopsy pancreas malignant neoplasm carcinoma pleomorphic
C4030423|biopsy of pancreas showed pleomorphic carcinoma
C4030528|biopsy of pancreas showed cystadenocarcinoma
C4030528|biopsy pancreas malignant neoplasm carcinoma cystadenocarcinoma
C4030528|biopsy of pancreas showed cystadenocarcinoma (procedure)
C4030496|biopsy of pancreas showed interdigitating dendritic cell sarcoma
C4030496|biopsy pancreas malig neoplasm sarcoma interdigitating dendritic cell
C4030496|biopsy of pancreas showed interdigitating dendritic cell sarcoma (procedure)
C4030439|biopsy of pancreas showed non-Hodgkin's lymphoma
C4030439|biopsy of pancreas showed non-Hodgkin's lymphoma (procedure)
C4030439|biopsy pancreas malignant neoplasm lymphoma non-hodgkin's
C4030503|biopsy of pancreas showed Hodgkin's lymphoma with lymphocytic depletion
C4030503|biopsy of pancreas showed Hodgkin's lymphoma with lymphocytic depletion (procedure)
C4030503|biopsy pancreas malig lymphoma hodgkin's lymphocytic depletion
C4030531|biopsy of pancreas showed comedocarcinoma (procedure)
C4030531|biopsy pancreas malignant neoplasm carcinoma comedocarcinoma
C4030531|biopsy of pancreas showed comedocarcinoma
C4030427|biopsy of pancreas showed papillary cystadenocarcinoma (procedure)
C4030427|biopsy pancreas malignant neoplasm cystadenocarcinoma papillary
C4030427|biopsy of pancreas showed papillary cystadenocarcinoma
C4030559|biopsy of pancreas showed adenocarcinoma with spindle cell metaplasia (procedure)
C4030559|biopsy of pancreas showed adenocarcinoma with spindle cell metaplasia
C4030559|biopsy pancreas malig neoplasm adenocarcinoma metaplastic spindle cell
C4030572|biopsy pancreas malignant neoplasm carcinoid tumor adenocarcinoid
C4030572|biopsy of pancreas showed adenocarcinoid tumor (procedure)
C4030572|biopsy of pancreas showed adenocarcinoid tumor
C4030466|biopsy of pancreas showed malignant mantle cell lymphoma
C4030466|biopsy of pancreas showed malignant mantle cell lymphoma (procedure)
C4030466|biopsy pancreas malignant neoplasm lymphoma mantle cell
C4030471|biopsy of pancreas showed malignant immunoblastic large B-cell diffuse lymphoma
C4030471|biopsy pancreas malig lymphoma large b-cell diffuse immunoblastic
C4030471|biopsy of pancreas showed malignant immunoblastic large B-cell diffuse lymphoma (procedure)
C4030522|biopsy of pancreas showed epithelioid leiomyosarcoma
C4030522|biopsy of pancreas showed epithelioid leiomyosarcoma (procedure)
C4030522|biopsy pancreas malig neoplasm myosarcoma leiomyosarcoma epithelioid
C4030454|biopsy of pancreas showed medullary carcinoma (procedure)
C4030454|biopsy of pancreas showed medullary carcinoma
C4030454|biopsy pancreas malignant neoplasm carcinoma medullary
C4030547|biopsy of pancreas showed basal cell adenocarcinoma (procedure)
C4030547|biopsy pancreas malignant neoplasm adenocarcinoma basal cell
C4030547|biopsy of pancreas showed basal cell adenocarcinoma
C4030451|biopsy pancreas malig mixed islet cell & exocrine adenocarcinoma
C4030451|biopsy of pancreas showed mixed islet cell and exocrine adenocarcinoma (procedure)
C4030451|biopsy of pancreas showed mixed islet cell and exocrine adenocarcinoma
C4030476|biopsy of pancreas showed malignant epithelioma (procedure)
C4030476|biopsy pancreas malignant neoplasm carcinoma epithelioma
C4030476|biopsy of pancreas showed malignant epithelioma
C4030462|biopsy of pancreas showed malignant small B-cell lymphocytic lymphoma (procedure)
C4030462|biopsy pancreas malignant neoplasm lymphoma small b-cell lymphocytic
C4030462|biopsy of pancreas showed malignant small B-cell lymphocytic lymphoma
C4030501|biopsy pancreas malignant neoplasm lymphoma hodgkin's nodular sclerosis
C4030501|biopsy of pancreas showed Hodgkin's lymphoma with nodular sclerosis (procedure)
C4030501|biopsy of pancreas showed Hodgkin's lymphoma with nodular sclerosis
C4030493|biopsy pancreas malig adenocarcinoma intraductal papillary w/ invasion
C4030493|biopsy of pancreas showed intraductal papillary adenocarcinoma with invasion (procedure)
C4030493|biopsy of pancreas showed intraductal papillary adenocarcinoma with invasion
C4030463|biopsy of pancreas showed malignant neoplasm
C4030463|biopsy pancreas malignant neoplasm
C4030463|biopsy of pancreas showed malignant neoplasm (procedure)
C4030490|biopsy pancreas malig carcinoma intraductal papillary-mucinous invasive
C4030490|biopsy of pancreas showed invasive intraductal papillary-mucinous carcinoma
C4030490|biopsy of pancreas showed invasive intraductal papillary-mucinous carcinoma (procedure)
C4030395|biopsy of pancreas showed tubular adenocarcinoma
C4030395|biopsy pancreas malignant neoplasm adenocarcinoma tubular
C4030395|biopsy of pancreas showed tubular adenocarcinoma (procedure)
C4030515|biopsy of pancreas showed giant cell sarcoma (procedure)
C4030515|biopsy of pancreas showed giant cell sarcoma
C4030515|biopsy pancreas malignant neoplasm sarcoma giant cell
C4030474|biopsy pancreas malignant neoplasm giant cell type
C4030474|biopsy of pancreas showed malignant giant cell type neoplasm (procedure)
C4030474|biopsy of pancreas showed malignant giant cell type neoplasm
C4030554|biopsy of pancreas showed anaplastic carcinoma (procedure)
C4030554|biopsy of pancreas showed anaplastic carcinoma
C4030554|biopsy pancreas malignant neoplasm carcinoma anaplastic
C4030397|biopsy pancreas malig carcinoma squamous cell with horn formation
C4030397|biopsy of pancreas showed squamous cell carcinoma with horn formation
C4030397|biopsy of pancreas showed squamous cell carcinoma with horn formation (procedure)
C4030535|biopsy pancreas malignant neoplasm carcinoma simplex
C4030535|biopsy of pancreas showed carcinoma simplex (procedure)
C4030535|biopsy of pancreas showed carcinoma simplex
C4030445|biopsy of pancreas showed mucoepidermoid carcinoma (procedure)
C4030445|biopsy pancreas malignant neoplasm carcinoma mucoepidermoid
C4030445|biopsy of pancreas showed mucoepidermoid carcinoma
C4030512|biopsy of pancreas showed grade 1 follicular lymphoma
C4030512|biopsy of pancreas showed grade 1 follicular lymphoma (procedure)
C4030512|biopsy pancreas malignant neoplasm lymphoma follicular grade 1
C4030550|biopsy pancreas malig neoplasm lymphoma mature t-cell angioimmunoblastic
C4030550|biopsy of pancreas showed angioimmunoblastic T-cell lymphoma (procedure)
C4030550|biopsy of pancreas showed angioimmunoblastic T-cell lymphoma
C4030549|biopsy of pancreas showed angiomyosarcoma (procedure)
C4030549|biopsy pancreas malignant neoplasm myosarcoma angiomyosarcoma
C4030549|biopsy of pancreas showed angiomyosarcoma
C4030540|biopsy of pancreas showed carcinoid tumor (procedure)
C4030540|biopsy pancreas malignant neoplasm carcinoid tumor
C4030540|biopsy of pancreas showed carcinoid tumor
C1409082|pancreas; islet cell adenocarcinoma with exocrine
C1386256|adenocarcinoma; islet cell with exocrine, unspecified site
C1391905|carcinoma; islet cell, met exocrine, unspecified site
C1396226|islet cell; adenocarcinoma, met exocrine, unspecified site
C1396227|islet cell; carcinoma with exocrine, unspecified site
C0279884|cellular diagnosis, pancreatic cancer
C0279884|pancreas cancer cellular diagnosis
C0279884|pancreatic cancer cellular diagnosis
C0280222|stage, pancreatic cancer
C0280222|pancreatic cancer stage
C1335307|malignant lymphoma of pancreatic lymph nodes (diagnosis)
C1335307|malignant lymphoma of pancreatic lymph nodes
C1335307|pancreatic lymphoma
C1335307|Lymphoma of Pancreas
C1335307|Lymphoma of the Pancreas
C1276580|T2: Tumor limited to pancreas and > 2 cm in greatest dimension (finding)
C1276580|T2: Tumor limited to pancreas and > 2 cm in greatest dimension
C1276580|T2: Tumour limited to pancreas and > 2 cm in greatest dimension
C1276580|T2: Tumor limited to pancreas and > 2 cm in greatest dimension (tumor staging)
C0341485|malignant cystic neoplasm of exocrine pancreas
C0341485|pancreatic neoplasm malignant exocrine cystic
C0341485|malignant cystic neoplasm of exocrine pancreas (diagnosis)
C0341485|Malignant cystic tumor of exocrine pancreas
C0341485|Malignant cystic tumour of exocrine pancreas
C0341485|Malignant cystic tumor of exocrine pancreas (disorder)
C0238337|cystadenocarcinoma of pancreas (diagnosis)
C0238337|cystadenocarcinoma of pancreas
C0238337|Cystadenocarcinoma - pancreas
C0238337|Cystadenocarcinoma of the pancreas
C0238337|Cystadenocarcinoma pancreas
C0238337|Cystadenocarcinoma of pancreas (disorder)
C0238337|Pancreatic Cystadenocarcinoma
C0345933|Pancreatic Carcinoid Tumor
C0345933|Carcinoid Neoplasm of Pancreas
C0345933|Carcinoid Neoplasm of the Pancreas
C0345933|Carcinoid Tumor of Pancreas
C0345933|Carcinoid Tumor of the Pancreas
C0345933|Pancreatic Serotonin Producing Neoplasm
C0345933|EC Cell, Serotonin Producing Pancreatic NET
C0345933|Pancreatic Serotonin Producing Tumor
C0345933|Enterochromaffin Cell Serotonin-Producing Pancreatic Neuroendocrine Tumor
C0345933|EC Cell, Serotonin Producing Pancreatic Neuroendocrine Tumor
C0345933|Carcinoid tumour of the pancreas
C0345933|Carcinoid tumour of pancreas
C0345933|Carcinoid tumor of pancreas (disorder)
C0345933|Serotonin-Producing Tumor of Pancreas
C0345933|Serotonin-Producing Tumor of the Pancreas
C2033026|lymphocyte-rich Hodgkin's lymphoma of pancreas (diagnosis)
C2033026|lymphocyte-rich Hodgkin's lymphoma of pancreas
C2033030|nodular sclerosing Hodgkin's lymphoma of pancreas (diagnosis)
C2033030|nodular sclerosing Hodgkin's lymphoma of pancreas
C2033048|grade 3 follicular lymphoma of pancreas (diagnosis)
C2033048|grade 3 follicular lymphoma of pancreas
C2033055|mature T-cell lymphoma of pancreas (diagnosis)
C2033055|mature T-cell lymphoma of pancreas
C2046512|pancreatic malignant lymphoma Hodgkin's and non-Hodgkin's
C2046512|composite Hodgkin's and non-Hodgkin's lymphoma of pancreas (diagnosis)
C2046512|composite Hodgkin's and non-Hodgkin's lymphoma of pancreas
C2033052|lymphoplasmacytic lymphoma of pancreas
C2033052|lymphoplasmacytic lymphoma of pancreas (diagnosis)
C2033045|follicular lymphoma of pancreas
C2033045|follicular lymphoma of pancreas (diagnosis)
C2033046|grade 1 follicular lymphoma of pancreas (diagnosis)
C2033046|grade 1 follicular lymphoma of pancreas
C2046585|Hodgkin's granuloma of pancreas
C2046585|Hodgkin's granuloma of pancreas (diagnosis)
C2033058|small B-cell lymphocytic lymphoma of pancreas
C2033058|small B-cell lymphocytic lymphoma of pancreas (diagnosis)
C2033053|mantle cell lymphoma of pancreas
C2033053|mantle cell lymphoma of pancreas (diagnosis)
C2033051|immunoblastic large B-cell diffuse lymphoma of pancreas (diagnosis)
C2033051|immunoblastic large B-cell diffuse lymphoma of pancreas
C2113717|precursor cell lymphoblastic lymphoma of pancreas (diagnosis)
C2113717|precursor cell lymphoblastic lymphoma of pancreas
C2205509|mast cell sarcoma of pancreas
C2205509|mast cell sarcoma of pancreas (diagnosis)
C2033050|large B-cell diffuse lymphoma of pancreas (diagnosis)
C2033050|large B-cell diffuse lymphoma of pancreas
C2033047|grade 2 follicular lymphoma of pancreas
C2033047|grade 2 follicular lymphoma of pancreas (diagnosis)
C2113646|precursor B-cell lymphoblastic lymphoma of pancreas (diagnosis)
C2113646|precursor B-cell lymphoblastic lymphoma of pancreas
C2113786|precursor T-cell lymphoblastic lymphoma of pancreas
C2113786|precursor T-cell lymphoblastic lymphoma of pancreas (diagnosis)
C2033029|mixed cellularity Hodgkin's lymphoma of pancreas
C2033029|mixed cellularity Hodgkin's lymphoma of pancreas (diagnosis)
C2033033|grade 2 nodular sclerosing Hodgkin's lymphoma of pancreas (diagnosis)
C2033033|grade 2 nodular sclerosing Hodgkin's lymphoma of pancreas
C2033054|marginal zone B-cell lymphoma of pancreas (diagnosis)
C2033054|marginal zone B-cell lymphoma of pancreas
C2033056|angioimmunoblastic T-cell lymphoma of pancreas
C2033056|angioimmunoblastic T-cell lymphoma of pancreas (diagnosis)
C2033056|angioimmunoblastic lymphadenopathy with dysproteinemia (AILD) of pancreas
C2033032|grade 1 nodular sclerosing Hodgkin's lymphoma of pancreas
C2033032|grade 1 nodular sclerosing Hodgkin's lymphoma of pancreas (diagnosis)
C2033057|NK/T-cell lymphoma of pancreas (diagnosis)
C2033057|NK/T-cell lymphoma of pancreas
C2033027|Hodgkin's disease, lymphocytic depletion of pancreas (diagnosis)
C2033027|Hodgkin's disease, lymphocytic depletion of pancreas
C2033028|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of pancreas
C2033028|Hodgkin's disease, lymphocytic depletion, diffuse fibrosis of pancreas (diagnosis)
C2033031|nodular sclerosing Hodgkin's lymphoma in cellular phase of pancreas
C2033031|nodular sclerosing Hodgkin's lymphoma in cellular phase of pancreas (diagnosis)
C2046725|Hodgkin's sarcoma of pancreas (diagnosis)
C2046725|Hodgkin's sarcoma of pancreas
C2033049|malignant histiocytosis of pancreas
C2033049|malignant histiocytosis of pancreas (diagnosis)
C2205522|Sezary syndrome of pancreas (diagnosis)
C2205522|Sezary syndrome of pancreas
C0153620|Urethra
C0153620|Malignant neoplasm of urethra
C0153620|malignant neoplasm of urethra (diagnosis)
C0153620|malignant tumor of urethra
C0153620|Malign neopl urethra
C0153620|Malignant tumour of urethra
C0153620|Malignant tumour of urethra (disorder)
C0153620|Malignant urethral tumor
C0153620|Malignant urethral tumour
C0153620|Malignant tumor of urethra (disorder)
C0153620|Malignant Neoplasm of the Urethra
C0153620|Malignant Tumor of the Urethra
C0153620|Malignant Urethra Neoplasm
C0153620|Malignant Urethra Tumor
C0153620|Malignant Urethral Neoplasm
C0153620|Neoplasm malig;urethra
C0153620|malignant neosplasm of the urethra
C0153621|Malignant neoplasm of paraurethral glands
C0153621|Paraurethral gland
C0153621|Malignant neoplasm of paraurethral gland
C0153621|malignant neoplasm of paraurethral gland (diagnosis)
C0153621|malignant tumor of paraurethral gland
C0153621|Mal neo paraurethral
C0153621|Malignant tumour of paraurethral gland
C0153621|Malignant tumor of paraurethral gland (disorder)
C0349055|Malignant neoplasm overlapping urinary organ site
C0349055|Overlapping lesion of urinary organs
C0349055|Malignant neoplasm of overlapping sites of urinary organs
C0349055|malignant neoplasm of urinary organs overlapping sites
C0349055|malignant neoplasm of overlapping sites of urinary organs (diagnosis)
C0349055|Malignant neoplasm of overlapping lesion of urinary organs
C0349055|Malignant neoplasm of overlapping lesion of urinary organs (disorder)
C0348371|Malignant neoplasm of urinary organ, unspecified
C0348371|Urinary organ, unspecified
C0348371|Mal neo urinary NOS
C0348371|Cancer of urinary organs
C0348371|Malignant neoplasm of urinary organ (disorder)
C0348371|Cancer of urinary organ
C0348371|Malignant neoplasm of urinary organ
C0348371|[X]Malignant neoplasm of urinary organ, unspecified
C0348371|[X]Malignant neoplasm of urinary organ, unspecified (disorder)
C0348371|Urinary organs--Cancer
C0348371|Malignant neoplasm of urinary organ, site unspecified
C0346890|Malignant neoplasm of other and unspecified urinary organs
C0346890|Cancer of other urinary organs
C0346890|Malignant neoplasm of other urinary organs (disorder)
C0346890|Malignant neoplasm of other urinary organs
C0700101|Urethral Carcinoma
C0700101|carcinoma of urethra (diagnosis)
C0700101|urethral carcinoma (diagnosis)
C0700101|carcinoma of urethra
C0700101|Cancers, Urethra
C0700101|Urethra Cancers
C0700101|Cancer, Urethral
C0700101|Cancers, Urethral
C0700101|Urethral Cancers
C0700101|Carcinoma;urethra
C0700101|Cancer, Urethra
C0700101|urethral cancer
C0700101|Urethra cancer
C0700101|Urethral cancer NOS
C0700101|Cancer of the Urethra
C0700101|CA - Cancer of urethra
C0700101|Urethral Ca
C0700101|Urethra Carcinoma
C0700101|Carcinoma of the Urethra
C0700101|Cancer of Urethra
C0153619|Malignant neoplasm of ureter
C0153619|URETER, CANCER OF
C0153619|malignant neoplasm of ureter (diagnosis)
C0153619|Ureter Cancers
C0153619|Cancer, Ureteral
C0153619|Cancers, Ureteral
C0153619|Ureteral Cancers
C0153619|malignant tumor of ureter
C0153619|ureteral cancer
C0153619|Malign neopl ureter
C0153619|Malignant tumour of ureter (disorder)
C0153619|Malignant tumour of ureter
C0153619|Ureters--Cancer
C0153619|Ureter cancer
C0153619|Ureteric cancer
C0153619|Ureteric cancer NOS
C0153619|Cancer of the Ureter
C0153619|Ureter Ca
C0153619|Cancer of ureter
C0153619|Malignant tumor of ureter (disorder)
C0153619|Malignant Neoplasm of the Ureter
C0153619|Malignant Tumor of the Ureter
C0153619|Malignant Ureter Neoplasm
C0153619|Malignant Ureter Tumor
C0153619|Malignant Ureteral Neoplasm
C0153619|Malignant Ureteral Tumor
C0153619|Neoplasm malig;ureter
C0153619|malignant neosplasm of the ureter
C0153618|Malignant neoplasm of renal pelvis
C0153618|malignant neoplasm of renal pelvis (diagnosis)
C0153618|malignant tumor of renal pelvis
C0153618|Malig neo renal pelvis
C0153618|Malignant neoplasm of renal pelvis NOS
C0153618|Malignant neoplasm of renal pelvis NOS (disorder)
C0153618|Renal pelvis cancer NOS
C0153618|Malignant tumour of renal pelvis
C0153618|Malignant tumor of renal pelvis (disorder)
C0153618|Malignant Neoplasm of the Renal Pelvis
C0153618|Malignant Renal Pelvis Neoplasm
C0153618|Malignant Renal Pelvis Tumor
C0153618|Malignant Tumor of the Renal Pelvis
C0153622|Malignant neoplasm of other specified sites of urinary organs
C0153622|Mal neo urinary NEC
C0494158|Malignant neoplasm of kidney, except renal pelvis
C0494158|Malig neopl kidney
C0494158|Malignant neoplasm of kidney, except pelvis
C0494158|Malignant neoplasm of kidney, excl pelvis
C0494158|Malignant neoplasm of kidney, excluding pelvis
C0494158|Malignant Neoplasm of Kidney Except Pelvis
C0494158|Malignant Kidney Neoplasm Except Pelvis
C0600079|carcinoma of ureter
C0600079|carcinoma of ureter (diagnosis)
C0600079|Ureter Carcinoma
C0600079|Carcinoma;ureter
C0600079|Ureteral Carcinoma
C0600079|Carcinoma of the Ureter
C0751571|Malignant Urinary System Neoplasm
C0751571|Malignant Urinary Tract Neoplasm
C0751571|Malignant neoplasm of urinary system
C0751571|malignant neoplasm of urinary organs (diagnosis)
C0751571|malignant neoplasm of urinary organs
C0751571|Malignant neoplasms of urinary tract
C0751571|Malignant tumor of urinary tract proper (disorder)
C0751571|Malignant tumor of urinary tract
C0751571|Malignant tumour of urinary tract
C0751571|Malignant tumor of urinary tract proper
C0751571|Malignant tumor of urinary tract (disorder)
C0751571|Malignant tumour of urinary tract proper
C0751571|Cancers, Urinary Tract
C0751571|Urinary Tract Cancers
C0751571|Cancer, Urologic
C0751571|Cancers, Urologic
C0751571|Urologic Cancers
C0751571|Cancer, Urological
C0751571|Cancers, Urological
C0751571|Urological Cancers
C0751571|Malignant neoplasm of urinary system NOS
C0751571|Cancer, Urinary Tract
C0751571|Malignant neoplasms of urinary tract (C64-C68)
C0751571|[X]Malignant neoplasm of urinary tract (disorder)
C0751571|[X]Malignant neoplasm of urinary tract
C0751571|malignant neoplasm of urinary tract proper (diagnosis)
C0751571|malignant neoplasm of urinary tract proper
C0751571|malignant neoplasm urinary system
C0751571|urinary neoplasm malignant of tract proper
C0751571|malignant neoplasm of urinary system (diagnosis)
C0751571|Urothelial/bladder cancer, NOS
C0751571|Urothelial tract/bladder cancer, NOS
C0751571|Malignant urinary tract neoplasm NOS
C0751571|Cancer of the Urinary Tract
C0751571|Urological Cancer
C0751571|Urologic Cancer
C0751571|Urinary Tract Cancer
C0751571|Malignant neoplasm of urinary system, NOS
C0751571|Cancer of Urinary Tract
C0751571|Neoplasm malig;urological
C0751571|malignant neosplasm of the urological system
C1276598|Ta: Noninvasive papillary carcinoma (urinary tract) (finding)
C1276598|Ta: Noninvasive papillary carcinoma (urinary tract)
C1276598|Ta: Noninvasive papillary carcinoma (urinary tract) (tumor staging)
C0023418|Leukemias
C0023418|Leukemia
C0023418|Leukemia of unspecified cell type
C0023418|Leukaemia
C0023418|Leukaemia of unspecified cell type
C0023418|Leukaemia, unspecified
C0023418|Leukemia, unspecified
C0023418|Leukemia, disease
C0023418|Leukaemia, disease
C0023418|leukemia (diagnosis)
C0023418|Leukaemia, no ICD-O subtype
C0023418|Leukemia, no ICD-O subtype
C0023418|Leukaemias
C0023418|Leukemia NOS
C0023418|Leukemia [Disease/Finding]
C0023418|Leucocythaemias
C0023418|Leucocythemias
C0023418|Leucocythaemia
C0023418|Leucocythemia
C0023418|Leukaemia of unspecified cell type (disorder)
C0023418|[M]Leukemia NOS
C0023418|Leukemia (disorder)
C0023418|[M]Leukaemia NOS
C0023418|Leukemia of unspecified cell type (disorder)
C0023418|[M]Leukemia unspecified, NOS
C0023418|[M]leukemia unspecified, NOS (morphologic abnormality)
C0023418|[M]Leukaemia NOS (disorder)
C0023418|Leukemia NOS (disorder)
C0023418|[M]leukemia NOS (morphologic abnormality)
C0023418|[M]Leukaemia unspecified, NOS
C0023418|Leukaemia NOS
C0023418|[M]Leukaemias unspecified
C0023418|[M]leukemias unspecified (morphologic abnormality)
C0023418|[M]Leukemias unspecified
C0023418|Leukemia, no ICD-O subtype (morphologic abnormality)
C0023418|Leukemia, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0023418|Leukemia, no International Classification of Diseases for Oncology subtype
C0023418|Leukemia, NOS
C0023418|LEUKEMIA, MALIGNANT
C0023418|-- Leukemia
C0023418|Blood (Leukemia)
C0023418|Leukemias, General
C0023418|Leukemia unspecified
C0023418|Unspecified leukemia without mention of remission
C0023418|Unspecified leukaemia without mention of remission
C0023418|Leukaemia unspecified
C0023418|Unspecified leukaemia
C0023418|Unspecified leukemia
C0023418|Leukaemia morphology
C0023418|Leukemia morphology
C0023418|Chronic leukaemia [obs]
C0023418|Chronic leukemia [obs]
C0023418|Leukemia, disease (disorder)
C0023418|Aleukaemic leukaemia [obs]
C0023418|Aleukemic leukemia [obs]
C0023418|Subacute leukaemia [obs]
C0023418|Subacute leukemia [obs]
C0023418|Leukaemia, NOS
C0023418|Leukaemia, NOS, without mention of remission
C0023418|Leukemia, NOS, without mention of remission
C0023418|Leukemia, morphology (morphologic abnormality)
C0026764|Multiple Myeloma
C0026764|Multiple Myelomas
C0026764|Myeloma, Plasma Cell
C0026764|Myelomas, Multiple
C0026764|plasma cell myeloma
C0026764|myelomatosis
C0026764|Myelomas, Plasma-Cell
C0026764|Plasma-Cell Myeloma
C0026764|Plasma-Cell Myelomas
C0026764|Multiple myeloma / Plasma cell neoplasm
C0026764|MYELOMA, MULTIPLE
C0026764|myeloma
C0026764|multiple myeloma (diagnosis)
C0026764|Multiple myeloma, no ICD-O subtype
C0026764|Cell Myeloma, Plasma
C0026764|Cell Myelomas, Plasma
C0026764|Plasma Cell Myelomas
C0026764|Myelomas, Plasma Cell
C0026764|Kahler's disease
C0026764|Multiple myeloma NOS
C0026764|Multiple Myeloma [Disease/Finding]
C0026764|Myeloma, Plasma-Cell
C0026764|Myelomatoses
C0026764|Disease, Kahler
C0026764|Myeloma-Multiples
C0026764|Myeloma Multiple
C0026764|Myeloma;multiple
C0026764|Myeloma-Multiple
C0026764|Kahler Disease
C0026764|Multiple myeloma myelomatosis
C0026764|Myeloma (disorder)
C0026764|Multiple myeloma (disorder)
C0026764|Multiple myeloma, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0026764|Multiple myeloma, no ICD-O subtype (morphologic abnormality)
C0026764|Multiple myeloma, no International Classification of Diseases for Oncology subtype
C0026764|MYELOMA, PLASMA CELL, MALIGNANT
C0026764|Myeloma, NOS
C0026764|[M]Plasma cell myeloma
C0026764|Peripheral plasma cell myeloma
C0026764|Myelomatosis multiple
C0026764|Plasmacytic myeloma
C0026764|plasma cell neoplasm
C0026764|neoplasm, plasma cell
C0026764|multiple myeloma and other plasma cell neoplasms
C0026764|plasma cell neoplasms
C0026764|Kahler
C0026764|myelomata; multiple
C0026764|Multiple myeloma (clinical)
C0026764|Multiple myeloma, morphology (morphologic abnormality)
C0019829|Disease, Hodgkin
C0019829|Hodgkin Disease
C0019829|Hodgkin's Disease
C0019829|Lymphogranulomas, Malignant
C0019829|Malignant Lymphogranuloma
C0019829|Malignant Lymphogranulomas
C0019829|Disease, Hodgkin's
C0019829|Disease, Hodgkins
C0019829|Hodgkin's disease, unspecified
C0019829|Hodgkin lymphoma
C0019829|HODGKIN DIS
C0019829|HODGKINS DIS
C0019829|Hodgkin's Lymphoma
C0019829|Lymphoma, Hodgkin's
C0019829|Lymphoma, Hodgkin
C0019829|Hodgkins Lymphoma
C0019829|Hodgkin's granuloma
C0019829|Hodgkin's sarcoma
C0019829|lymphogranulomatosis (malignant)
C0019829|Hodgkin's paragranuloma, NOS
C0019829|Hodgkin's disease, NOS
C0019829|Hodgkin lymphoma, no ICD-O subtype
C0019829|Hodgkin's paragranuloma -RETIRED-
C0019829|Lymphomas Hodgkin's disease
C0019829|Hodgins
C0019829|Hodgkin sarcoma
C0019829|Hodgkin granuloma
C0019829|Hodgkin lymphoma, unspecified
C0019829|Hodgkin Disease [Disease/Finding]
C0019829|Granuloma, Hodgkins
C0019829|Granuloma, Hodgkin
C0019829|Hodgkins Disease
C0019829|Lymphogranuloma, Malignant
C0019829|Granuloma, Hodgkin's
C0019829|Granuloma, Malignant
C0019829|Disease;Hodgkins
C0019829|Lymphoma;Hodgkins
C0019829|Sarcoma;Hodgkins
C0019829|Hodgkins Granuloma
C0019829|Malignant Granulomas
C0019829|Malignant Granuloma
C0019829|lymphogranulomatosis
C0019829|Hodgkin's paragranuloma (morphologic abnormality)
C0019829|[M]Hodgkin's disease NOS
C0019829|Hodgkin's disease NOS
C0019829|Hodgkin's sarcoma of unspecified site
C0019829|Hodgkin's paragranuloma of unspecified site
C0019829|Hodgkin's sarcoma NOS
C0019829|Hodgkin's granuloma NOS (disorder)
C0019829|[M]Hodgkin's paragranuloma (morphologic abnormality)
C0019829|[M]Hodgkin's disease NOS (morphologic abnormality)
C0019829|[M]Hodgkin's paragranuloma
C0019829|[M]Lymphogranuloma, malignant (morphologic abnormality)
C0019829|Hodgkin's paragranuloma (disorder)
C0019829|[M]Hodgkin's disease NOS (& [lymphogranuloma malignant])
C0019829|Hodgkin's disease NOS, unspecified site (disorder)
C0019829|Hodgkin's paragranuloma NOS (disorder)
C0019829|Hodgkin's granuloma of unspecified site
C0019829|Hodgkin's sarcoma NOS (disorder)
C0019829|Hodgkin's disease NOS, unspecified site
C0019829|Hodgkin's disease NOS (disorder)
C0019829|Hodgkin's paragranuloma
C0019829|[M]Lymphogranuloma, malignant
C0019829|Hodgkin's paragranuloma of unspecified site (disorder)
C0019829|[M]Hodgkin's disease NOS (& [lymphogranuloma malignant]) (disorder)
C0019829|Hodgkin's paragranuloma NOS
C0019829|Hodgkin's granuloma NOS
C0019829|Hodgkin's sarcoma of unspecified site (disorder)
C0019829|[M]Hodgkin's disease NOS (disorder)
C0019829|Hodgkin's disease (disorder)
C0019829|Hodgkin's granuloma of unspecified site (disorder)
C0019829|Hodgkin lymphoma, no ICD-O subtype (morphologic abnormality)
C0019829|Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype
C0019829|Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0019829|Hodgkin lymphoma, NOS
C0019829|Hodgkin disease (diagnosis)
C0019829|Hodgkin disease sarcoma (diagnosis)
C0019829|Hodgkin disease sarcoma
C0019829|Hodgkin disease granuloma
C0019829|Hodgkin disease granuloma (diagnosis)
C0019829|Hodgkin disease paragranuloma
C0019829|Hodgkin disease paragranuloma (diagnosis)
C0019829|[M]Hodgkin's disease
C0019829|[M]Hodgkin's granuloma
C0019829|[M]Hodgkin's sarcoma
C0019829|CHL
C0019829|LYMPHOMA, HODGKIN, CLASSIC
C0019829|Lymphoma, Hodgkins
C0019829|Hodgkin's disease, unspecified type
C0019829|Hodgkin`s disease
C0019829|Malignant Hodgkin's lymphoma
C0019829|Malignant lymphoma, Hodgkin's
C0019829|HD - Hodgkin's disease
C0019829|Hodgkin granuloma [obs] (morphologic abnormality)
C0019829|Hodgkin granuloma [obs]
C0019829|Hodgkin paragranuloma [obs]
C0019829|Hodgkin paragranuloma, nodular [obs]
C0019829|Hodgkin sarcoma [obs] (morphologic abnormality)
C0019829|Hodgkin sarcoma [obs]
C0019829|Hodgkin's disease (clinical)
C0019829|Hodgkin's granuloma (clinical)
C0019829|Hodgkin's granuloma (disorder)
C0019829|Hodgkin's paragranuloma (clinical)
C0019829|Hodgkin's sarcoma (clinical)
C0019829|Hodgkin's sarcoma (disorder)
C0019829|Hodgkin; granuloma
C0019829|Hodgkin; lymphoma
C0019829|Hodgkin; paragranuloma
C0019829|Hodgkin; sarcoma
C0019829|Hodgkin
C0019829|disease; Hodgkin
C0019829|granuloma; Hodgkin
C0019829|granuloma; malignant
C0019829|lymphoma; Hodgkin
C0019829|malignant; granuloma
C0019829|paragranuloma; Hodgkin
C0019829|sarcoma; Hodgkin
C0019829|Hodgkin's paragranuloma, nodular
C0019829|HL
C0019829|Hodgkin's lymphoma NOS
C0019829|Malignant lymphogranulomatosis
C0019829|Hodgkins sarcoma
C0023448|Lymphoid Leukemias
C0023448|Leukemias, Lymphocytic
C0023448|Leukemias, Lymphoid
C0023448|Lymphocytic Leukemias
C0023448|LEUKEMIA LYMPHATIC
C0023448|LEUKEMIA LYMPHOCYTIC
C0023448|LEUKEMIA LYMPHOID
C0023448|Lymphoid leukemia
C0023448|lymphocytic leukemia
C0023448|Lymphoid leukaemia
C0023448|Lymphoid leukaemia, unspecified
C0023448|Lymphoid leukemia, unspecified
C0023448|Leukemia, Lymphoid
C0023448|lymphatic leukemia
C0023448|lymphoblastic leukemia
C0023448|lymphogenous leukemia
C0023448|lymphocytic leukemia (diagnosis)
C0023448|Lymphoid leukaemia, no ICD-O subtype
C0023448|Lymphoid leukemia, no ICD-O subtype
C0023448|Lymphocytic leukaemia
C0023448|Lymphoid leukemia NOS
C0023448|Leukemia, Lymphocytic
C0023448|Leukemia, Lymphoid [Disease/Finding]
C0023448|[M]Lymphoid leukaemias
C0023448|[M]Lymphoid leukemias
C0023448|Lymphoid leukemia, disease (disorder)
C0023448|Lymphoid leukaemia NOS
C0023448|Lymphoid leukemia NOS (disorder)
C0023448|[M]Lymphoid leukemias (morphologic abnormality)
C0023448|Lymphoid leukemia, no ICD-O subtype (morphologic abnormality)
C0023448|Lymphoid leukemia, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0023448|Lymphoid leukemia, no International Classification of Diseases for Oncology subtype
C0023448|LEUKEMIA, LYMPHOCYTIC, MALIGNANT
C0023448|[M]Lymphoid leukemia NOS
C0023448|[M]Lymphoid leukaemia NOS
C0023448|Leukaemia lymphocytic
C0023448|Leukaemia lymphoid
C0023448|Unspecified lymphoid leukemia
C0023448|Lymphoblastic leukemia NOS
C0023448|Lymphatic leukaemia
C0023448|Leukaemia lymphatic
C0023448|Lymphoblastic leukaemia NOS
C0023448|Unspecified lymphoid leukaemia
C0023448|Aleukaemic lymphatic leukaemia [obs]
C0023448|Aleukaemic lymphocytic leukaemia [obs]
C0023448|Aleukaemic lymphoid leukaemia [obs]
C0023448|Aleukemic lymphatic leukemia [obs]
C0023448|Aleukemic lymphocytic leukemia [obs]
C0023448|Aleukemic lymphoid leukemia [obs]
C0023448|Lymphoid leukemia (disorder)
C0023448|Lymphosarcoma cell leukaemia [obs]
C0023448|Lymphosarcoma cell leukemia [obs]
C0023448|leukemia; lymphatic
C0023448|leukemia; lymphoblastic
C0023448|lymphatic; leukemia
C0023448|lymphoblastic; leukemia
C0023448|Lymphatic leukemia, NOS
C0023448|Lymphocytic leukemia, NOS
C0023448|Lymphoid leukemia, NOS
C0023448|Lymphoid leukemia, disease [Ambiguous]
C0598894|Monocytic leukemia
C0598894|LEUKEMIA MONOCYTIC
C0598894|Monocytic leukaemia
C0598894|Monocytic leukaemia, unspecified
C0598894|Monocytic leukemia, unspecified
C0598894|Schilling's leukemia
C0598894|monocytic leukemia (diagnosis)
C0598894|Monocytic leukaemia -RETIRED-
C0598894|Monocytic leukemia -RETIRED-
C0598894|monocytoid leukemia
C0598894|Monocytic leukemia, unspecified NOS
C0598894|Monocytic leukemia (morphologic abnormality)
C0598894|Monocytic leukemia NOS
C0598894|[M]Monocytic leukaemias
C0598894|Monocytic leukemia (disorder)
C0598894|[M]Monocytic leukemias
C0598894|[M]Monocytic leukaemia NOS
C0598894|[M]Monocytic leukemias (morphologic abnormality)
C0598894|Monocytic leukemia NOS (disorder)
C0598894|[M]Monocytic leukaemia NOS (disorder)
C0598894|Monocytic leukaemia NOS
C0598894|[M]Monocytic leukemia NOS
C0598894|Leukaemia monocytic NOS
C0598894|Unspecified monocytic leukemia
C0598894|Leukemia monocytic NOS
C0598894|Unspecified monocytic leukaemia
C0598894|Leukaemia monocytic
C0598894|Schilling-type monocytic leukemia
C0598894|Schilling-type monocytic leukaemia
C0598894|leukemia; monocytic
C0598894|monocytic; leukemia
C0598894|Monocytic leukemia, NOS
C0023470|Myeloid Leukemias
C0023470|Granulocytic Leukemias
C0023470|Leukemia, Myeloid
C0023470|Leukemias, Granulocytic
C0023470|Leukemias, Myelocytic
C0023470|Leukemias, Myelogenous
C0023470|Leukemias, Myeloid
C0023470|Myelocytic Leukemias
C0023470|Myelogenous Leukemias
C0023470|Myeloid Leukemia
C0023470|LEUKEMIA GRANULOCYTIC
C0023470|LEUKEMIA MYELOGENOUS
C0023470|LEUKEMIA MYELOID
C0023470|myelogenous leukemia
C0023470|Myeloid leukaemia
C0023470|Myeloid leukaemia, unspecified
C0023470|Myeloid leukemia, unspecified
C0023470|myelocytic leukemia
C0023470|myelosis
C0023470|granulocytic leukemia
C0023470|myeloid granulocytic leukemia
C0023470|myelogenous leukemia (diagnosis)
C0023470|Myeloid leukemia - category
C0023470|Myeloid leukaemia - category
C0023470|Leukemic granulocytic
C0023470|Myeloid leukemia, unspecified NOS
C0023470|Leukemia, Granulocytic
C0023470|Leukemia, Myelocytic
C0023470|Leukemia, Myelogenous
C0023470|Leukemia, Myeloid [Disease/Finding]
C0023470|Myeloid leukemia NOS (disorder)
C0023470|Myeloid leukaemia NOS
C0023470|Myeloid leukemia NOS
C0023470|[M]Myeloid leukemias (morphologic abnormality)
C0023470|[M]Myeloid leukaemias
C0023470|Myeloid leukemia, disease (disorder)
C0023470|[M]Myeloid leukemias
C0023470|Granulocytic leukemia (disorder)
C0023470|Myeloid leukemia, no ICD-O subtype (morphologic abnormality)
C0023470|Myeloid leukemia, no International Classification of Diseases for Oncology subtype
C0023470|Myeloid leukemia, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0023470|LEUKEMIA, GRANULOCYTIC, MALIGNANT
C0023470|[M]Myeloid leukaemia NOS
C0023470|[M]Myeloid leukemia NOS
C0023470|Non-lymphoblastic Leukemia
C0023470|Non-lymphocytic Leukemia
C0023470|Leukemia granulocytic NOS
C0023470|Non-lymphoblastic leukemia NOS
C0023470|Unspecified myeloid leukemia
C0023470|Leukaemia granulocytic
C0023470|Myelocytic leukaemia
C0023470|Unspecified myeloid leukaemia
C0023470|Leukaemia myelogenous
C0023470|Leukaemia myeloid
C0023470|Non-lymphoblastic leukaemia NOS
C0023470|Leukaemia granulocytic NOS
C0023470|Granulocytic leukaemia
C0023470|Aleukaemic monocytic leukaemia [obs]
C0023470|Aleukemic monocytic leukemia [obs]
C0023470|Myelogenous leukaemia
C0023470|Myeloid leukaemia (category)
C0023470|Myeloid leukemia (category)
C0023470|Myeloid leukemia (disorder)
C0023470|Myeloid leukemia - category (morphologic abnormality)
C0023470|Non-lymphocytic leukaemia
C0023470|granulocytic; leukemia
C0023470|leukemia; granulocytic
C0023470|leukemia; myelocytic
C0023470|leukemia; myeloid
C0023470|myelocytic; leukemia
C0023470|myeloid; leukemia
C0023470|Granulocytic leukemia, NOS
C0023470|Myelocytic leukemia, NOS
C0023470|Myelogenous leukemia, NOS
C0023470|Myeloid leukemia, NOS
C0023470|Myeloid leukaemia, NOS
C0023470|Myeloid leukemia, disease [Ambiguous]
C0023470|Myeloid leukemia, morphology (morphologic abnormality)
C0348394|Diffuse non-Hodgkin's lymphoma, unspecified
C0348394|Diffuse non-Hodgkin's lymphoma
C0348394|Diffuse non-Hodgkin lymphoma
C0348394|Nonfollicular lymphoma
C0348394|[X]Diffuse non-Hodgkin's lymphoma, unspecified (disorder)
C0348394|[X]Diffuse non-Hodgkin's lymphoma, unspecified
C0348394|Diffuse non-Hodgkin's lymphoma (disorder)
C0024301|Brill Symmers Disease
C0024301|Follicular Lymphomas
C0024301|Follicular Lymphomas, Giant
C0024301|Giant Follicular Lymphomas
C0024301|Lymphoma, Follicular
C0024301|Lymphomas, Follicular
C0024301|Lymphomas, Giant Follicular
C0024301|Lymphomas, Nodular
C0024301|Nodular Lymphomas
C0024301|Disease, Brill-Symmers
C0024301|Nodular Lymphoma
C0024301|Follicular [nodular] non-Hodgkin's lymphoma
C0024301|Follicular non-Hodgkin's lymphoma, unspecified
C0024301|Follicular non-Hodgkin lymphoma
C0024301|GIANT FOLLIC LYMPHOMA
C0024301|FOLLIC LYMPHOMA
C0024301|FOLLIC LYMPHOMA GIANT
C0024301|LYMPHOMA FOLLIC
C0024301|LYMPHOMA GIANT FOLLIC
C0024301|BRILL SYMMERS DIS
C0024301|follicular lymphoma
C0024301|nodular malignant lymphoma (diagnosis)
C0024301|nodular malignant lymphoma
C0024301|Malignant lymphoma, centroblastic-centrocytic, follicular -RETIRED-
C0024301|giant follicular lymphosarcoma (diagnosis)
C0024301|nodular lymphosarcoma
C0024301|giant follicular lymphosarcoma
C0024301|nodular lymphosarcoma (diagnosis)
C0024301|Follicular lymphoma, unspecified
C0024301|Lymphoma, Nodular
C0024301|Brill-Symmers Disease
C0024301|Lymphoma, Giant Follicular
C0024301|Lymphoma, Follicular [Disease/Finding]
C0024301|Follicular Lymphoma, Giant
C0024301|Giant Follicular Lymphoma
C0024301|follicular lymphoma (diagnosis)
C0024301|malignant neoplasm nodular lymphoma follicular
C0024301|(Nodular lymphoma: Brill-Symmers disease) or (reticulosarcoma - follicular or nodular) (disorder)
C0024301|Nodular lymphoma NOS (disorder)
C0024301|Follicular lymphoma NOS
C0024301|Follicular lymphoma: [non-Hodgkin's] or [NOS] (disorder)
C0024301|Nodular lymphoma (Brill - Symmers disease)
C0024301|[M]Malignant lymphoma, centroblastic-centrocytic, follicular
C0024301|(Nodular lymphoma: Brill-Symmers disease) or (reticulosarcoma - follicular or nodular)
C0024301|Nodular lymphoma of unspecified site
C0024301|[M]Malignant lymphoma, centroblastic-centrocytic, follicular (morphologic abnormality)
C0024301|[M]Malignant lymphoma, nodular NOS (& [Brill - Symmers' disease])
C0024301|[M]Malignant lymphoma, nodular NOS
C0024301|[M]Follicular lymphosarcoma NOS
C0024301|[M]Malignant lymphoma, nodular NOS (& [Brill - Symmers' disease]) (disorder)
C0024301|[M]Giant follicular lymphoma
C0024301|Nodular lymphoma NOS
C0024301|Follicular non-Hodgkin's lymphoma
C0024301|[M]Brill - Symmers' disease
C0024301|Follicular lymphoma: [non-Hodgkin's] or [NOS]
C0024301|Malignant lymphoma, centroblastic-centrocytic, follicular (morphologic abnormality)
C0024301|Nodular lymphoma of unspecified site (disorder)
C0024301|Reticulosarcoma - follicular or nodular
C0024301|Malignant lymphoma, centroblastic-centrocytic, follicular
C0024301|[M]Malignant lymphoma, nodular NOS (morphologic abnormality)
C0024301|[M]Nodular lymphosarcoma NOS
C0024301|follicular malignant lymphoma - centroblastic-centrocytic
C0024301|malignant neoplasm lymphoma follicular - centroblastic-centrocytic
C0024301|malignant neoplasm lymphoma b-cell low grade follicular
C0024301|follicular malignant lymphoma - centroblastic-centrocytic (diagnosis)
C0024301|Follicular low grade B-cell lymphoma (diagnosis)
C0024301|Follicular low grade B-cell lymphoma
C0024301|LYMPHOMA, FOLLICULAR, MALIGNANT
C0024301|Lymphoma, Follicular Centre Cell
C0024301|Follicular Centre Cell Lymphoma
C0024301|Follicle Center Lymphoma
C0024301|Nodular (follicular) lymphoma
C0024301|Malignant lymphoma, nodular
C0024301|Malignant lymphoma, follicular
C0024301|Follicular lymphosarcoma
C0024301|Brill - Symmers' disease
C0024301|Germinoblastoma, follicular
C0024301|Follicular low grade B-cell lymphoma (disorder)
C0024301|Follicular lymphoma (morphologic abnormality)
C0024301|Follicular non-Hodgkin's lymphoma (disorder)
C0024301|Malignant lymphoma, centroblastic-centrocytic, follicular (disorder)
C0024301|Malignant lymphoma, follicle center, follicular
C0024301|Malignant lymphoma, follicle center
C0024301|Malignant lymphoma, follicle centre, follicular
C0024301|Malignant lymphoma, follicle centre
C0024301|Malignant lymphoma, lymphocytic, nodular
C0024301|Nodular lymphoma (disorder)
C0024301|follicular; germinoblastoma
C0024301|follicular; lymphosarcoma
C0024301|germinoblastoma; follicular
C0024301|Brill-Symmers
C0024301|lymphocytic; lymphoma, nodular
C0024301|lymphoma; follicular
C0024301|lymphoma; lymphocytic, nodular
C0024301|lymphoma; nodular, lymphocytic
C0024301|lymphoma; nodular
C0024301|lymphosarcoma; follicular
C0024301|nodular; lymphoma, lymphocytic
C0024301|nodular; lymphoma
C0024301|Malignant lymphoma, follicular, NOS
C0024301|Malignant lymphoma, lymphocytic, nodular, NOS
C0024301|Malignant lymphoma, nodular, NOS
C0024301|Nodular lymphocytic lymphoma
C1264191|Malignant immunoproliferative disease, unspecified
C1264191|Malignant immunoproliferative diseases
C1264191|Malignant immunoproliferative disease
C1264191|malignant immunoproliferative disease (diagnosis)
C1264191|Malignant immunoproliferative disease (clinical)
C1264191|Malignant immunoproliferative disease (disorder)
C0494174|Multiple myeloma and malignant plasma cell neoplasms
C0494176|Other and unspecified malignant neoplasms of lymphoid, haematopoietic and related tissue
C0494176|Other and unspecified malignant neoplasms of lymphoid, hematopoietic and related tissue
C0494172|Other and unspecified types of non-Hodgkin's lymphoma
C0494172|Other specified and unspecified types of non-Hodgkin lymphoma
C0494175|Other leukaemias of specified cell type
C0494175|Other leukemias of specified cell type
C0456860|Peripheral and cutaneous T-cell lymphomas
C0456860|malignant neoplasm lymphoma cutaneous / peripheral t-cell
C0456860|cutaneous / peripheral T-cell lymphoma
C0456860|cutaneous / peripheral T-cell lymphoma (diagnosis)
C0456860|Cutaneous/peripheral T-cell lymphoma
C0456860|Cutaneous/peripheral T-cell lymphoma (disorder)
C2853945|Non-follicular lymphoma
C0079774|Lymphoma, Peripheral T-Cell
C0079774|Lymphoma, T-Cell, Peripheral
C0079774|Lymphomas, Peripheral T-Cell
C0079774|Peripheral T Cell Lymphoma
C0079774|Peripheral T-Cell Lymphomas
C0079774|T Cell Lymphoma, Peripheral
C0079774|T-Cell Lymphomas, Peripheral
C0079774|Peripheral T-cell lymphoma
C0079774|Mature T-Cell and NK-Cell Non-Hodgkin's Lymphoma
C0079774|Mature T-Cell and NK-Cell Non-Hodgkin Lymphoma
C0079774|mature T-cell lymphoma
C0079774|mature T-cell lymphoma (diagnosis)
C0079774|Peripheral T-cell lymphoma, no ICD-O subtype
C0079774|Peripheral T-Cell Lymphoma, Not Otherwise Specified
C0079774|Peripheral T-Cell Lymphoma, NOS
C0079774|Mature T/NK-cell lymphomas, unspecified
C0079774|Mature T/NK-cell lymphomas
C0079774|Lymphoma, T-Cell, Peripheral [Disease/Finding]
C0079774|T-Cell Lymphoma, Peripheral
C0079774|Lymphoma, T Cell, Peripheral
C0079774|[M] Peripheral T-cell lymphoma NOS (morphologic abnormality)
C0079774|Peripheral T-cell lymphoma (disorder)
C0079774|[M] Peripheral T-cell lymphoma NOS
C0079774|mature NK/T-cell lymphoma (diagnosis)
C0079774|mature NK/T-cell lymphoma
C0079774|malignant neoplasm lymphoma mature nk/t-cell
C0079774|Peripheral T-cell lymphoma, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0079774|Peripheral T-cell lymphoma, no ICD-O subtype (morphologic abnormality)
C0079774|Peripheral T-cell lymphoma, no International Classification of Diseases for Oncology subtype
C0079774|Peripheral T-cell lymphoma unspecified
C0079774|Peripheral T-cell lymphoma unspecified NOS
C0079774|Peripheral T-cell lymphoma (clinical)
C0079774|T-cell; lymphoma, peripheral
C0079774|lymphoma; T-cell, peripheral
C0079774|lymphoma; peripheral T-cell
C0079774|peripheral; T-cell lymphoma
C0079774|Mature T-Cell Non-Hodgkin's Lymphoma
C0079774|Mature T-Cell and NK-Cell Lymphoma
C0079774|Mature T-and NK-Cell Lymphoma
C0079774|PTCL
C0079774|Peripheral T-cell lymphoma (morphologic abnormality)
C2854064|Other specified types of T/NK-cell lymphoma
C2854069|Malignant immunoproliferative diseases and certain other B-cell lymphomas
C0085165|Bovine Leukoses
C0085165|Bovine Leukoses, Enzootic
C0085165|Bovine Leukosis, Enzootic
C0085165|Enzootic Bovine Leukoses
C0085165|Enzootic Bovine Leukosis
C0085165|Leukoses, Bovine
C0085165|Leukoses, Enzootic Bovine
C0085165|Leukosis, Enzootic Bovine
C0085165|Bovine Leukosis
C0085165|Enzootic Bovine Leukosis [Disease/Finding]
C0085165|Leukosis, Bovine
C0085165|Bovine viral leukosis
C0085165|Bovine viral leukosis (disorder)
C0085165|Malignant lymphoma of cattle
C0152276|Myeloid sarcoma
C0152276|Chloroma
C0152276|Sarcomas, Myeloid
C0152276|Myeloid Sarcomas
C0152276|Sarcoma, Myeloid
C0152276|Myeloid sarcoma, morphology
C0152276|Myeloid sarcoma, disease
C0152276|chloroma (diagnosis)
C0152276|granulocytic sarcoma (diagnosis)
C0152276|leukemia myeloid sarcoma
C0152276|leukemia myeloid sarcoma granulocytic sarcoma
C0152276|granulocytic sarcoma
C0152276|myeloid sarcoma (diagnosis)
C0152276|leukemia myeloid sarcoma chloroma
C0152276|Myeloid sarcoma NOS
C0152276|Myeloid Cell Tumor, Extramedullary
C0152276|Extramedullary Myeloid Cell Tumor
C0152276|Sarcoma, Granulocytic
C0152276|Sarcoma, Myeloid [Disease/Finding]
C0152276|Chloromas
C0152276|Granulocytic Sarcomas
C0152276|Sarcomas, Granulocytic
C0152276|Myeloid sarcoma NOS (disorder)
C0152276|SARCOMA, GRANULOCYTIC, MALIGNANT
C0152276|SARCOMA, MYELOID, MALIGNANT
C0152276|[M]Myeloid sarcoma
C0152276|[M]Chloroma
C0152276|[M]Granulocytic sarcoma
C0152276|Extramedullary Myeloid Tumor
C0152276|Chloroma (disorder)
C0152276|Granulocytic sarcoma (disorder)
C0152276|Myeloid sarcoma, disease (disorder)
C0152276|Myeloid sarcoma, morphology (morphologic abnormality)
C0152276|myelosarcoma
C0152276|granulocytic; sarcoma
C0152276|myeloid; sarcoma
C0152276|sarcoma; granulocytic
C0152276|sarcoma; myeloid
C0348393|Malignant neoplasm of lymphoid, haematopoietic and related tissue, unspecified
C0348393|Malignant neoplasm of lymphoid, hematopoietic and related tissue, unspecified
C0348393|Malignant neoplasms of lymphoid, haematopoietic and related tissue
C0348393|Malignant neoplasms of lymphoid, hematopoietic and related tissue
C0348393|Cancer of lymphatic and hematopoietic tissue
C0348393|Malignant neoplasms of lymphoid, hematopoietic and related tissue (C81-C96)
C0348393|Malignant tumor of lymphoid hemopoietic and related tissue
C0348393|Malig neoplm of lymphoid, hematpoetc and rel tissue, unsp
C0348393|[X]Malignant neoplasm of lymphoid, haematopoietic and related tissue, unspecified
C0348393|Malignant neoplasm of lymphatic and hemopoietic tissue
C0348393|[X]Malignant neoplasms of lymphoid, hematopoietic and related tissue (disorder)
C0348393|[X]Malignant neoplasms of lymphoid, hematopoietic and related tissue
C0348393|[X]Malignant neoplasm of lymphoid, hematopoietic and related tissue, unspecified
C0348393|[X]Malignant neoplasm of lymphoid, hematopoietic and related tissue, unspecified (disorder)
C0348393|[X]Malignant neoplasms of lymphoid, haematopoietic and related tissue
C0348393|Malignant neoplasm of lymphatic and haemopoietic tissue
C0348393|malignant neoplasm of lymphoid, hemopoietic and/or related tissue (diagnosis)
C0348393|malignant neoplasm of lymphoid, hemopoietic and/or related tissue
C0348393|Malignant tumor of lymphoid, hemopoietic AND/OR related tissue
C0348393|Malignant tumour of lymphoid haemopoietic and related tissue
C0348393|hematopoietic/lymphoid cancer
C0348393|Malignant tumor of lymphoid, hemopoietic AND/OR related tissue (disorder)
C0348393|Malignant tumor of lymphoid hemopoietic and related tissue (disorder)
C0348393|MALIGNANT NEOPLASM OF LYMPHATIC AND HEMATOPOIETIC TISSUE
C0021071|alpha Chain Disease
C0021071|Immunoproliferative Small Intestinal Disease
C0021071|Disease, alpha-Chain
C0021071|Diseases, alpha-Chain
C0021071|alpha-Chain Diseases
C0021071|Alpha heavy chain disease
C0021071|ALPHA CHAIN DIS
C0021071|HEAVY CHAIN DIS IGA TYPE
C0021071|IMMUNOPROLIFERATIVE SMALL INTESTINAL DIS
C0021071|Mediterraneanl Lymphoma
C0021071|Alpha heavy chain disease, NOS
C0021071|immunoproliferative small intestinal disease (diagnosis)
C0021071|Alpha heavy chain disease -RETIRED-
C0021071|immunoproliferative intestinal disease
C0021071|Mediterranean lymphoma
C0021071|Immunoproliferative Small Intestinal Disease [Disease/Finding]
C0021071|Lymphoma, Mediterranean
C0021071|Heavy Chain Disease, IgA Type
C0021071|alpha-Chain Disease
C0021071|IPSID
C0021071|[M] Immunoproliferative small intestinal disease
C0021071|[M] Alpha heavy chain disease
C0021071|Alpha heavy chain disease (disorder)
C0021071|[M] Alpha heavy chain disease (morphologic abnormality)
C0021071|[M] Immunoproliferative small intestinal disease (morphologic abnormality)
C0021071|Alpha heavy chain disease (diagnosis)
C0021071|Alpha heavy chain disease, enteric form (diagnosis)
C0021071|heavy chain disease alpha, enteric form
C0021071|Alpha heavy chain disease, enteric form
C0021071|heavy chain disease alpha
C0021071|Immunoproliferative small intestinal disease (clinical)
C0021071|Immunoproliferative small intestinal disease (disorder)
C0021071|Immunoproliferative small intestinal disease (morphologic abnormality)
C0021071|Alpha heavy chain disease (clinical)
C0021071|Alpha heavy chain disease, enteric form (disorder)
C0021071|Mediterranean lymphoma (clinical)
C0021071|IgA heavy chain disease
C0021071|disease (or disorder); alpha heavy chain
C0021071|disease (or disorder); heavy chain, alpha
C0021071|disease (or disorder); immunoproliferative, small intestine
C0021071|disease; alpha heavy chain
C0021071|heavy chain alpha
C0021071|lymphoma; mediterranean
C0021071|mediterranean; lymphoma
C0021071|alpha heavy chain; disease
C0021071|alpha; alpha heavy chain disease
C0021071|IgA heavy chain disease, NOS
C0021071|Alpha heavy chain disease [dup] (disorder)
C0021071|Mediterranean Abdominal Lymphoma
C0021071|immunoproliferative; disease, small intestine
C0376545|Hematologic Neoplasm
C0376545|Hematologic Neoplasms
C0376545|Hematological Malignancy
C0376545|Hematological Neoplasm
C0376545|Malignancies, Hematological
C0376545|Malignancy, Hematological
C0376545|Neoplasm, Hematologic
C0376545|Neoplasm, Hematological
C0376545|Neoplasms, Hematological
C0376545|Haematological malignancy
C0376545|NEOPL HEMATOL
C0376545|MALIGNANCY HEMATOL
C0376545|HEMATOL NEOPL
C0376545|HEMATOL MALIGNANCY
C0376545|MALIGNANCIES HEMATOL
C0376545|HEMATOL MALIGNANCIES
C0376545|Hematologic Malignancy
C0376545|Malignancy, Hematologic
C0376545|Hematologic Malignancies
C0376545|Hematological Neoplasms
C0376545|Hematological Malignancies
C0376545|Hematologic Neoplasms [Disease/Finding]
C0376545|Malignancies, Hematologic
C0376545|Neoplasms, Hematologic
C0376545|Carcinoma;blood
C0376545|Carcinoma;bone;marrow
C0376545|blood cancer
C0376545|Hematologic malignancy (disorder)
C0376545|Haematologic malignancy
C0376545|hematologic cancer
C0376545|Haematologic neoplasm
C0376545|Hematologic neoplasm (disorder)
C0376545|Hematological Tumor
C0376545|Malignant Hematologic Neoplasm
C0018854|Franklins Disease
C0018854|Franklin's disease
C0018854|gamma Chain Disease
C0018854|gamma-Chain Diseases
C0018854|Gamma heavy chain disease
C0018854|FRANKLINS DIS
C0018854|FRANKLIN DIS
C0018854|Gamma heavy chain disease -RETIRED-
C0018854|Franklin disease
C0018854|Gamma heavy chain disease (disorder)
C0018854|[M] Gamma heavy chain disease
C0018854|Gamma heavy chain disease (morphologic abnormality)
C0018854|[M] Gamma heavy chain disease (morphologic abnormality)
C0018854|:: Gamma heavy chain disease
C0018854|heavy chain disease gamma
C0018854|Gamma heavy chain disease (diagnosis)
C0018854|Gamma heavy chain disease (clinical)
C0018854|Franklin
C0018854|disease; gamma heavy chain
C0018854|gamma heavy chain; disease
C0018854|heavy chain gamma
C0018854|IgG heavy chain disease
C0018854|Gamma heavy chain disease [dup] (disorder)
C0018854|gamma-Chain Disease
C0543670|malignant white blood cell disorder
C0543670|malignant white blood cell disorder (diagnosis)
C0543670|malignant neoplasm white blood cell disorder
C0543670|Malignant white blood cell disorder (disorder)
C0474969|Malignant neoplasm of lymphatic or hematopoietic tissue otherwise specified (disorder)
C0474969|Malignant neoplasm of lymphatic or hematopoietic tissue otherwise specified
C0474969|Malignant neoplasm of lymphatic or haematopoietic tissue otherwise specified
C0474970|lymphatic/hematopoietic neoplasm
C0474970|neoplasm of lymphatic or hematopoietic tissue
C0474970|Malignant neoplasm lymphatic or haematopoietic tissue NOS
C0474970|Malignant neoplasm lymphatic or hematopoietic tissue NOS (disorder)
C0474970|Malignant neoplasm lymphatic or hematopoietic tissue NOS
C0474970|malignant lymphatic/hematopoietic neoplasm (diagnosis)
C0474970|malignant lymphatic/hematopoietic neoplasm
C0348391|Other malignant immunoproliferative diseases
C0348391|[X]Other malignant immunoproliferative diseases
C0348391|[X]Other malignant immunoproliferative diseases (disorder)
C0348392|Other specified malignant neoplasms of lymphoid, haematopoietic and related tissue
C0348392|Other specified malignant neoplasms of lymphoid, hematopoietic and related tissue
C0348392|Oth malig neoplm of lymphoid, hematpoetc and related tissue
C0348392|[X]Other specified malignant neoplasms of lymphoid, hematopoietic and related tissue (disorder)
C0348392|[X]Other specified malignant neoplasms of lymphoid, hematopoietic and related tissue
C0348392|[X]Other specified malignant neoplasms of lymphoid, haematopoietic and related tissue
C0024299|Lymphomas
C0024299|Germinoblastic Sarcomas
C0024299|Germinoblastomas
C0024299|Lymphoma
C0024299|Reticulolymphosarcomas
C0024299|Sarcomas, Germinoblastic
C0024299|Lymphomas, Malignant
C0024299|Malignant Lymphomas
C0024299|Germinoblastic Sarcoma
C0024299|Malignant Lymphoma
C0024299|Lymphoma (Hodgkin and Non-Hodgkin)
C0024299|Malignant lymphoma - category
C0024299|Malignant lymphoma (category)
C0024299|malignant lymphoma (diagnosis)
C0024299|Malignant lymphoma, no ICD-O subtype
C0024299|Lymphoma NOS
C0024299|Malignant lymphoma NOS
C0024299|Germinoblastoma
C0024299|Reticulolymphosarcoma
C0024299|Sarcoma, Germinoblastic
C0024299|Lymphoma, Malignant
C0024299|Lymphoma [Disease/Finding]
C0024299|Lymphomatous
C0024299|Malignant lymphoma NOS of unspecified site
C0024299|Malignant lymphoma NOS (disorder)
C0024299|[M]Reticulolymphosarcoma NOS
C0024299|[M]Malignant lymphoma NOS (disorder)
C0024299|Malignant lymphoma NOS of unspecified site (disorder)
C0024299|Lymphoma morphology
C0024299|[M]Malignant lymphoma NOS
C0024299|Lymphoma morphology (morphologic abnormality)
C0024299|Lymphosarcoma
C0024299|Malignant lymphoma, no ICD-O subtype (morphologic abnormality)
C0024299|Malignant lymphoma, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0024299|Malignant lymphoma, no International Classification of Diseases for Oncology subtype
C0024299|Lymphoma, NOS
C0024299|Lymphoma (Hodgkin's and Non-Hodgkin's)
C0024299|Lymphoma malignant
C0024299|Lymphoma (clinical)
C0024299|Malignant lymphoma (clinical)
C0024299|Malignant lymphoma (disorder)
C0024299|Malignant lymphoma - category (morphologic abnormality)
C0024299|Malignant lymphoma, NOS
C1306621|Primary malignant neoplasm of spleen
C1306621|splenic neoplasm malignant primary
C1306621|Primary malignant neoplasm of spleen (diagnosis)
C1306621|Primary malignant neoplasm of spleen (disorder)
C0040028|Essential Thrombocythemias
C0040028|Hemorrhagic Thrombocythemias
C0040028|Idiopathic Thrombocythemias
C0040028|Primary Thrombocythemias
C0040028|Thrombocythemias, Essential
C0040028|Thrombocythemias, Hemorrhagic
C0040028|Thrombocythemias, Idiopathic
C0040028|Thrombocythemias, Primary
C0040028|Essential Thrombocythemia
C0040028|Idiopathic Thrombocythemia
C0040028|hemorrhagic thrombocythemia
C0040028|Essential (haemorrhagic) thrombocythaemia
C0040028|Essential (hemorrhagic) thrombocythemia
C0040028|Essential thrombocythaemia
C0040028|Essential thrombocytosis
C0040028|Essential hemorrhagic thrombocythemia
C0040028|Idiopathic (hemorrhagic) thrombocythemia
C0040028|Primary thrombocytosis
C0040028|primary thrombocythemia
C0040028|Essential thrombocythaemia (clinical disorder)
C0040028|Essential thrombocythemia (clinical)
C0040028|essential thrombocytosis (diagnosis)
C0040028|essential thrombocythemia (diagnosis)
C0040028|primary thrombocytosis (diagnosis)
C0040028|idiopathic thrombocythemia (diagnosis)
C0040028|Idiopathic thrombocythaemia -RETIRED-
C0040028|Idiopathic thrombocythemia -RETIRED-
C0040028|essential hemorrhagic thrombocythemia (diagnosis)
C0040028|Thrombocythemia, Essential
C0040028|Ideopathic thrombocytosis
C0040028|Essntial thrombocythemia
C0040028|Idiopathic hemorrhagic thrombocythemia
C0040028|Thrombocythemia, Primary
C0040028|Thrombocythemia, Idiopathic
C0040028|Thrombocythemia, Essential [Disease/Finding]
C0040028|Thrombocythemia, Hemorrhagic
C0040028|Thrombocytosis;essential
C0040028|Thrombocytoses, Primary
C0040028|Primary Thrombocytoses
C0040028|Thrombocytosis, Primary
C0040028|Idiopathic thrombocythaemia
C0040028|Essential thrombocytosis (disorder)
C0040028|ET - Essential thrombocythaemia
C0040028|Essential thrombocythaemia (disorder)
C0040028|Idiopathic thrombocythemia (disorder)
C0040028|ET - Essential thrombocythemia
C0040028|Idiopathic thrombocythaemia (disorder)
C0040028|Idiopathic thrombocythemia (morphologic abnormality)
C0040028|[M]Idiopathic thrombocythaemia
C0040028|[M]Idiopathic thrombocythemia
C0040028|Primary thrombocythaemia
C0040028|Idiopathic thrombocytosis
C0040028|Essential haemorrhagic thrombocythaemia
C0040028|Idiopathic haemorrhagic thrombocythaemia
C0040028|Essential thrombocythemia (disorder)
C0040028|Essential thrombocythemia (morphologic abnormality)
C0040028|thrombocytosis; essential
C0040028|Essential thrombocythaemia (clinical)
C0040028|Essential Thrombocytemia
C0040028|Essential thrombocythemia (clinical disorder)
C3463824|Dysmyelopoietic Syndrome
C3463824|Myelodysplastic Syndromes
C3463824|Syndrome, Dysmyelopoietic
C3463824|Syndromes, Dysmyelopoietic
C3463824|Syndromes, Myelodysplastic
C3463824|Myelodysplastic Syndrome
C3463824|Syndrome, Myelodysplastic
C3463824|Myelodysplastic syndrome, unspecified
C3463824|Oligoblastic Leukemia
C3463824|Myelodysplasia
C3463824|Myelodysplastic syndrome (morphology) -Retired-
C3463824|Myelodysplastic syndrome (morphology)
C3463824|myelodysplasia (diagnosis)
C3463824|Myelodysplastic synd NOS
C3463824|Myelodysplastic Syndrome/Neoplasm
C3463824|Myelodysplastic Neoplasm
C3463824|Hematopoeitic - Myelodysplastic Syndrome (MDS)
C3463824|Myelodysplastic Syndromes [Disease/Finding]
C3463824|Dysmyelopoietic Syndromes
C3463824|MDS
C3463824|Preleukemia
C3463824|Smoldering leukemia
C3463824|[X]Myelodysplastic syndrome, unspecified
C3463824|Smouldering leukaemia
C3463824|Myelodysplastic syndrome (disorder)
C3463824|Preleukaemia
C3463824|Myelodysplastic syndrome (morphologic abnormality)
C3463824|Preleukemic syndrome
C3463824|Myelodysplasia (disorder)
C3463824|Preleukaemic syndrome
C3463824|[X]Myelodysplastic syndrome, unspecified (disorder)
C3463824|[M]Myelodysplastic syndrome
C3463824|myelodysplastic syndrome (diagnosis)
C3463824|Myelodysplastic syndrome, NOS
C3463824|MYELODYSPLASTIC SYNDROME, SUSCEPTIBILITY TO
C3463824|Myeloid dysplasia
C3463824|Myelodysplastic syndrome NOS
C3463824|MDS - Myelodysplastic syndrome
C3463824|Myelodysplastic syndrome (clinical)
C3463824|dysmyelopoiesis
C3463824|myelodysplastic; syndrome
C3463824|preleukemic; syndrome
C3463824|syndrome; myelodysplastic
C3463824|syndrome; preleukemic
C0019613|Disorder, Malignant Histiocytic
C0019613|Disorders, Malignant Histiocytic
C0019613|Histiocytic Disorder, Malignant
C0019613|Histiocytic Disorders, Malignant
C0019613|Malignant Histiocytic Disorder
C0019613|Malignant Histiocytic Disorders
C0019613|Histiocytic Disorders, Malignant [Disease/Finding]
C0019613|malig neoplasm histiocytic disorder
C0019613|malignant histiocytic disorder (diagnosis)
C0019613|Malignant histiocytic disorder (disorder)
C0341713|Leukemic infiltrate of kidney (diagnosis)
C0341713|Leukemic infiltrate of kidney
C0341713|renal neoplasm malignant leukemic infiltrate
C0341713|Leukaemic infiltrate of kidney
C0341713|Leukemic infiltrate of kidney (disorder)
C1301145|mast cell malignancy (diagnosis)
C1301145|Mast cell malignancy
C1301145|Mast cell malignancy (disorder)
C0024305|Lymphoma, Non Hodgkin's
C0024305|Lymphoma, Non-Hodgkin
C0024305|Lymphoma, Nonhodgkin
C0024305|Non Hodgkin's Lymphoma
C0024305|Non-Hodgkins Lymphoma
C0024305|Nonhodgkin's Lymphoma
C0024305|Non-Hodgkin's lymphoma, unspecified type
C0024305|Lymphoma, Non Hodgkin
C0024305|Lymphoma, Non Hodgkins
C0024305|Non Hodgkin Lymphoma
C0024305|Nonhodgkins Lymphoma
C0024305|Small cleaved cell (diffuse)
C0024305|Small cleaved cell (diffuse) non-Hodgkin's lymphoma
C0024305|LYMPHOMA, NON-HODGKIN, FAMILIAL
C0024305|Non-Hodgkin lymphoma
C0024305|NHL
C0024305|NONHODGKIN LYMPHOMA
C0024305|Non-Hodgkin's Lymphoma
C0024305|Diffuse Small Cleaved Cell Lymphoma
C0024305|LYMPHOMA SMALL CLEAVED DIFFUSE
C0024305|Small Cleaved Cell Lymphoma, Diffuse
C0024305|DIFFUSE SMALL CLEAVED LYMPHOMA
C0024305|SMALL CLEAVED LYMPHOMA DIFFUSE
C0024305|Malignant lymphoma, non-Hodgkin's, NOS
C0024305|non-Hodgkin's lymphoma (diagnosis)
C0024305|Non-Hodgkin lymphoma - category
C0024305|Malignant lymphoma, small cleaved cell, diffuse -RETIRED-
C0024305|Non-Hodgkin lymphoma, no ICD-O subtype
C0024305|Non-Hodgkin's Lymphoma (NHL)
C0024305|Non-Hodgkin lymphoma NOS
C0024305|Lymphoma, Nonhodgkins
C0024305|Lymphoma, Non-Hodgkin's
C0024305|Lymphoma, Nonhodgkin's
C0024305|Lymphoma, Non-Hodgkin [Disease/Finding]
C0024305|Lymphoma, Non-Hodgkins
C0024305|Small Cleaved-Cell Lymphoma, Diffuse
C0024305|Lymphoma, Atypical Diffuse Small Lymphoid
C0024305|Diffuse Small Cleaved-Cell Lymphoma
C0024305|Lymphoma, Small Cleaved Cell, Diffuse
C0024305|Lymphoma, Small Cleaved-Cell, Diffuse
C0024305|Lymphoma;non Hodgkins
C0024305|[X]Non-Hodgkin's lymphoma, unspecified type (disorder)
C0024305|[X]Non-Hodgkin's lymphoma, unspecified type
C0024305|Non-Hodgkin's lymphoma NOS
C0024305|[M]Malignant lymphoma, small cleaved cell, diffuse (morphologic abnormality)
C0024305|[M]Malignant lymphoma, small cleaved cell, diffuse
C0024305|Non-Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C0024305|Non-Hodgkin lymphoma, no ICD-O subtype (morphologic abnormality)
C0024305|Non-Hodgkin lymphoma, no International Classification of Diseases for Oncology subtype
C0024305|NHL, NOS
C0024305|Non-Hodgkin lymphoma, NOS
C0024305|[M]Non-Hodgkin's lymphoma
C0024305|[M]Malignant lymphoma, non-Hodgkin's type
C0024305|Lymphoma (non-Hodgkin's)
C0024305|Non-Hodgkin`s lymphoma
C0024305|Diffuse non-Hodgkin's small cleaved cell (diffuse) lymphoma
C0024305|Malignant lymphoma, non-Hodgkin's type
C0024305|NHL - Non-Hodgkin's lymphoma
C0024305|Malignant lymphoma, cleaved cell [obs]
C0024305|Malignant lymphoma, non-Hodgkin's
C0024305|Malignant lymphoma, non-Hodgkin
C0024305|Malignant lymphoma, small cell, noncleaved, diffuse [obs]
C0024305|Malignant lymphoma, small cleaved cell [obs]
C0024305|Malignant lymphoma, small cleaved cell, diffuse [obs]
C0024305|Malignant lymphoma, undifferentiated cell type [obs]
C0024305|Malignant lymphoma, undifferentiated cell, non-Burkitt [obs]
C0024305|Non-Hodgkin lymphoma (category)
C0024305|Non-Hodgkin lymphoma - category (morphologic abnormality)
C0024305|Non-Hodgkin's lymphoma (clinical)
C0024305|Non-Hodgkin's lymphoma (disorder)
C0024305|Non-Hodgkin's lymphoma - disorder
C0024305|diffuse; lymphoma, small cell, cleaved
C0024305|lymphoma; diffuse, small cell, cleaved
C0024305|lymphoma; non-Hodgkin's
C0024305|lymphoma; small cell, cleaved (diffuse)
C0024305|non-Hodgkin's; lymphoma
C0024305|small cell; lymphoma, cleaved (diffuse)
C0024305|Non-Hodgkin's lymphoma, NOS
C0024305|non hodgkins lymphoma
C1292778|Chronic myeloproliferative disease
C1292778|Myeloproliferative disease (chronic) NOS
C1292778|Chronic myeloproliferative disorder
C1292778|Chronic myeloproliferative disease -RETIRED-
C1292778|Chronic myeloproliferative disease, no ICD-O subtype
C1292778|MPN
C1292778|Myeloproliferative Disorder
C1292778|Myeloproliferative Neoplasm
C1292778|Chronic Myeloproliferative Neoplasm
C1292778|Myeloproliferative Tumor
C1292778|chronic myeloproliferative syndrome (diagnosis)
C1292778|chronic myeloproliferative syndrome
C1292778|myeloproliferative syndrome chronic
C1292778|Chronic myeloproliferative disease, no International Classification of Diseases for Oncology subtype
C1292778|Chronic myeloproliferative disease, no International Classification of Diseases for Oncology subtype (morphologic abnormality)
C1292778|Chronic myeloproliferative disease, no ICD-O subtype (morphologic abnormality)
C1292778|Myeloproliferative neoplasm, no ICD-O subtype
C1292778|Chronic myeloproliferative disorder (morphology)
C1292778|MPD
C1292778|Chronic myeloproliferative disorder (clinical) (disorder)
C1292778|Chronic myeloproliferative disorder (clinical)
C1292778|Chronic myeloproliferative disorder (morphologic abnormality)
C1292778|chronic myeloproliferative disorders
C1292778|disease (or disorder); myeloproliferative (chronic)
C1292778|myeloproliferative; disease (chronic)
C1292778|CMPD
C1292778|Chronic myeloproliferative disease (morphologic abnormality)
C1292778|Chronic myeloproliferative disease NOS
C1301355|Disease, Myeloproliferative-Myelodisplastic
C1301355|Diseases, Myeloproliferative-Myelodisplastic
C1301355|Myelodysplastic-Myeloproliferative Diseases
C1301355|Myelodysplastic-Myeloproliferative Disease
C1301355|Disease, Myelodysplastic-Myeloproliferative
C1301355|Myelodysplastic Myeloproliferative Diseases
C1301355|Myeloproliferative-Myelodisplastic Disease
C1301355|Diseases, Myelodysplastic-Myeloproliferative
C1301355|Myeloproliferative Myelodisplastic Diseases
C1301355|Myelodysplastic/Myeloproliferative Neoplasm
C1301355|Myelodysplastic/Myeloproliferative Disease
C1301355|MDS/MPN
C1301355|Myeloproliferative-Myelodisplastic Diseases
C1301355|Myelodysplastic-Myeloproliferative Diseases [Disease/Finding]
C1301355|Myelodysplastic/myeloproliferative disease (disorder)
C1301355|myelodysplastic / myeloproliferative disease
C1301355|myelodysplastic / myeloproliferative disease (diagnosis)
C1301355|bone marrow neoplasm myelodysplastic / myeloproliferative disease
C1301355|Myelodysplastic/myeloproliferative disease (morphologic abnormality)
C1301355|MDS/MPD
C1301355|myelodysplastic/myeloproliferative diseases
C1301355|MDS-MPD
C1301355|MPD-MDS
C1301355|MPD/MDS
C1301355|Myelodysplastic/Myeloproliferative Disorders
C1301355|Myelodysplastic/Myeloproliferative Disorder
C1301355|Myeloproliferative/Myelodysplastic Disorders
C1301355|Myeloproliferative/Myelodysplastic Syndromes
C0029812|Other specified leukaemias
C0029812|Other specified leukemias
C0029812|Other specified leukemia (disorder)
C0029812|Other specified leukemias NOS
C0029812|Other specified leukemia NOS (disorder)
C0029812|[X]Other specified leukaemias
C0029812|Other specified leukemia
C0029812|Other specified leukaemia
C0029812|Other specified leukemia NOS
C0029812|[X]Other specified leukemias
C0029812|[X]Other specified leukemias (disorder)
C0029812|Other specified leukaemia NOS
C1955727|Lymphosarcoma and reticulosarcoma and other specified malignant tumors of lymphatic tissue
C0153867|Multiple myeloma and immunoproliferative neoplasms
C0153867|Multiple myeloma and immunoproliferative disease
C0153867|Multiple myeloma and immunoproliferative disease (disorder)
C0153793|Other malignant neoplasms of lymphoid and histiocytic tissue
C0153793|Other malignant neoplasm of lymphoid and histiocytic tissue (disorder)
C0153793|Other malignant neoplasm of lymphoid and histiocytic tissue
C0432564|malignant neoplasm of lymphoid and histiocytic tissue
C0432564|malignant neoplasm of lymphoid and histiocytic tissue (diagnosis)
C0432564|Malignant neoplasm of lymphoid AND/OR histiocytic tissue -RETIRED-
C0432564|malignant tumor of lymphoid and histiocytic tissue
C0432564|Malignant neoplasm of lymphoid AND/OR histiocytic tissue
C0432564|Malignant neoplasm of lymphoid AND/OR histiocytic tissue (disorder)
C0432564|Unspecified malignant neoplasm of lymphoid and histiocytic tissue of unspecified site (disorder)
C0432564|Unspecified malignant neoplasm of lymphoid and histiocytic tissue of unspecified site
C0432564|Malignant neoplasms of lymphoid and histiocytic tissue NOS (disorder)
C0432564|Malignant neoplasms of lymphoid and histiocytic tissue NOS
C0432564|Malignant neoplasm of lymphoid and histiocytic tissue, NOS
C2217148|malignant neoplasm of lymphoid and histiocytic tissue of head, face, or neck (diagnosis)
C2217148|malignant neoplasm of lymphoid and histiocytic tissue of head, face, or neck
C2217148|malignant tumor of lymphoid and histiocytic tissue of head, face, or neck
C2217152|malignant neoplasm of lymphoid and histiocytic tissue of intrathoracic region (diagnosis)
C2217152|malignant neoplasm of lymphoid and histiocytic tissue of intrathoracic region
C2217152|malignant neoplasm of intrathoracic lymphoid and histiocytic tissue
C2217152|malignant tumor of lymphoid and histiocytic tissue of intrathoracic region
C2217150|malignant neoplasm of lymphoid and histiocytic tissue of intra-abdominal region (diagnosis)
C2217150|malignant neoplasm of lymphoid and histiocytic tissue of intra-abdominal region
C2217150|malignant neoplasm of intra-abdominal lymphoid and histiocytic tissue
C2217150|malignant tumor of lymphoid and histiocytic tissue of intra-abdominal region
C2217147|malignant neoplasm of lymphoid and histiocytic tissue of axilla or upper limb
C2217147|malignant neoplasm of lymphoid and histiocytic tissue of axilla or upper limb (diagnosis)
C2217147|malignant tumor of lymphoid and histiocytic tissue of axilla or upper limb
C2217149|malignant neoplasm of lymphoid and histiocytic tissue of inguinal region or lower limb (diagnosis)
C2217149|malignant neoplasm of lymphoid and histiocytic tissue of inguinal region or lower limb
C2217149|malignant tumor of lymphoid and histiocytic tissue of inguinal region or lower limb
C2217151|malignant neoplasm of lymphoid and histiocytic tissue of intrapelvic region (diagnosis)
C2217151|malignant neoplasm of lymphoid and histiocytic tissue of intrapelvic region
C2217151|malignant neoplasm of intrapelvic lymphoid and histiocytic tissue
C2217151|malignant tumor of lymphoid and histiocytic tissue of intrapelvic region
C2217154|malignant neoplasm of lymphoid and histiocytic tissue of spleen
C2217154|malignant neoplasm of lymphoid and histiocytic tissue of spleen (diagnosis)
C2217154|malignant neoplasm of splenic lymphoid and histiocytic tissue
C2217154|malignant tumor of lymphoid and histiocytic tissue of spleen
C2217153|malignant neoplasm of lymphoid and histiocytic tissue of multiple sites (diagnosis)
C2217153|malignant neoplasm of lymphoid and histiocytic tissue of multiple sites
C2217153|malignant tumor of lymphoid and histiocytic tissue of multiple sites
C0936223|Prostate cancer metastatic
C0936223|Metastatic Prostate Carcinoma
C0936223|Metastatic Prostate Cancer
C0936223|Carcinoma of the prostate metastatic
C0936223|Prostatic cancer metastatic
C0936223|Prostate Carcinoma Metastatic
C0278838|Prostate cancer recurrent
C0278838|Recurrent Prostate Cancer
C0278838|Recurrent Prostate Carcinoma
C0278838|Carcinoma of the prostate recurrent
C0278838|Prostatic cancer recurrent
C0278838|prostate cancer, recurrent
C0278838|Recurrent Cancer of Prostate
C0278838|Recurrent Cancer of the Prostate
C0854969|Prostate cancer stage 0
C0854969|Prostatic cancer stage 0
C0278834|Prostate cancer stage I
C0278834|Stage I Prostate Carcinoma
C0278834|Stage I Prostate Cancer AJCC v6
C0278834|Stage I Prostatic Cancer AJCC v6
C0278834|Prostate Carcinoma Stage I AJCC v6
C0278834|Prostate Cancer Stage I AJCC v6
C0278834|Stage I Prostate Carcinoma AJCC v6
C0278834|Cancer of Prostate Stage I AJCC v6
C0278834|Cancer of the Prostate Stage I AJCC v6
C0278834|Stage I Cancer of the Prostate AJCC v6
C0278834|Stage I Cancer of Prostate AJCC v6
C0278834|Stage I Prostatic Carcinoma AJCC v6
C0278834|stage I prostate cancer
C0278834|Prostatic cancer stage I
C0278834|Carcinoma of the prostate stage I
C0278834|cancer of the prostate, stage I
C0278834|carcinoma of the prostate, stage I
C0278834|prostate cancer, stage I
C0278834|stage I cancer of the prostate
C0278834|stage I carcinoma of the prostate
C0278835|Prostate cancer stage II
C0278835|Stage II Prostate Carcinoma
C0278835|Cancer of the Prostate Stage II AJCC v6
C0278835|Prostate Cancer Stage II AJCC v6
C0278835|Stage II Cancer of Prostate AJCC v6
C0278835|Stage II Cancer of the Prostate AJCC v6
C0278835|Stage II Prostate Carcinoma AJCC v6
C0278835|Prostate Carcinoma Stage II AJCC v6
C0278835|Stage II Prostate Cancer AJCC v6
C0278835|Stage II Prostatic Carcinoma AJCC v6
C0278835|Stage II Prostatic Cancer AJCC v6
C0278835|Cancer of Prostate Stage II AJCC v6
C0278835|stage II prostate cancer
C0278835|Prostatic cancer stage II
C0278835|Carcinoma of the prostate stage II
C0278835|cancer of the prostate, stage II
C0278835|carcinoma of the prostate, stage II
C0278835|prostate cancer, stage II
C0278835|stage II cancer of the prostate
C0278835|stage II carcinoma of the prostate
C0278836|Prostate cancer stage III
C0278836|Stage III Prostate Carcinoma
C0278836|Stage III Prostate Carcinoma AJCC v6
C0278836|Stage III Cancer of Prostate AJCC v6
C0278836|Cancer of Prostate Stage III AJCC v6
C0278836|Prostate Cancer Stage III AJCC v6
C0278836|Stage III Cancer of the Prostate AJCC v6
C0278836|Prostate Carcinoma Stage III AJCC v6
C0278836|Stage III Prostate Cancer AJCC v6
C0278836|Cancer of the Prostate Stage III AJCC v6
C0278836|Stage III Prostatic Cancer AJCC v6
C0278836|Stage III Prostatic Carcinoma AJCC v6
C0278836|stage III prostate cancer
C0278836|Carcinoma of the prostate stage III
C0278836|Prostatic cancer stage III
C0278836|cancer of the prostate, stage III
C0278836|carcinoma of the prostate, Stage III
C0278836|prostate cancer, stage III
C0278836|stage III cancer of the prostate
C0278836|stage III carcinoma of the prostate
C0278837|Prostate cancer stage IV
C0278837|Stage IV Prostate Carcinoma
C0278837|Stage IV Prostate Cancer AJCC v6
C0278837|Prostate Cancer Stage IV AJCC v6
C0278837|Stage IV Cancer of Prostate AJCC v6
C0278837|Stage IV Cancer of the Prostate AJCC v6
C0278837|Prostate Carcinoma Stage IV AJCC v6
C0278837|Stage IV Prostatic Cancer AJCC v6
C0278837|Cancer of Prostate Stage IV AJCC v6
C0278837|Cancer of the Prostate Stage IV AJCC v6
C0278837|Stage IV Prostate Carcinoma AJCC v6
C0278837|Stage IV Prostatic Carcinoma AJCC v6
C0278837|stage IV prostate cancer
C0278837|Carcinoma of the prostate stage IV
C0278837|Prostatic cancer stage IV
C0278837|cancer of the prostate, stage IV
C0278837|carcinoma of the prostate, stage IV
C0278837|prostate cancer, stage IV
C0278837|stage IV cancer of the prostate
C0278837|stage IV carcinoma of the prostate
C1297952|malignant neoplasm involving prostate by direct extension from bladder (diagnosis)
C1297952|prostate gland malignant by direct extension from bladder
C1297952|malignant neoplasm involving prostate by direct extension from bladder
C1297952|Malignant tumor involving prostate by direct extension from bladder (disorder)
C1297952|Malignant tumor involving prostate by direct extension from bladder
C1297952|Malignant tumour involving prostate by direct extension from bladder
C2007082|carcinosarcoma of prostate gland (diagnosis)
C2007082|carcinosarcoma of prostate gland
C2212269|malignant small cell neoplasm of prostate gland
C2212269|prostate gland neoplasm malignant small cell type
C2212269|malignant small cell neoplasm of prostate gland (diagnosis)
C2011401|giant cell type neoplasm of prostate gland (diagnosis)
C2011401|prostate gland neoplasm malignant giant cell type
C2011401|giant cell type neoplasm of prostate gland
C2018684|spindle cell type neoplasm of prostate gland
C2018684|spindle cell type neoplasm of prostate gland (diagnosis)
C2018684|prostate gland neoplasm malignant spindle cell type
C2075644|prostate gland neoplasm malignant clear cell type
C2075644|clear cell type neoplasm of prostate gland
C2075644|clear cell type neoplasm of prostate gland (diagnosis)
C0600139|CARCINOMA OF PROSTATE
C0600139|carcinoma of prostate gland
C0600139|carcinoma of prostate gland (diagnosis)
C0600139|prostatic carcinoma
C0600139|Carcinoma;prostate
C0600139|Cancer of prostate
C0600139|Carcinoma of prostate (disorder)
C0600139|Prostate cancer, NOS
C0600139|prostate cancer
C0600139|Prostate Carcinoma
C0600139|Carcinoma prostate
C0600139|Carcinoma prostatic
C0600139|CA - Carcinoma of prostate
C0600139|carcinoma, prostatic
C0600139|Cancer of the Prostate
C0600139|Carcinoma of the Prostate
C2212291|sarcoma of prostate gland (diagnosis)
C2212291|sarcoma of prostate gland
C2212294|fibrosarcoma of prostate gland
C2212294|fibrosarcoma of prostate gland (diagnosis)
C2212297|myosarcoma of prostate gland
C2212297|myosarcoma of prostate gland (diagnosis)
C2142688|marginal zone B-cell lymphoma of prostate gland
C2142688|marginal zone B-cell lymphoma of prostate gland (diagnosis)
C2217386|malignant neoplasm of prostate gland staging
C2217386|malignant neoplasm of prostate gland staging (diagnosis)
C2217386|malignant prostatic neoplasm staging
C2217386|prostatic cancer staging
C2217386|malignant tumor of prostate gland staging
C0007112|adenocarcinoma of prostate gland
C0007112|adenocarcinoma of prostate gland (diagnosis)
C0007112|prostatic adenocarcinoma
C0007112|Prostate adenocarcinoma
C0007112|Adenocarcinoma of prostate
C0007112|Adenocarcinoma of prostate (disorder)
C0007112|adenocarcinoma of the prostate
C0007112|adenocarcinoma, prostatic
C0007112|prostate cancer, adenocarcinoma
C2146665|acinar cell carcinoma of prostate gland (diagnosis)
C2146665|acinar cell carcinoma of prostate gland
C2146677|acinar cell cystadenocarcinoma of prostate gland
C2146677|prostate malignant carcinoma acinar cell cystadenocarcinoma
C2146677|acinar cell cystadenocarcinoma of prostate gland (diagnosis)
C2033179|papillary carcinoma in situ of prostate gland
C2033179|papillary carcinoma in situ of prostate gland (diagnosis)
C2142680|noninvasive papillary squamous cell carcinoma in situ of prostate gland
C2142680|prostate gland CIS papillary squamous cell noninvasive
C2142680|noninvasive papillary squamous cell carcinoma in situ of prostate gland (diagnosis)
C2019399|squamous cell carcinoma in situ of prostate gland
C2019399|squamous cell carcinoma in situ of prostate gland (diagnosis)
C2019400|squamous cell carcinoma in situ of prostate gland with questionable stromal invasion (diagnosis)
C2019400|prostate carcinoma in situ squamous cell with questionable stromal invasion
C2019400|squamous cell carcinoma in situ of prostate gland with questionable stromal invasion
C2145436|transitional cell carcinoma in situ of prostate gland
C2145436|transitional cell carcinoma in situ of prostate gland (diagnosis)
C2142681|noninvasive papillary transitional cell carcinoma in situ of prostate gland
C2142681|prostate gland CIS papillary transitional cell noninvasive
C2142681|noninvasive papillary transitional cell carcinoma in situ of prostate gland (diagnosis)
C2142714|noninfiltrating intraductal papillary adenocarcinoma in situ of prostate gland
C2142714|noninfiltrating intraductal papillary adenocarcinoma in situ of prostate gland (diagnosis)
C2142714|prostate noninfiltrating intraductal papillary adenocarcinoma in situ
C2142679|prostate gland CIS noninfiltrating intracystic carcinoma
C2142679|noninfiltrating intracystic carcinoma in situ of prostate gland
C2142679|noninfiltrating intracystic carcinoma in situ of prostate gland (diagnosis)
C2142677|prostate gland carcinoma in situ intraductal micropapillary
C2142677|intraductal micropapillary carcinoma in situ of prostate gland (diagnosis)
C2142677|intraductal micropapillary carcinoma in situ of prostate gland
C2212270|malignant epithelioma of prostate gland (diagnosis)
C2212270|malignant epithelioma of prostate gland
C2111662|large cell carcinoma of prostate gland
C2111662|large cell carcinoma of prostate gland (diagnosis)
C2111743|large cell neuroendocrine carcinoma of prostate gland (diagnosis)
C2111743|large cell neuroendocrine carcinoma of prostate gland
C2111663|large cell carcinoma of prostate gland with rhabdoid phenotype
C2111663|large cell carcinoma of prostate gland with rhabdoid phenotype (diagnosis)
C2111663|prostate malignant carcinoma large cell with rhabdoid phenotype
C2012107|glassy cell carcinoma of prostate gland
C2012107|glassy cell carcinoma of prostate gland (diagnosis)
C2188081|undifferentiated carcinoma of prostate gland
C2188081|undifferentiated carcinoma of prostate gland (diagnosis)
C2212271|anaplastic carcinoma of prostate gland
C2212271|anaplastic carcinoma of prostate gland (diagnosis)
C2082456|pleomorphic carcinoma of prostate gland (diagnosis)
C2082456|pleomorphic carcinoma of prostate gland
C2011261|giant cell carcinoma of prostate gland (diagnosis)
C2011261|giant cell carcinoma of prostate gland
C2018401|spindle cell carcinoma of prostate gland (diagnosis)
C2018401|spindle cell carcinoma of prostate gland
C2011226|giant cell and spindle cell carcinoma of prostate gland (diagnosis)
C2011226|giant cell and spindle cell carcinoma of prostate gland
C2011226|prostate malignant carcinoma giant cell and spindle cell
C2142931|pseudosarcomatous carcinoma of prostate gland (diagnosis)
C2142931|pseudosarcomatous carcinoma of prostate gland
C2111813|polygonal cell carcinoma of prostate gland
C2111813|polygonal cell carcinoma of prostate gland (diagnosis)
C2142712|carcinoma of prostate gland with osteoclast-like giant cells (diagnosis)
C2142712|carcinoma of prostate gland with osteoclast-like giant cells
C2142712|prostatic carcinoma with osteoclast-like giant cells
C2033229|papillary carcinoma of prostate gland
C2033229|papillary carcinoma of prostate gland (diagnosis)
C2033307|papillary squamous cell carcinoma of prostate gland (diagnosis)
C2033307|papillary squamous cell carcinoma of prostate gland
C2189358|verrucous carcinoma of prostate gland (diagnosis)
C2189358|verrucous carcinoma of prostate gland
C2109317|prostate malignant carcinoma squamous cell keratinizing
C2109317|keratinizing squamous cell carcinoma of prostate gland (diagnosis)
C2109317|keratinizing squamous cell carcinoma of prostate gland
C2212272|nonkeratinizing large cell squamous carcinoma cell of prostate gland
C2212272|prostate malignant carcinoma squamous cell large cell nonkeratinizing
C2212272|nonkeratinizing large cell squamous carcinoma cell of prostate gland (diagnosis)
C2212273|nonkeratinizing small cell squamous cell carcinoma of prostate gland (diagnosis)
C2212273|prostate malignant carcinoma squamous cell small cell nonkeratinizing
C2212273|nonkeratinizing small cell squamous cell carcinoma of prostate gland
C2018564|spindle cell squamous cell carcinoma of prostate gland (diagnosis)
C2018564|spindle cell squamous cell carcinoma of prostate gland
C2018564|prostate malignant carcinoma squamous cell spindle cell
C2212275|microinvasive squamous cell carcinoma of prostate gland (diagnosis)
C2212275|prostate malignant carcinoma squamous cell microinvasive
C2212275|microinvasive squamous cell carcinoma of prostate gland
C2019492|prostate malignant carcinoma squamous cell with horn formation
C2019492|squamous cell carcinoma of prostate gland with horn formation
C2019492|squamous cell carcinoma with horn formation of prostate gland
C2019492|squamous cell carcinoma of prostate gland with horn formation (diagnosis)
C2009885|fusiform type small cell carcinoma of prostate gland
C2009885|fusiform type small cell carcinoma of prostate gland (diagnosis)
C2182974|duct carcinoma, desmoplastic type, of prostate gland (diagnosis)
C2182974|duct carcinoma, desmoplastic type, of prostate gland
C2145466|transitional cell carcinoma of prostate gland (diagnosis)
C2145466|transitional cell carcinoma of prostate gland
C2018609|spindle cell transitional cell carcinoma of prostate gland (diagnosis)
C2018609|prostate malignant carcinoma transitional cell spindle cell
C2018609|spindle cell transitional cell carcinoma of prostate gland
C2212276|prostate gland malignant carcinoma Schneiderian
C2212276|Schneiderian carcinoma of prostate gland
C2212276|Schneiderian carcinoma of prostate gland (diagnosis)
C2212277|basaloid carcinoma of prostate gland
C2212277|basaloid carcinoma of prostate gland (diagnosis)
C2075845|cloacogenic carcinoma of prostate gland (diagnosis)
C2075845|cloacogenic carcinoma of prostate gland
C2033335|prostate malignant carcinoma transitional cell papillary
C2033335|papillary transitional cell carcinoma of prostate gland
C2033335|papillary transitional cell carcinoma of prostate gland (diagnosis)
C2212278|micropapillary transitional cell carcinoma of prostate gland (diagnosis)
C2212278|micropapillary transitional cell carcinoma of prostate gland
C2212279|adenoid cystic carcinoma of prostate gland
C2212279|adenoid cystic carcinoma of prostate gland (diagnosis)
C2138458|cribriform carcinoma of prostate gland (diagnosis)
C2138458|cribriform carcinoma of prostate gland
C2142686|prostate gland malignant carcinoma intracystic
C2142686|prostate gland malignant carcinoma intracystic (diagnosis)
C2212280|adenosquamous carcinoma of prostate gland
C2212280|adenosquamous carcinoma of prostate gland (diagnosis)
C2212281|epithelial-myoepithelial carcinoma of prostate gland
C2212281|epithelial-myoepithelial carcinoma of prostate gland (diagnosis)
C2212282|medullary carcinoma of prostate gland
C2212282|medullary carcinoma of prostate gland (diagnosis)
C2212283|scirrhous adenocarcinoma of prostate gland
C2212283|scirrhous adenocarcinoma of prostate gland (diagnosis)
C2212283|prostate gland malignant adenocarcinoma scirrhous
C2037349|superficial spreading adenocarcinoma of prostate (diagnosis)
C2037349|superficial spreading adenocarcinoma of prostate
C2033129|papillary adenocarcinoma of prostate gland
C2033129|papillary adenocarcinoma of prostate gland (diagnosis)
C2189645|villous adenocarcinoma of prostate gland
C2189645|villous adenocarcinoma of prostate gland (diagnosis)
C2212285|mucinous adenocarcinoma of prostate gland
C2212285|mucinous adenocarcinoma of prostate gland (diagnosis)
C2212286|mucin-producing adenocarcinoma of prostate gland
C2212286|mucin-producing adenocarcinoma of prostate gland (diagnosis)
C2018507|spindle cell sarcoma of prostate gland (diagnosis)
C2018507|spindle cell sarcoma of prostate gland
C2011321|giant cell sarcoma of prostate gland
C2011321|giant cell sarcoma of prostate gland (diagnosis)
C2212292|small cell sarcoma of prostate gland (diagnosis)
C2212292|small cell sarcoma of prostate gland
C2212293|epithelioid sarcoma of prostate gland (diagnosis)
C2212293|epithelioid sarcoma of prostate gland
C2188144|undifferentiated sarcoma of prostate gland (diagnosis)
C2188144|undifferentiated sarcoma of prostate gland
C2142687|desmoplastic small round cell tumor of prostate gland
C2142687|desmoplastic small round cell tumor of prostate gland (diagnosis)
C2170822|tubular adenocarcinoma of prostate gland
C2170822|tubular adenocarcinoma of prostate gland (diagnosis)
C2212295|fibromyxosarcoma of prostate gland
C2212295|fibromyxosarcoma of prostate gland (diagnosis)
C2212296|fascial fibrosarcoma of prostate gland (diagnosis)
C2212296|fascial fibrosarcoma of prostate gland
C2142682|infantile fibrosarcoma of prostate gland
C2142682|infantile fibrosarcoma of prostate gland (diagnosis)
C2142689|malignant solitary fibrous tumor of prostate gland (diagnosis)
C2142689|malignant solitary fibrous tumor of prostate gland
C2168295|leiomyosarcoma of prostate gland (diagnosis)
C2168295|leiomyosarcoma of prostate gland
C2168263|prostate gland neoplasm malignant leiomyosarcoma epithelioid
C2168263|epithelioid leiomyosarcoma of prostate gland (diagnosis)
C2168263|epithelioid leiomyosarcoma of prostate gland
C2212298|myxoid leiomyosarcoma of prostate gland (diagnosis)
C2212298|myxoid leiomyosarcoma of prostate gland
C1335518|rhabdomyosarcoma of prostate (diagnosis)
C1335518|prostate gland neoplasm malignant rhabdomyosarcoma
C1335518|rhabdomyosarcoma of prostate
C1335518|Prostate Rhabdomyosarcoma
C1335518|Rhabdomyosarcoma of the Prostate
C2212299|adult type pleomorphic rhabdomyosarcoma of prostate (diagnosis)
C2212299|prostate gland rhabdomyosarcoma pleomorphic, adult type
C2212299|adult type pleomorphic rhabdomyosarcoma of prostate
C1335508|prostate gland rhabdomyosarcoma embryonal
C1335508|embryonal rhabdomyosarcoma of prostate
C1335508|embryonal rhabdomyosarcoma of prostate (diagnosis)
C1335508|Embryonal Rhabdomyosarcoma of the Prostate
C1335508|Prostate Embryonal Rhabdomyosarcoma
C2018449|spindle cell rhabdomyosarcoma of prostate
C2018449|prostate gland rhabdomyosarcoma spindle cell
C2018449|spindle cell rhabdomyosarcoma of prostate (diagnosis)
C2212300|alveolar rhabdomyosarcoma of prostate (diagnosis)
C2212300|alveolar rhabdomyosarcoma of prostate
C2212300|prostate gland rhabdomyosarcoma alveolar
C2200364|rhabdomyosarcoma of prostate with ganglionic differentiation
C2200364|rhabdomyosarcoma of prostate with ganglionic differentiation (diagnosis)
C2200364|prostate rhabdomyosarcoma with ganglionic differentiation
C2212301|angiomyosarcoma of prostate gland (diagnosis)
C2212301|angiomyosarcoma of prostate gland
C2078063|intraductal papillary adenocarcinoma of prostate with invasion (diagnosis)
C2078063|intraductal papillary adenocarcinoma of prostate with invasion
C2212302|prostate gland rhabdomyosarcoma mixed type
C2212302|mixed type rhabdomyosarcoma of prostate
C2212302|mixed type rhabdomyosarcoma of prostate (diagnosis)
C2212303|embryonal carcinosarcoma of prostate gland (diagnosis)
C2212303|embryonal carcinosarcoma of prostate gland
C2212304|malignant myoepithelioma of prostate gland
C2212304|malignant myoepithelioma of prostate gland (diagnosis)
C2217396|malignant neoplasm of prostate TNM staging (diagnosis)
C2217396|malignant prostate neoplasm TNM staging
C2217396|malignant neoplasm of prostate TNM staging
C2217396|malignant prostatic neoplasm TNM staging
C2217396|prostatic cancer TNM staging
C2217396|malignant tumor of prostate TNM staging
C2217394|malignant neoplasm of prostate stage III
C2217394|malignant neoplasm of prostate stage III (diagnosis)
C2217394|malignant prostatic neoplasm stage III
C2217394|prostatic cancer stage III
C2217394|malignant tumor of prostate stage III
C2217408|malignant neoplasm of prostate TNM staging histiopathic grade (G) GX
C2217408|malignant neoplasm of prostate TNM staging histiopathic grade (G) GX (diagnosis)
C2217408|malignant prostatic neoplasm GX
C2217408|prostatic cancer TNM staging histiopathic grade (G) GX
C2217408|malignant tumor of prostate TNM staging histiopathic grade (G) GX
C2217405|malignant neoplasm of prostate TNM staging histiopathic grade (G) G1 (diagnosis)
C2217405|malignant neoplasm of prostate TNM staging histiopathic grade (G) G1
C2217405|malignant prostatic neoplasm G1
C2217405|prostatic cancer TNM staging histiopathic grade (G) G1
C2217405|malignant tumor of prostate TNM staging histiopathic grade (G) G1
C2217406|malignant neoplasm of prostate TNM staging histiopathic grade (G) G2 (diagnosis)
C2217406|malignant neoplasm of prostate TNM staging histiopathic grade (G) G2
C2217406|malignant prostatic neoplasm G2
C2217406|malignant tumor of prostate TNM staging histiopathic grade (G) G2
C2217406|prostatic cancer TNM staging histiopathic grade (G) G2
C2217407|malignant neoplasm of prostate TNM staging histiopathic grade (G) G3-4
C2217407|malignant neoplasm of prostate TNM staging histiopathic grade (G) G3-4 (diagnosis)
C2217407|malignant prostatic neoplasm G3-4
C2217407|prostatic cancer TNM staging histiopathic grade (G) G3-4
C2217407|malignant tumor of prostate TNM staging histiopathic grade (G) G3-4
C2217387|malignant neoplasm of prostate Jewett staging system
C2217387|malignant neoplasm of prostate Jewett staging system (diagnosis)
C2217387|malignant prostatic neoplasm Jewett staging system
C2217387|malignant tumor of prostate Jewett staging system
C2217387|prostatic cancer Jewett staging system
C2217388|malignant neoplasm of prostate Jewett staging system stage A (diagnosis)
C2217388|malignant neoplasm of prostate Jewett staging system stage A
C2217388|malignant prostatic neoplasm stage A
C2217388|prostatic cancer Jewett staging system stage A
C2217388|malignant tumor of prostate Jewett staging system stage A
C2217389|malignant neoplasm of prostate Jewett staging system stage B
C2217389|malignant neoplasm of prostate Jewett staging system stage B (diagnosis)
C2217389|malignant prostatic neoplasm stage B
C2217389|prostatic cancer Jewett staging system stage B
C2217389|malignant tumor of prostate Jewett staging system stage B
C2217390|malignant neoplasm of prostate Jewett staging system stage C
C2217390|malignant neoplasm of prostate Jewett staging system stage C (diagnosis)
C2217390|malignant prostatic neoplasm stage C
C2217390|malignant tumor of prostate Jewett staging system stage C
C2217390|prostatic cancer Jewett staging system stage C
C2217391|malignant neoplasm of prostate Jewett staging system stage D (diagnosis)
C2217391|malignant neoplasm of prostate Jewett staging system stage D
C2217391|malignant prostatic neoplasm stage D
C2217391|malignant tumor of prostate Jewett staging system stage D
C2217391|prostatic cancer Jewett staging system stage D
C3469524|prostate cancer susceptibility
C3469524|prostate cancer susceptibility (diagnosis)
C3469524|PROSTATE CANCER, SUSCEPTIBILITY TO
C1328504|Hormone refractory prostate cancer (disorder)
C1328504|Hormone refractory prostate cancer
C1328504|Hormone-refractory prostate cancer
C1328504|prostate gland malignant hormone refractory cancer
C1328504|Hormone refractory prostate cancer (diagnosis)
C1328504|HRPC
C3160891|Hormone-dependent prostate cancer
C1330959|primary malignant neoplasm of prostate (diagnosis)
C1330959|primary malignant neoplasm of prostate
C1330959|Primary malignant neoplasm of prostate (disorder)
C0347001|Metastatic Neoplasm to the Prostate
C0347001|Metastases to prostate
C0347001|secondary malignant neoplasm of prostate
C0347001|secondary malignant neoplasm of prostate (diagnosis)
C0347001|Metastatic Malignant Neoplasm to the Prostate Gland
C0347001|Metastatic Malignant Neoplasm in the Prostate Gland
C0347001|Cancer metastatic to prostate
C0347001|Metastasis to prostate
C0347001|Metastatic tumor to prostate
C0347001|Metastatic tumour to prostate
C0347001|Metastatic malignant neoplasm to prostate
C0347001|Secondary malignant neoplasm of prostate (disorder)
C0347001|Metastases to the Prostate
C0347001|Metastasis to the Prostate
C0347001|Metastatic Tumor to the Prostate
C1282482|local recurrence of malignant neoplasm of prostate
C1282482|local recurrence of malignant neoplasm of prostate (diagnosis)
C1282482|Local recurrence of malignant tumor of prostate (disorder)
C1282482|Local recurrence of malignant tumor of prostate
C1282482|Local recurrence of malignant tumour of prostate
C4030346|biopsy of prostate showed cribriform carcinoma (procedure)
C4030346|biopsy of prostate showed malignant carcinoma cribriform
C4030346|biopsy of prostate showed cribriform carcinoma
C4030340|biopsy of prostate showed giant cell and spindle cell carcinoma (procedure)
C4030340|biopsy of prostate showed giant cell and spindle cell carcinoma
C4030340|biopsy of prostate showed malignant carcinoma giant cell and spindle cell
C4030339|biopsy of prostate showed giant cell carcinoma
C4030339|biopsy of prostate showed malignant carcinoma giant cell
C4030339|biopsy of prostate showed giant cell carcinoma (procedure)
C4030286|biopsy of prostate showed malignant small cell type (procedure)
C4030286|biopsy of prostate showed malignant small cell type
C4030304|biopsy of prostate showed malignant fibrosarcoma solitary fibrous tumor (procedure)
C4030304|biopsy of prostate showed malignant fibrosarcoma solitary fibrous tumor
C4030342|biopsy of prostate showed malignant carcinoma epithelial-myoepithelial
C4030342|biopsy of prostate showed epithelial-myoepithelial carcinoma
C4030342|biopsy of prostate showed epithelial-myoepithelial carcinoma (procedure)
C4030293|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma mixed type
C4030293|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma mixed type (procedure)
C4030309|biopsy of prostate showed malignant clear cell type
C4030309|biopsy of prostate showed malignant clear cell type (procedure)
C4030355|biopsy of prostate showed basal cell adenocarcinoma
C4030355|biopsy of prostate showed malignant adenocarcinoma basal cell
C4030355|biopsy of prostate showed basal cell adenocarcinoma (procedure)
C4030300|biopsy of prostate showed malignant myosarcoma angiomyosarcoma (procedure)
C4030300|biopsy of prostate showed malignant myosarcoma angiomyosarcoma
C4030348|biopsy of prostate showed clear cell adenocarcinoma (procedure)
C4030348|biopsy of prostate showed clear cell adenocarcinoma
C4030348|biopsy of prostate showed malignant adenocarcinoma clear cell
C4030333|biopsy of prostate showed malignant adenocarcinoma in tubulovillous adenoma (procedure)
C4030333|biopsy of prostate showed malignant adenocarcinoma in tubulovillous adenoma
C4030297|biopsy of prostate showed malignant myosarcoma leiomyosarcoma myxoid
C4030297|biopsy of prostate showed malignant myosarcoma leiomyosarcoma myxoid (procedure)
C4030275|biopsy of prostate showed scirrhous adenocarcinoma (procedure)
C4030275|biopsy of prostate showed malignant adenocarcinoma scirrhous
C4030275|biopsy of prostate showed scirrhous adenocarcinoma
C4030325|biopsy of prostate showed malignant carcinoma small cell fusiform cell
C4030325|biopsy of prostate showed malignant carcinoma small cell fusiform cell (procedure)
C4030307|biopsy of prostate showed malignant fibrosarcoma fascial (procedure)
C4030307|biopsy of prostate showed malignant fibrosarcoma fascial
C4030305|biopsy of prostate showed malignant fibrosarcoma infantile
C4030305|biopsy of prostate showed malignant fibrosarcoma infantile (procedure)
C4030302|biopsy of prostate showed malignant marginal zone b-cell lymphoma
C4030302|biopsy of prostate showed malignant marginal zone b-cell lymphoma (procedure)
C4030368|biopsy of prostate showed acinar cell cystadenocarcinoma (procedure)
C4030368|biopsy of prostate showed acinar cell cystadenocarcinoma
C4030368|biopsy of prostate showed malignant carcinoma acinar cell cystadenocarcinoma
C4030295|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma alveolar (procedure)
C4030295|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma alveolar
C4030287|biopsy of prostate showed malignant sarcoma undifferentiated
C4030287|biopsy of prostate showed malignant sarcoma undifferentiated (procedure)
C4030283|biopsy of prostate showed malignant adenocarcinoma mucinous
C4030283|biopsy of prostate showed mucinous adenocarcinoma
C4030283|biopsy of prostate showed mucinous adenocarcinoma (procedure)
C4030330|biopsy of prostate showed malignant carcinoma large cell with rhabdoid phenotype
C4030330|biopsy of prostate showed malignant carcinoma large cell with rhabdoid phenotype (procedure)
C4030288|biopsy of prostate showed malignant sarcoma small cell (procedure)
C4030288|biopsy of prostate showed malignant sarcoma small cell
C4030285|biopsy of prostate showed malignant spindle cell type (procedure)
C4030285|biopsy of prostate showed malignant spindle cell type
C4030277|biopsy of prostate showed pleomorphic carcinoma (procedure)
C4030277|biopsy of prostate showed malignant carcinoma pleomorphic
C4030277|biopsy of prostate showed pleomorphic carcinoma
C4030322|biopsy of prostate showed malignant carcinoma squamous cell large cell, nonkerat (procedure)
C4030322|biopsy of prostate showed malignant carcinoma squamous cell large cell, nonkerat
C4030312|biopsy of prostate showed malignant carcinosarcoma (procedure)
C4030312|biopsy of prostate showed malignant carcinosarcoma
C4030334|biopsy of prostate showed malignant carcinoma large cell neuroendocrine
C4030334|biopsy of prostate showed large cell neuroendocrine carcinoma (procedure)
C4030334|biopsy of prostate showed large cell neuroendocrine carcinoma
C4030298|biopsy of prostate showed malignant myosarcoma leiomyosarcoma epithelioid (procedure)
C4030298|biopsy of prostate showed malignant myosarcoma leiomyosarcoma epithelioid
C4030294|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma embryonal
C4030294|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma embryonal (procedure)
C4030271|biopsy of prostate showed superficial spreading adenocarcinoma
C4030271|biopsy of prostate showed malignant adenocarcinoma superficial spreading
C4030271|biopsy of prostate showed superficial spreading adenocarcinoma (procedure)
C4030267|biopsy of prostate showed villous adenocarcinoma (procedure)
C4030267|biopsy of prostate showed villous adenocarcinoma
C4030267|biopsy of prostate showed malignant adenocarcinoma villous
C4030323|biopsy of prostate showed malignant carcinoma squamous cell keratinizing
C4030323|biopsy of prostate showed malignant carcinoma squamous cell keratinizing (procedure)
C4030308|biopsy of prostate showed malignant fibrosarcoma (procedure)
C4030308|biopsy of prostate showed malignant fibrosarcoma
C4030363|biopsy of prostate showed adenocarcinoma with metaplasia (procedure)
C4030363|biopsy of prostate showed adenocarcinoma with metaplasia
C4030363|biopsy of prostate showed malignant adenocarcinoma with metaplasia
C4030344|biopsy of prostate showed duct carcinoma, desmoplastic type (procedure)
C4030344|biopsy of prostate showed duct carcinoma, desmoplastic type
C4030344|biopsy of prostate showed malignant carcinoma duct, desmoplastic type
C4030296|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma
C4030296|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma (procedure)
C4030278|biopsy of prostate showed malignant carcinoma papillary
C4030278|biopsy of prostate showed papillary carcinoma (procedure)
C4030278|biopsy of prostate showed papillary carcinoma
C4030269|biopsy of prostate showed tubular adenocarcinoma
C4030269|biopsy of prostate showed tubular adenocarcinoma (procedure)
C4030269|biopsy of prostate showed malignant adenocarcinoma tubular
C4030328|biopsy of prostate showed malignant carcinoma pseudosarcomatous
C4030328|biopsy of prostate showed malignant carcinoma pseudosarcomatous (procedure)
C4030318|biopsy of prostate showed malignant carcinoma squamous cell with horn formation
C4030318|biopsy of prostate showed malignant carcinoma squamous cell with horn formation (procedure)
C4030303|biopsy of prostate showed malignant giant cell type
C4030303|biopsy of prostate showed malignant giant cell type (procedure)
C4030356|biopsy of prostate showed anaplastic carcinoma (procedure)
C4030356|biopsy of prostate showed malignant carcinoma anaplastic
C4030356|biopsy of prostate showed anaplastic carcinoma
C4030331|biopsy of prostate showed malignant carcinoma epithelioma
C4030331|biopsy of prostate showed malignant carcinoma epithelioma (procedure)
C4030281|biopsy of prostate showed myosarcoma rhabdomyosarcoma pleomorphic, adult type
C4030281|biopsy of prostate showed myosarcoma rhabdomyosarcoma pleomorphic, adult type (procedure)
C4030279|biopsy of prostate showed malignant adenocarcinoma papillary
C4030279|biopsy of prostate showed papillary adenocarcinoma
C4030279|biopsy of prostate showed papillary adenocarcinoma (procedure)
C4030268|biopsy of prostate showed malignant carcinoma verrucous
C4030268|biopsy of prostate showed verrucous carcinoma
C4030268|biopsy of prostate showed verrucous carcinoma (procedure)
C4030301|biopsy of prostate showed malignant myosarcoma
C4030301|biopsy of prostate showed malignant myosarcoma (procedure)
C4030299|biopsy of prostate showed malignant myosarcoma leiomyosarcoma
C4030299|biopsy of prostate showed malignant myosarcoma leiomyosarcoma (procedure)
C4030292|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma spindle cell
C4030292|biopsy of prostate showed malignant myosarcoma rhabdomyosarcoma spindle cell (procedure)
C4030291|biopsy of prostate showed a malignant neoplasm
C4030291|biopsy of prostate showed malignant neoplasm (procedure)
C4030291|biopsy of prostate showed malignant neoplasm
C4030290|biopsy of prostate showed malignant sarcoma (procedure)
C4030290|biopsy of prostate showed malignant sarcoma
C4030273|biopsy of prostate showed spindle cell sarcoma
C4030273|biopsy of prostate showed spindle cell sarcoma (procedure)
C4030273|biopsy of prostate showed malignant sarcoma spindle cell
C4030324|biopsy of prostate showed malignant carcinoma squamous cell adenoid
C4030324|biopsy of prostate showed malignant carcinoma squamous cell adenoid (procedure)
C4030317|biopsy of prostate showed malignant carcinoma transitional cell micropapillary (procedure)
C4030317|biopsy of prostate showed malignant carcinoma transitional cell micropapillary
C4030338|biopsy of prostate showed malignant carcinoma glassy cell
C4030338|biopsy of prostate showed glassy cell carcinoma
C4030338|biopsy of prostate showed glassy cell carcinoma (procedure)
C4030276|biopsy of prostate showed polygonal cell carcinoma
C4030276|biopsy of prostate showed malignant carcinoma polygonal cell
C4030276|biopsy of prostate showed polygonal cell carcinoma (procedure)
C4030274|biopsy of prostate showed malignant carcinoma spindle cell
C4030274|biopsy of prostate showed spindle cell carcinoma
C4030274|biopsy of prostate showed spindle cell carcinoma (procedure)
C4030321|biopsy of prostate showed malignant carcinoma squamous cell microinvasive
C4030321|biopsy of prostate showed malignant carcinoma squamous cell microinvasive (procedure)
C4030313|biopsy of prostate showed malignant carcinoma with osteoclast-like cells (procedure)
C4030313|biopsy of prostate showed malignant carcinoma with osteoclast-like cells
C4030280|biopsy of prostate showed myosarcoma rhabdomyosarcoma with ganglionic differentiation
C4030280|biopsy of prostate showed myosarcoma rhabdomyosarcoma with ganglionic differentiation (procedure)
C4030289|biopsy of prostate showed malignant sarcoma giant cell (procedure)
C4030289|biopsy of prostate showed malignant sarcoma giant cell
C4030327|biopsy of prostate showed malignant carcinoma schneiderian (procedure)
C4030327|biopsy of prostate showed malignant carcinoma schneiderian
C4030311|biopsy of prostate showed malignant carcinosarcoma embryonal type
C4030311|biopsy of prostate showed malignant carcinosarcoma embryonal type (procedure)
C4030310|biopsy of prostate showed malignant carcinosarcoma myoepithelioma (procedure)
C4030310|biopsy of prostate showed malignant carcinosarcoma myoepithelioma
C4030345|biopsy of prostate showed desmoplastic small round cell sarcoma (procedure)
C4030345|biopsy of prostate showed desmoplastic small round cell sarcoma
C4030345|biopsy of prostate showed malignant sarcoma desmoplastic small round cell
C4030272|biopsy of prostate showed malignant carcinoma squamous cell
C4030272|biopsy of prostate showed squamous cell carcinoma
C4030272|biopsy of prostate showed squamous cell carcinoma (procedure)
C4030270|biopsy of prostate showed malignant carcinoma transitional cell
C4030270|biopsy of prostate showed transitional cell carcinoma (procedure)
C4030270|biopsy of prostate showed transitional cell carcinoma
C4030316|biopsy of prostate showed malignant carcinoma transitional cell papillary
C4030316|biopsy of prostate showed malignant carcinoma transitional cell papillary (procedure)
C4030358|biopsy of prostate showed malignant carcinoma adenosquamous
C4030358|biopsy of prostate showed adenosquamous carcinoma
C4030358|biopsy of prostate showed adenosquamous carcinoma (procedure)
C4030357|biopsy of prostate showed malignant adenocarcinoma alveolar
C4030357|biopsy of prostate showed alveolar adenocarcinoma (procedure)
C4030357|biopsy of prostate showed alveolar adenocarcinoma
C4030341|biopsy of prostate showed malignant sarcoma epithelioid
C4030341|biopsy of prostate showed epithelioid sarcoma (procedure)
C4030341|biopsy of prostate showed epithelioid sarcoma
C4030332|biopsy of prostate showed malignant adenocarcinoma in villous adenoma (procedure)
C4030332|biopsy of prostate showed malignant adenocarcinoma in villous adenoma
C4030319|biopsy of prostate showed malignant carcinoma squamous cell spindle cell (procedure)
C4030319|biopsy of prostate showed malignant carcinoma squamous cell spindle cell
C4030314|biopsy of prostate showed malignant carcinoma undifferentiated
C4030314|biopsy of prostate showed malignant carcinoma undifferentiated (procedure)
C4030359|biopsy of prostate showed malignant carcinoma adenoid cystic
C4030359|biopsy of prostate showed adenoid cystic carcinoma (procedure)
C4030359|biopsy of prostate showed adenoid cystic carcinoma
C4030354|biopsy of prostate showed malignant carcinoma basaloid
C4030354|biopsy of prostate showed basaloid carcinoma (procedure)
C4030354|biopsy of prostate showed basaloid carcinoma
C4030335|biopsy of prostate showed large cell carcinoma
C4030335|biopsy of prostate showed malignant carcinoma large cell
C4030335|biopsy of prostate showed large cell carcinoma (procedure)
C4030366|biopsy of prostate showed adenocarcinoma intraductal papillary, with invasion
C4030366|biopsy of prostate showed adenocarcinoma intraductal papillary, with invasion (procedure)
C4030284|biopsy of prostate showed medullary carcinoma
C4030284|biopsy of prostate showed malignant carcinoma medullary
C4030284|biopsy of prostate showed medullary carcinoma (procedure)
C4030282|biopsy of prostate showed malignant adenocarcinoma mucin-producing
C4030282|biopsy of prostate showed mucin-producing adenocarcinoma
C4030282|biopsy of prostate showed mucin-producing adenocarcinoma (procedure)
C4030369|biopsy of prostate showed acinar cell carcinoma
C4030369|biopsy of prostate showed malignant carcinoma acinar cell
C4030369|biopsy of prostate showed acinar cell carcinoma (procedure)
C4030347|biopsy of prostate showed malignant carcinoma cloacogenic
C4030347|biopsy of prostate showed cloacogenic carcinoma
C4030347|biopsy of prostate showed cloacogenic carcinoma (procedure)
C4030329|biopsy of prostate showed malignant carcinoma papillary squamous cell (procedure)
C4030329|biopsy of prostate showed malignant carcinoma papillary squamous cell
C4030320|biopsy of prostate showed malignant carcinoma squamous cell small cell, nonkerat (procedure)
C4030320|biopsy of prostate showed malignant carcinoma squamous cell small cell, nonkerat
C4030315|biopsy of prostate showed malignant carcinoma transitional cell spindle cell
C4030315|biopsy of prostate showed malignant carcinoma transitional cell spindle cell (procedure)
C4030306|biopsy of prostate showed malignant fibrosarcoma fibromyxosarcoma
C4030306|biopsy of prostate showed malignant fibrosarcoma fibromyxosarcoma (procedure)
C1282496|metastasis from malignant neoplasm of prostate (diagnosis)
C1282496|metastasis from malignant neoplasm of prostate
C1282496|Cancer of the prostate with metastasis
C1282496|Metastatic prostate cancer
C1282496|Metastasis from malignant tumor of prostate
C1282496|Metastasis from malignant tumor of prostate (disorder)
C1282496|Metastasis from malignant tumour of prostate
C4081803|Prostate cancer metastatic to eye (disorder)
C4081803|Prostate cancer metastatic to eye
C1302530|squamous cell carcinoma of prostate gland
C1302530|squamous cell carcinoma of prostate gland (diagnosis)
C1302530|Squamous cell carcinoma of prostate (disorder)
C1302530|Squamous cell carcinoma of prostate
C1302530|Prostate Squamous Cell Carcinoma
C1302530|Squamous Cell Carcinoma of the Prostate
C0154088|Prostate
C0154088|Carcinoma in situ of prostate
C0154088|carcinoma in situ of prostate gland (diagnosis)
C0154088|carcinoma in situ of prostate gland
C0154088|Ca in situ prostate
C0154088|CIS - Carcinoma in situ of prostate
C0154088|Cancer in situ of prostate
C0154088|CIS (Carcinoma in situ) of prostate
C0154088|Carcinoma in situ of prostate (disorder)
C0154088|PIN III
C0154088|Prostatic intraepithelial neoplasia, grade III
C0154088|Adenocarcinoma in situ of Prostate
C0154088|Adenocarcinoma in situ of the Prostate
C0154088|Grade 3 PIN
C0154088|Grade 3 Prostatic Intraepithelial Neoplasia
C0154088|Grade III PIN
C0154088|Grade III Prostatic Intraepithelial Neoplasia
C0154088|Prostate Adenocarcinoma in situ
C1386259|endometrioid; adenocarcinoma, unspecified site, male
C1386259|adenocarcinoma; endometrioid, unspecified site, male
C1391907|carcinoma; endometrioid, unspecified site, male
C1391907|endometrioid; carcinoma, unspecified site, male
C1394298|cystadenocarcinoma; endometrioid, unspecified site, male
C1394298|endometrioid; cystadenocarcinoma, unspecified site, male
C0279882|cellular diagnosis, prostate cancer
C0279882|prostate cancer cellular diagnosis
C0280280|stage, prostate cancer
C0280280|prostate cancer stage
C1335514|Extramedullary Myeloid Neoplasm of Prostate
C1335514|Extramedullary Myeloid Neoplasm of the Prostate
C1335514|Extramedullary Myeloid Tumor of Prostate
C1335514|Extramedullary Myeloid Tumor of the Prostate
C1335514|Prostate Extramedullary Myeloid Neoplasm
C1335514|Prostate Extramedullary Myeloid Tumor
C1335514|Prostate Myeloid Sarcoma
C1335514|Prostatic Chloroma
C1335514|Prostatic Extramedullary Myeloid Neoplasm
C1335514|Prostatic Extramedullary Myeloid Tumor
C1335514|Prostatic Myeloid Sarcoma
C0238393|Prostate Sarcoma
C0238393|Sarcoma of Prostate
C0238393|Sarcoma of the Prostate
C1334615|Malignant Phyllodes Tumor of Prostate
C1334615|Phyllodes Tumor of the Prostate
C1334615|Malignant Phyllodes Neoplasm of Prostate
C1334615|Malignant Phyllodes Neoplasm of the Prostate
C1334615|Malignant Phyllodes Tumor of the Prostate
C1334615|Malignant Prostate Phyllodes Neoplasm
C1334615|Malignant Prostate Phyllodes Tumor
C1335512|Primary Prostate Lymphoma
C1335512|Lymphoma of Prostate
C1335512|Lymphoma of the Prostate
C1335512|Prostate Lymphoma
C1276489|T3a: Prostate tumor with extracapsular extension (unilateral or bilateral) (finding)
C1276489|T3a: Prostate tumor with extracapsular extension (unilateral or bilateral)
C1276489|T3a: Prostate tumour with extracapsular extension (unilateral or bilateral)
C1276489|T3a: Prostate tumor with extracapsular extension (unilateral or bilateral) (tumor staging)
C1720586|Extraprostatic extension of tumor present, non-focal (finding)
C1720586|Extraprostatic extension of tumor present, non-focal
C1720586|Extraprostatic extension of tumour present, non-focal
C1300585|small cell carcinoma of prostate gland (diagnosis)
C1300585|small cell carcinoma of prostate gland
C1300585|Prostate Small Cell NEC
C1300585|Prostate Small Cell Neuroendocrine Carcinoma
C1300585|Oat Cell Carcinoma of Prostate
C1300585|Small cell carcinoma of prostate (disorder)
C1300585|Small cell carcinoma of prostate
C1300585|Oat Cell Carcinoma of the Prostate
C1300585|Prostate Oat Cell Carcinoma
C1300585|Prostate Small Cell Carcinoma
C1300585|Small Cell Carcinoma of the Prostate
C1276487|T2a: Prostate tumor involves one lobe (finding)
C1276487|T2a: Prostate tumor involves one lobe
C1276487|T2a: Prostate tumour involves one lobe
C1276487|T2a: Prostate tumor involves one lobe (tumor staging)
C0349672|Endometrioid carcinoma of prostate
C0349672|prostate gland malignant carcinoma endometrioid
C0349672|Endometrioid carcinoma of prostate (diagnosis)
C0349672|Endometrioid carcinoma of prostate (disorder)
C0349672|Ductal Adenocarcinoma of Prostate
C0349672|Ductal Adenocarcinoma of the Prostate
C0349672|Endometrioid Adenocarcinoma of Prostate
C0349672|Endometrioid Adenocarcinoma of the Prostate
C0349672|Endometrioid Carcinoma of the Prostate
C0349672|Prostate Ductal Adenocarcinoma
C0349672|Prostate Endometrioid Adenocarcinoma
C0349672|Prostate Endometrioid Carcinoma
C0349672|Prostatic Endometrioid Carcinoma
C1276488|T3: Prostate tumor extends through the prostatic capsule (finding)
C1276488|T3: Prostate tumor extends through the prostatic capsule
C1276488|T3: Prostate tumour extends through the prostatic capsule
C1276488|T3: Prostate tumor extends through the prostatic capsule (tumor staging)
C1276626|T2: Tumor confined within the prostate (finding)
C1276626|T2: Tumor confined within the prostate
C1276626|T2: Tumour confined within the prostate
C1276626|T2: Tumor confined within the prostate (tumor staging)
C0392920|Cancer chemotherapy
C0392920|Chemotherapy Regimen
C0392920|chemotherapeutics regimen
C0392920|chemotherapeutics regimen (treatment)
C0392920|neoplasm/cancer chemotherapy
C0392920|neoplasm chemotherapy
C0392920|Chemotherapy
C0392920|Cancer chemotherapy (regime/therapy)
C0392920|Chemotherapy (procedure)
C0392920|Cancer chemotherapy regimen
C0392920|Antineoplastic chemotherapy regimen (procedure)
C0392920|Antineoplastic chemotherapy regimen
C0392920|neoplasm/cancer pharmacotherapy
C0392920|neoplasm pharmacotherapy
C0392920|cancer pharmacotherapy
C0392920|cancer; chemotherapy
C0392920|chemotherapy; cancer
C0392920|chemotherapy; neoplasm
C0392920|neoplasm; chemotherapy
C0392920|Chemotherapy, NOS
C0392920|Antineoplastic chemotherapy regimen (regime/therapy)
C0280024|mercaptopurine/methotrexate/prednisolone/vincristine
C0280024|POMP
C0280024|MP/MTX/PRDL/VCR
C0280024|mercaptopurine/methotrexate/prednisolone/vincristine protocol
C0280075|mercaptopurine/methotrexate/methylprednisolone/vincristine
C0280075|POMP
C0280075|MePRDL/MP/MTX/VCR
C0280075|mercaptopurine/methotrexate/methylprednisolone/vincristine protocol
C0280580|doxorubicin/fluorouracil
C0280580|AFA
C0280580|FA
C0280580|DOX/5-FU
C0280580|doxorubicin/fluorouracil protocol
C0280593|doxorubicin/fluorouracil/semustine
C0280593|MEFA
C0280593|FAME
C0280593|DOX/5-FU/MeCCNU
C0280593|doxorubicin/fluorouracil/semustine protocol
C0338272|CL
C0338272|cyclophosphamide/losoxantrone
C0338272|CTX/DuP-941
C2045825|chemotherapeutics regimen first line of treatment
C2045825|chemotherapeutics regimen first line of treatment (treatment)
C2045828|chemotherapeutics regimen second line of treatment
C2045828|chemotherapeutics regimen second line of treatment (treatment)
C2045827|oral chemotherapeutics regimen
C2045827|oral chemotherapeutics regimen (treatment)
C2045826|intravenous chemotherapeutics regimen
C2045826|intravenous chemotherapeutics regimen (treatment)
C3179010|Induction Chemotherapy
C3179010|Chemotherapy, Induction
C3179010|Chemotherapies, Induction
C3179010|Induction Chemotherapies
C3179010|Induction chemotherapy (procedure)
C0374470|CHEMO INTRALESIONAL OVER 7
C0374470|intralesional chemotherapy administration for more than 7 lesions
C0374470|intralesional chemotherapy administration for more than 7 lesions (treatment)
C0374470|CHEMOTHERAPY ADMINISTRATION INTRALESIONAL >7
C0374470|Chemotherapy administration; intralesional, more than 7 lesions
C0199953|Chemotherapy administration, intra-arterial; push technique
C0199953|chemotherapy by intra-arterial push technique
C0199953|chemotherapy by intra-arterial push technique (treatment)
C0199953|CHEMO IA PUSH TECNIQUE
C0199953|CHEMOTHERAPY ADMIN INTRA-ARTERIAL PUSH TQ
C0199953|Intra-arterial, push technique chemotherapy administration
C0199953|Injection of chemotherapy using push technique into an artery
C0199953|Retired procedure (procedure) [P2-67050]
C0199953|Retired procedure [P2-67050]
C0580690|TB chemotherapy (procedure)
C0580690|Tuberculosis chemotherapy (procedure)
C0580690|Tuberculosis chemotherapy
C0580690|TB chemotherapy
C0580690|TB chemotherapy (regime/therapy)
C1302181|chemotherapeutics regimen cycle (treatment)
C1302181|chemotherapeutics regimen cycle
C1302181|Chemotherapy cycle
C1302181|Chemotherapy cycle (procedure)
C1302181|Chemotherapy cycle (regime/therapy)
C0413365|Intravenous chemotherapy
C0413365|Intravenous drug therapy
C0413365|Intravenous chemotherapy (procedure)
C0413365|Intravenous therapy: [chemo-] or [drug] (procedure)
C0413365|Intravenous therapy: [chemo-] or [drug]
C0413365|Intravenous chemotherapy (treatment)
C0260835|Chemotherapy follow-up (procedure)
C0260835|Chemotherapy follow-up
C0260835|Chemotherapy follow-up (regime/therapy)
C0199957|Chemotherapy administration, subcutaneous, with local anesthesia
C0199957|Chemotherapy administration, subcutaneous, with local anaesthesia
C0199957|Chemotherapy administration, subcutaneous, with local anesthesia (procedure)
C0199957|Chemotherapy administration, subcutaneous, with local anesthesia (regime/therapy)
C0198526|Chemotherapy administration into peritoneal cavity requiring paracentesis
C0198526|Chemotherapy administration into peritoneal cavity requiring paracentesis (procedure)
C0198526|Chemotherapy administration into peritoneal cavity requiring paracentesis (regime/therapy)
C0189560|Chemotherapy administration into pleural cavity, requiring and including thoracentesis
C0189560|Chemotherapy administration into pleural cavity requiring thoracentesis (procedure)
C0189560|CHEMOTHERAPY INTRACAVITARY
C0189560|Chemotherapy administration into pleural cavity with thoracentesis
C0189560|Chemotherapy administration into pleural cavity requiring thoracentesis
C0189560|Chemotherapy administration into pleural cavity requiring thoracentesis (regime/therapy)
C0189560|CHEMOTX ADMN PLEURAL CAVITY REQ&W/THORACNTS
C0419073|Oral cytotoxic drug therapy
C0419073|Oral chemotherapy
C0419073|Oral chemotherapy (procedure)
C0419073|Oral chemotherapy (regime/therapy)
C0199948|Chemotherapy for non-neoplastic disease
C0199948|Chemotherapy for non-neoplastic disease (procedure)
C0199948|Chemotherapy for non-neoplastic disease, NOS
C0199948|Chemotherapy for non-neoplastic disease (regime/therapy)
C0282515|Chemoprevention
C0282515|CHEMOPREV
C0282515|Prescription of a prophylactic chemotherapeutic agent
C0282515|Prescription of a prophylactic chemotherapeutic agent (procedure)
C0282515|Prophylactic chemotherapy
C0282515|Chemoprophylaxis
C0282515|Prophylactic chemotherapy (procedure)
C0282515|Prophylactic chemotherapy NOS
C0282515|Prophylactic chemotherapy NOS (procedure)
C0282515|chemotherapy prophylactic
C0282515|prophylactic chemotherapy (treatment)
C0282515|Chemoprophylaxis NOS
C0282515|Prescription of a prophylactic chemotherapeutic agent, NOS
C0282515|Prophylactic chemotherapy (regime/therapy)
C0282515|Prophylactic chemotherapy NOS (regime/therapy)
C1276154|Ambulatory chemotherapy (procedure)
C1276154|Ambulatory chemotherapy
C1276154|ambulatory chemotherapy administration (medication)
C1276154|chemotherapy administration ambulatory
C1276154|ambulatory chemotherapy administration
C1276154|Ambulatory chemotherapy (regime/therapy)
C3695058|chemotherapeutics regimen intracavitary (treatment)
C3695058|chemotherapeutics regimen intracavitary
C3665477|Chemotherapy Regimen or Agent Combination
C3665477|Combination Chemotherapy Regimen
C0476658|Chemotherapy session for neoplasm
C0476658|[V]Chemotherapy session for neoplasm (context-dependent category)
C0476658|Encounter for antineoplastic chemotherapy and immunotherapy
C0476658|[V]Chemotherapy session for neoplasm
C0476658|[V]Chemotherapy session for neoplasm (situation)
C0476658|Encounter due to Chemotherapy session for neoplasm
C0476658|Encounter or admission for chemotherapy
C0178200|Inject ca chemother NEC
C0178200|Injection or infusion of cancer chemotherapeutic substance
C0178200|Injection or infusion of antineoplastic agent
C0374469|intralesional chemotherapy administration up to and including 7 lesions
C0374469|intralesional chemotherapy administration up to and including 7 lesions (treatment)
C0374469|CHEMO INTRALESIONAL UP TO 7
C0374469|CHEMOTHERAPY ADMINISTRATION INTRALESIONAL </7
C0374469|Chemotherapy administration; intralesional, up to and including 7 lesions
C0374473|CHEMOTHERAPY INTO CNS
C0374473|CHEMOTX ADMN CNS REQ SPINAL PUNCTURE
C0374473|Chemotherapy administration, into CNS (eg, intrathecal), requiring and including spinal puncture
C0199944|oral chemotherapeutics regimen for malignant neoplasm (treatment)
C0199944|oral chemotherapeutics regimen for malignant neoplasm
C0199944|chemotherapeutics regimen oral for malignant neoplasm
C0199944|Oral chemotherapy for malignant neoplasm
C0199944|Oral chemotherapy for malignant neoplasm (procedure)
C0199944|Oral chemotherapy for malignant neoplasm (regime/therapy)
C0278925|Chemoprevention of Cancer
C0278925|Cancer Chemoprevention
C0278925|chemoprevention
C0279023|potentiation
C0279023|chemosensitization/potentiation
C0279023|potentiation/chemosensitization
C0279023|Chemosensitization
C0281488|In Vitro Sensitivity-Directed Chemotherapy
C0199946|topical chemotherapy for malignant neoplasm (treatment)
C0199946|Topical chemotherapy for malignant neoplasm
C0199946|Topical chemotherapy for malignant neoplasm (procedure)
C0199946|Topical chemotherapy for malignant neoplasm (regime/therapy)
C0189561|Pleurodesis with cancer chemotherapy substance
C0189561|Pleurodesis with cancer chemotherapy substance (procedure)
C0199942|Perfusion chemotherapy for malignant neoplasm
C0199942|perfusion chemotherapy for malignant neoplasm (treatment)
C0199942|Perfusion chemotherapy for malignant neoplasm (procedure)
C0199942|Perfusion chemotherapy for malignant neoplasm (regime/therapy)
C0199940|Parenteral chemotherapy for malignant neoplasm
C0199940|parenteral chemotherapy for malignant neoplasm (treatment)
C0199940|Parenteral chemotherapy for malignant neoplasm (procedure)
C0199940|Parenteral chemotherapy for malignant neoplasm (regime/therapy)
C0199943|chemotherapeutics regimen intracavitary for malignant neoplasm
C0199943|intracavitary chemotherapeutics regimen for malignant neoplasm (treatment)
C0199943|intracavitary chemotherapeutics regimen for malignant neoplasm
C0199943|Intracavitary chemotherapy for malignant neoplasm
C0199943|Intracavitary chemotherapy for malignant neoplasm (procedure)
C0199943|Intracavitary chemotherapy for malignant neoplasm (regime/therapy)
C0199941|intravenous chemotherapy for malignant neoplasm (treatment)
C0199941|intravenous chemotherapy for malignant neoplasm
C0199941|chemotherapy intravenous for malignant neoplasm
C0199941|Infusion chemotherapy for malignant neoplasm
C0199941|Infusion chemotherapy for malignant neoplasm (procedure)
C0199941|Infusion chemotherapy for malignant neoplasm (regime/therapy)
C0191103|Intravenous, push technique chemotherapy administration
C0191103|Intravenous chemotherapy administration by push technique
C0191103|Intravenous chemotherapy administration by push technique (procedure)
C0199945|local chemotherapy for malignant neoplasm (treatment)
C0199945|Local chemotherapy for malignant neoplasm
C0199945|Local chemotherapy for malignant neoplasm (procedure)
C0199945|Local chemotherapy for malignant neoplasm (regime/therapy)
C0436299|Radiomimetic chemotherapy (procedure)
C0436299|Radiomimetic chemotherapy
C0436299|radiomimetic chemotherapy (treatment)
C0436299|Radiomimetic chemotherapy (regime/therapy)
C0199947|Chemotherapy for non-malignant neoplasm
C0199947|Chemotherapy for non-malignant neoplasm (procedure)
C0199947|Chemotherapy for non-malignant neoplasm, NOS
C0199947|Chemotherapy for non-malignant neoplasm (regime/therapy)
C0279512|cytarabine/daunorubicin/prednisone/thioguanine
C0279512|TRAP
C0279512|ARA-C/DNR/PRED/TG
C1521869|CTX/IFF/VP-16
C1521869|Ifosfamide/Cyclophosphamide/Etoposide
C1327770|CCI-779/IFN-A
C1327770|interferon alfa/temsirolimus
C1327770|CCI-779/Interferon Alfa
C1327912|galiximab/rituximab
C1327912|IDEC-114 Monoclonal Antibody/Rituximab
C1327912|MOAB IDEC-114/MOAB IDEC-C2B8
C1327970|letrozole/temsirolimus
C1327970|CCI-779/LTZ
C1327970|CCI-779/Letrozole
C1328116|captopril/recombinant tissue plasminogen activator
C1328116|Captopril/Tissue Plasminogen Activator
C1328116|CPT/t-PA
C0935858|ARA-C/ASP/DNR/MTX/PRDL/VCR
C0935858|asparaginase/cytarabine/daunorubicin/methotrexate/prednisolone/vincristine
C1134539|APC8015 vaccine/bevacizumab
C1134539|APC8015/Bevacizumab
C1134539|APC 8015/MOAB VEGF
C1134602|fowlpox virus vaccine vector/gp100 antigen/interleukin-2
C1134602|Fowlpox Virus Vaccine/gp100 Antigen/Interleukin-2
C1134602|FOWLVAC/gp100/IL-2
C0278888|interleukin-2/recombinant interferon beta
C0278888|IFN-B/IL-2
C0278888|Interferon Beta/Interleukin-2
C0278889|interferon gamma/recombinant interferon beta
C0278889|IFN-B/IFN-G
C0278889|Interferon Beta/Interferon Gamma
C0279257|recombinant interferon beta/zidovudine
C0279257|IFN-B/ZDV
C0279257|Interferon Beta/Zidovudine
C0279438|fluorouracil/recombinant interferon beta
C0279438|5-FU/IFN-B
C0279438|Fluorouracil/Interferon Beta
C0281419|isotretinoin/recombinant interferon beta
C0281419|13-CRA/IFN-B
C0281419|Interferon Beta/Isotretinoin
C0281420|Beta CT/VIT-A
C0281420|beta carotene/vitamin A regimen
C0281420|beta carotene/vitamin A
C0281420|beta carotene/VIT-A
C0281711|cisplatin/dihydrosphingosine
C0281711|CDDP/safingol
C0281711|Cisplatin/Safingol
C0393027|Ethynyluracil/Fluorouracil
C0393027|Eniluracil / 5-FU Combination Tablet
C0393027|GW776/5-FU
C0393027|GW776/5-Fluorouracil
C0393027|776C85/5-FU
C0393027|Eniluracil/Fluorouracil
C0393028|ethynyluracil/fluorouracil/leucovorin calcium
C0393028|776C85/CF/5-FU
C0393028|Eniluracil/Fluorouracil/Leucovorin Calcium
C0796602|fowlpox virus vaccine vector/interleukin-2
C0796602|FOWLVAC/IL-2
C0796602|Fowlpox Virus Vaccine/Interleukin-2
C0796658|fowlpox virus vaccine vector/interleukin-2/vaccinia-tyrosinase vaccine
C0796658|Fowlpox Virus Vaccine/Interleukin-2/Vaccinia-Tyrosinase Vaccine
C0796658|FOWLVAC/IL-2/VACTYROS
C0879332|HER-2/neu peptide vaccine/Montanide ISA-51
C0879332|HER-2-neu peptide vaccine/Montanide ISA-51
C0879332|HER-2/ISA-51
C0879358|HER-2/neu peptide vaccine/sargramostim
C0879358|HER-2-Neu Peptide Vaccine/Sargramostim
C0879358|GM-CSF/HER-2
C1831695|CTX/DOX/MOAB VEGF/TXT
C1831695|bevacizumab/cyclophosphamide/docetaxel/doxorubicin
C1831713|cisplatin/doxorubicin/etoposide/ifosfamide/methotrexate
C1831713|CDDP/DOX/IFF/MTX/VP-16
C1880034|Chemotherapy Regimen Used to Treat Malignant Brain Neoplasm
C1880033|Chemotherapy Regimen Used to Treat Acute Myeloid Leukemia
C1880060|Chemotherapy Regimen Used to Treat Plasma Cell Myeloma
C1880065|Chemotherapy Regimen Used to Treat Small Cell Lung Carcinoma
C1880051|Chemotherapy Regimen Used to Treat Malignant Mesothelioma
C1880043|Chemotherapy Regimen Used to Treat Chronic Lymphocytic Leukemia
C1880064|Chemotherapy Regimen Used to Treat Sarcoma
C1880052|Chemotherapy Regimen Used to Treat Malignant Renal Neoplasm
C1880052|Chemotherapy Regimen Used to Treat Kidney Cancer
C1880055|Chemotherapy Regimen Used to Treat Non-Hodgkin Lymphoma
C1880056|Chemotherapy Regimen Used to Treat Non-Small Cell Lung Carcinoma
C1880053|Chemotherapy Regimen Used to Treat Malignant Testicular Neoplasm
C1880053|Chemotherapy Regimen Used to Treat Testicular Cancer
C1880035|Chemotherapy Regimen Used to Treat Bladder Carcinoma
C1880032|Chemotherapy Regimen Used to Treat Acute Lymphoblastic Leukemia
C1880036|Chemotherapy Regimen Used to Treat Breast Carcinoma
C1880054|Chemotherapy Regimen Used to Treat Melanoma
C1880044|Chemotherapy Regimen Used to Treat Colorectal Carcinoma
C1880037|Chemotherapy Regimen Used to Treat Cervical Carcinoma
C1880048|Chemotherapy Regimen Used to Treat Gastric Carcinoma
C1880058|Chemotherapy Regimen Used to Treat Malignant Ovarian Neoplasm
C1880050|Chemotherapy Regimen Used to Treat Malignant Head and Neck Neoplasm
C1880049|Chemotherapy Regimen Used to Treat Hodgkins Lymphoma
C1880045|Chemotherapy Regimen Used to Treat Endometrial Carcinoma
C1880061|Chemotherapy Regimen Used to Treat Liver Cancer
C1880061|Chemotherapy Regimen Used to Treat Primary Malignant Neoplasm of Liver
C1880046|Chemotherapy Regimen Used to Treat Esophageal Carcinoma
C1880059|Chemotherapy Regimen Used to Treat Pancreatic Carcinoma
C1880059|Chemotherapy Regimen Used to Treat Pancreatic Cancer
C1880062|Chemotherapy Regimen Used to Treat Prostate Carcinoma
C2347611|Chemotherapy Regimen Used to Treat Gestational Trophoblastic Tumor
C0152018|CARCINOMA OF ESOPHAGUS
C0152018|ESOPHAGEAL CARCINOMA
C0152018|ESOPHAGEAL CANCER
C0152018|carcinoma of esophagus (diagnosis)
C0152018|Carcinoma;oesophagus
C0152018|Carcinoma of oesophagus
C0152018|Carcinoma of oesophagus (disorder)
C0152018|Cancer of oesophagus
C0152018|Carcinoma of esophagus (disorder)
C0152018|Esophageal cancer, NOS
C0152018|Esophageal carcinoma NOS
C0152018|Carcinoma of oesophagus NOS
C0152018|Carcinoma of esophagus NOS
C0152018|Oesophageal carcinoma
C0152018|Oesophageal carcinoma NOS
C0152018|Cancer of Esophagus
C0152018|Cancer of the Esophagus
C0152018|Esophagus Carcinoma
C0152018|Carcinoma of the Esophagus
C0152018|Carcinoma;esophagus
C0152018|carcinoma of the oesophagus
C0496775|Abdominal part of esophagus
C0496775|Abdominal part of oesophagus
C0496775|Malignant neoplasm of abdominal part of esophagus
C0496775|Malignant neoplasm of abdominal part of oesophagus
C0496775|malignant neoplasm of abdominal esophagus
C0496775|malignant neoplasm of abdominal esophagus (diagnosis)
C0496775|malignant tumor of abdominal esophagus
C0496775|Mal neo abdomin esophag
C0496775|Malignant neoplasm of abdominal oesophagus
C0496775|Malignant tumor of abdominal part of esophagus
C0496775|Malignant tumour of abdominal part of oesophagus
C0496775|Malignant tumor of abdominal part of esophagus (disorder)
C0496775|Malignant Neoplasm of the Abdominal Esophagus
C0496775|Malignant Tumor of the Abdominal Esophagus
C0496773|Cervical part of esophagus
C0496773|Cervical part of oesophagus
C0496773|Malignant neoplasm of cervical part of esophagus
C0496773|Malignant neoplasm of cervical part of oesophagus
C0496773|malignant neoplasm of cervical esophagus (diagnosis)
C0496773|malignant neoplasm of cervical esophagus
C0496773|malignant tumor of cervical esophagus
C0496773|Mal neo cervical esophag
C0496773|Malignant neoplasm of cervical oesophagus
C0496773|Malignant tumor of cervical part of esophagus
C0496773|Malignant tumour of cervical part of oesophagus
C0496773|Malignant tumor of cervical part of esophagus (disorder)
C0496773|Malignant Neoplasm of the Cervical Esophagus
C0153411|Malignant neoplasm of thoracic esophagus
C0153411|Malignant neoplasm of thoracic part of esophagus
C0153411|Malignant neoplasm of thoracic part of oesophagus
C0153411|Thoracic part of esophagus
C0153411|Thoracic part of oesophagus
C0153411|malignant neoplasm of thoracic esophagus (diagnosis)
C0153411|malignant tumor of thoracic esophagus
C0153411|Mal neo thoracic esophag
C0153411|Malignant neoplasm of thoracic oesophagus
C0153411|Malignant tumor of thoracic part of esophagus
C0153411|Malignant tumour of thoracic part of oesophagus
C0153411|Malignant tumor of thoracic part of esophagus (disorder)
C0153411|Malignant Neoplasm of the Thoracic Esophagus
C0153416|Malignant neoplasm of other specified part of esophagus
C0153416|Malignant neoplasm of other specified part of oesophagus
C0153416|Mal neo esophagus NEC
C0153416|Malignant neoplasm of other specified part of esophagus (disorder)
C0153413|Malignant neoplasm of upper third of esophagus
C0153413|Upper third of esophagus
C0153413|Malignant neoplasm of upper third of oesophagus
C0153413|Upper third of oesophagus
C0153413|Malignant neoplasm of upper third esophagus
C0153413|malignant neoplasm of upper third of esophagus (diagnosis)
C0153413|malignant tumor of upper third of esophagus
C0153413|Mal neo upper 3rd esoph
C0153413|Malignant tumour of upper third of oesophagus
C0153413|Malignant tumor of upper third of esophagus (disorder)
C0153413|Malignant Neoplasm of Proximal Third of Esophagus
C0153413|Malignant Neoplasm of the Proximal Third of the Esophagus
C0153413|Malignant Neoplasm of the Upper Third of the Esophagus
C0153413|Malignant Tumor of Proximal Third of Esophagus
C0153413|Malignant Tumor of the Proximal Third of the Esophagus
C0153413|Malignant Tumor of the Upper Third of the Esophagus
C0153415|Malignant neoplasm of lower third of esophagus
C0153415|Lower third of esophagus
C0153415|Lower third of oesophagus
C0153415|Malignant neoplasm of lower third of oesophagus
C0153415|malignant neoplasm of lower third of esophagus (diagnosis)
C0153415|malignant tumor of lower third of esophagus
C0153415|Mal neo lower 3rd esoph
C0153415|Ca lower third esophagus (disorder)
C0153415|Ca lower third esophagus
C0153415|Ca lower third oesophagus
C0153415|Ca lower third oesophagus (disorder)
C0153415|Malignant tumour of lower third of oesophagus
C0153415|Malignant tumor of lower third of esophagus (disorder)
C0153415|Malignant Lower Third of Esophagus Neoplasm
C0153415|Malignant Lower Third of Esophagus Tumor
C0153415|Malignant Lower Third of the Esophagus Neoplasm
C0153415|Malignant Lower Third of the Esophagus Tumor
C0153415|Malignant Neoplasm of Distal Third of Esophagus
C0153415|Malignant Neoplasm of the Distal Third of the Esophagus
C0153415|Malignant Neoplasm of the Lower Third of the Esophagus
C0153415|Malignant Tumor of Distal Third of Esophagus
C0153415|Malignant Tumor of the Distal Third of the Esophagus
C0153415|Malignant Tumor of the Lower Third of the Esophagus
C0153414|Malignant neoplasm of middle third of esophagus
C0153414|Middle third of esophagus
C0153414|Malignant neoplasm of middle third of oesophagus
C0153414|Middle third of oesophagus
C0153414|malignant neoplasm of middle third of esophagus (diagnosis)
C0153414|malignant tumor of middle third of esophagus
C0153414|Mal neo middle 3rd esoph
C0153414|Ca middle third esophagus (disorder)
C0153414|Ca middle third oesophagus
C0153414|Ca middle third oesophagus (disorder)
C0153414|Ca middle third esophagus
C0153414|Malignant tumour of middle third of oesophagus
C0153414|Malignant tumor of middle third of esophagus (disorder)
C0153414|Malignant Middle Third of Esophagus Neoplasm
C0153414|Malignant Middle Third of Esophagus Tumor
C0153414|Malignant Middle Third of the Esophagus Neoplasm
C0153414|Malignant Middle Third of the Esophagus Tumor
C0153414|Malignant Neoplasm of the Middle Third of the Esophagus
C0153414|Malignant Tumor of the Middle Third of the Esophagus
C0546837|Malignant neoplasm of esophagus
C0546837|Cancer of esophagus
C0546837|Malignant neoplasm of esophagus, unspecified
C0546837|Esophagus, unspecified
C0546837|Malignant neoplasm of oesophagus
C0546837|Malignant neoplasm of oesophagus, unspecified
C0546837|Oesophagus, unspecified
C0546837|malignant neoplasm of esophagus (diagnosis)
C0546837|esophageal cancer
C0546837|esophageal cancer (diagnosis)
C0546837|malignant esophageal neoplasm
C0546837|Ca esophagus
C0546837|Oesophageal neoplasms malignant
C0546837|Cancer, Esophageal
C0546837|Cancers, Esophageal
C0546837|Esophageal Cancers
C0546837|Cancers, Esophagus
C0546837|Esophagus Cancers
C0546837|malignant tumor of esophagus
C0546837|Mal neo esophagus NOS
C0546837|Cancer, Esophagus
C0546837|Malignant neoplasm of esophagus, unspecified site
C0546837|Oesophageal cancer
C0546837|Malignant neoplasm of oesophagus NOS
C0546837|Ca esophagus NOS (disorder)
C0546837|Ca esophagus NOS
C0546837|(Malignant neoplasm of oesophagus NOS or oesophageal cancer
C0546837|Malignant neoplasm of esophagus NOS
C0546837|Ca oesophagus NOS
C0546837|Ca oesophagus NOS (disorder)
C0546837|CA - Cancer of esophagus
C0546837|CA - Cancer of oesophagus
C0546837|Cancer of oesophagus
C0546837|Malignant tumour of oesophagus
C0546837|Malignant tumour of oesophagus (disorder)
C0546837|(Malignant neoplasm of esophagus NOS or esophageal cancer
C0546837|(Malignant neoplasm of oesophagus NOS or oesophageal cancer (disorder)
C0546837|Malignant neoplasm of esophagus NOS (disorder)
C0546837|Esophagus--Cancer
C0546837|-- Esophageal Cancer
C0546837|Oesophageal cancer NOS
C0546837|Esophageal cancer NOS
C0546837|Esophagus Cancer
C0546837|Cancer of the Esophagus
C0546837|Ca oesophagus
C0546837|Malignant tumor of esophagus (disorder)
C0546837|Malignant neoplasm of esophagus, NOS
C0546837|Malignant Esophageal Tumor
C0546837|Malignant Esophagus Tumor
C0546837|Malignant Neoplasm of the Esophagus
C0546837|Malignant Tumor of the Esophagus
C0546837|Esophageal neoplasms malignant
C0546837|Neoplasm malig;esophagus
C0546837|Neoplasm malig;oesophagus
C0546837|malignant neosplasm of the esophagus
C0546837|malignant neosplasm of the oesophagus
C0496776|Malignant neoplasm overlapping esophagus site
C0496776|Malignant neoplasm overlapping oesophagus site
C0496776|Overlapping lesion of esophagus
C0496776|Overlapping lesion of oesophagus
C0496776|Malignant neoplasm of overlapping sites of esophagus
C0496776|esophageal neoplasm malignant overlapping sites of esophagus
C0496776|malignant neoplasm of overlapping sites of esophagus (diagnosis)
C0279628|adenocarcinoma of esophagus (diagnosis)
C0279628|adenocarcinoma of esophagus
C0279628|esophageal adenocarcinoma
C0279628|Adenocarcinoma - esophagus
C0279628|Adenocarcinoma of the esophagus
C0279628|Esophageal adenocarcinoma NOS
C0279628|Oesophageal adenocarcinoma
C0279628|Oesophageal adenocarcinoma NOS
C0279628|Adenocarcinoma of oesophagus
C0279628|Adenocarcinoma of esophagus (disorder)
C0279628|esophageal cancer, adenocarcinoma
C0279628|esophagus cancer, adenocarcinoma
C0279628|Esophagus Adenocarcinoma
C0854762|Oesophageal adenocarcinoma recurrent
C0854762|Esophageal adenocarcinoma recurrent
C0854762|Esophageal Adenocarcinoma, Recurrent
C0854762|Recurrent Adenocarcinoma of Esophagus
C0854762|Recurrent Adenocarcinoma of the Esophagus
C0854762|Recurrent Esophageal Adenocarcinoma
C0854762|Recurrent Esophagus Adenocarcinoma
C0854762|Relapsed Adenocarcinoma of Esophagus
C0854762|Relapsed Adenocarcinoma of the Esophagus
C0854762|Relapsed Esophageal Adenocarcinoma
C0854762|Relapsed Esophagus Adenocarcinoma
C0854764|adenocarcinoma in situ of esophagus (diagnosis)
C0854764|adenocarcinoma in situ of esophagus
C0854764|Oesophageal adenocarcinoma stage 0
C0854764|Stage 0 Esophageal Adenocarcinoma AJCC v7
C0854764|Stage 0 Esophageal Adenocarcinoma
C0854764|Oesophageal adenocarcinoma site unspecified stage 0
C0854764|Esophageal adenocarcinoma in situ
C0854764|Oesophageal adenocarcinoma site unspecified in situ
C0854764|Esophageal adenocarcinoma site unspecified stage 0
C0854764|Esophageal adenocarcinoma stage 0
C0854764|Esophageal adenocarcinoma site unspecified in situ
C0854764|Oesophageal adenocarcinoma in situ
C0854764|Esophageal Adenocarcinoma, Stage 0
C0854764|Adenocarcinoma in situ of the Esophagus
C0854764|Esophagus Adenocarcinoma in situ
C0854764|Stage 0 Adenocarcinoma of Esophagus
C0854764|Stage 0 Adenocarcinoma of the Esophagus
C0854764|Stage 0 Esophagus Adenocarcinoma
C0854765|Oesophageal adenocarcinoma stage I
C0854765|Stage I Esophageal Adenocarcinoma AJCC v7
C0854765|Stage I Esophageal Adenocarcinoma
C0854765|Esophageal adenocarcinoma site unspecified stage I
C0854765|Esophageal adenocarcinoma stage I
C0854765|Oesophageal adenocarcinoma site unspecified stage I
C0854765|Esophageal Adenocarcinoma, Stage I
C0854765|Stage I Adenocarcinoma of Esophagus
C0854765|Stage I Adenocarcinoma of the Esophagus
C0854765|Stage I Esophagus Adenocarcinoma
C0854763|Oesophageal adenocarcinoma stage II
C0854763|Stage II Esophageal Adenocarcinoma AJCC v7
C0854763|Stage II Esophageal Adenocarcinoma
C0854763|Esophageal adenocarcinoma site unspecified stage II
C0854763|Esophageal adenocarcinoma stage II
C0854763|Oesophageal adenocarcinoma site unspecified stage II
C0854763|Esophageal Adenocarcinoma, Stage II
C0854763|Stage II Adenocarcinoma of Esophagus
C0854763|Stage II Adenocarcinoma of the Esophagus
C0854763|Stage II Esophagus Adenocarcinoma
C0854766|Oesophageal adenocarcinoma stage III
C0854766|Stage III Esophageal Adenocarcinoma AJCC v7
C0854766|Stage III Esophageal Adenocarcinoma
C0854766|Esophageal adenocarcinoma stage III
C0854766|Oesophageal adenocarcinoma site unspecified stage III
C0854766|Esophageal adenocarcinoma site unspecified stage III
C0854766|Esophageal Adenocarcinoma, Stage III
C0854766|Stage III Adenocarcinoma of Esophagus
C0854766|Stage III Adenocarcinoma of the Esophagus
C0854766|Stage III Esophagus Adenocarcinoma
C1142347|Oesophageal adenocarcinoma stage IV
C1142347|Stage IV Esophageal Adenocarcinoma AJCC v7
C1142347|Stage IV Esophageal Adenocarcinoma
C1142347|Oesophageal adenocarcinoma metastatic
C1142347|Esophageal adenocarcinoma metastatic
C1142347|Esophageal adenocarcinoma site unspecified stage IV
C1142347|Oesophageal adenocarcinoma site unspecified stage IV
C1142347|Esophageal adenocarcinoma stage IV
C1142347|Esophageal Adenocarcinoma, Stage IV
C1142347|Metastatic Adenocarcinoma of Esophagus
C1142347|Metastatic Adenocarcinoma of the Esophagus
C1142347|Metastatic Esophageal Adenocarcinoma
C1142347|Metastatic Esophagus Adenocarcinoma
C1142347|Stage IV Adenocarcinoma of Esophagus
C1142347|Stage IV Adenocarcinoma of the Esophagus
C1142347|Stage IV Esophagus Adenocarcinoma
C0854761|Oesophageal carcinoma recurrent
C0854761|Recurrent Esophageal Cancer
C0854761|Recurrent Esophageal Carcinoma
C0854761|Oesophageal carcinoma site unspecified recurrent
C0854761|Esophageal carcinoma recurrent
C0854761|Esophageal carcinoma site unspecified recurrent
C0854761|esophageal cancer, recurrent
C0854761|esophagus cancer, recurrent
C0854761|Esophageal Carcinoma, Recurrent
C0854761|Recurrent Cancer of Esophagus
C0854761|Recurrent Cancer of the Esophagus
C0854761|Recurrent Carcinoma of Esophagus
C0854761|Recurrent Carcinoma of the Esophagus
C0854761|Recurrent Esophagus Cancer
C0854761|Relapsed Cancer of Esophagus
C0854761|Relapsed Cancer of the Esophagus
C0854761|Relapsed Carcinoma of Esophagus
C0854761|Relapsed Carcinoma of the Esophagus
C0854761|Relapsed Esophageal Cancer
C0854761|Relapsed Esophagus Carcinoma
C0154059|Esophagus
C0154059|Carcinoma in situ of esophagus
C0154059|Carcinoma in situ of oesophagus
C0154059|Oesophagus
C0154059|carcinoma in situ of esophagus (diagnosis)
C0154059|Ca in situ esophagus
C0154059|Esophageal Carcinoma in situ AJCC v7
C0154059|Severe Esophageal Dysplasia AJCC v7
C0154059|Severe Esophageal Dysplasia
C0154059|Stage 0 Esophageal Cancer AJCC v7
C0154059|Esophageal Carcinoma in situ
C0154059|Stage 0 Esophageal Cancer
C0154059|Carcinoma in situ of esophagus NOS
C0154059|Carcinoma in situ of oesophagus NOS
C0154059|Carcinoma in situ of esophagus NOS (disorder)
C0154059|stage 0 esophageal carcinoma in situ
C0154059|Cancer in situ of esophagus
C0154059|Cancer in situ of oesophagus
C0154059|Oesophageal carcinoma NOS stage 0
C0154059|Esophageal carcinoma stage 0
C0154059|Esophageal carcinoma site unspecified stage 0
C0154059|Oesophageal carcinoma site unspecified stage 0
C0154059|Oesophageal carcinoma in situ
C0154059|Oesophageal carcinoma stage 0
C0154059|Esophageal carcinoma NOS stage 0
C0154059|Severe oesophageal dysplasia
C0154059|Carcinoma in situ of esophagus (disorder)
C0154059|Severe esophageal dysplasia (disorder)
C0154059|esophageal cancer, stage 0
C0154059|esophagus cancer, stage 0
C0154059|Carcinoma in situ of esophagus, NOS
C0854769|Oesophageal squamous cell carcinoma recurrent
C0854769|Esophageal squamous cell carcinoma site unspecified recurrent
C0854769|Esophageal squamous cell carcinoma recurrent
C0854769|Oesophageal squamous cell carcinoma site unspecified recurrent
C0854769|Recurrent Esophageal Squamous Cell Carcinoma
C0854769|Recurrent Squamous Cell Carcinoma of Esophagus
C0854769|Recurrent Squamous Cell Carcinoma of the Esophagus
C0854770|squamous cell carcinoma in situ of esophagus (diagnosis)
C0854770|squamous cell carcinoma in situ of esophagus
C0854770|Oesophageal squamous cell carcinoma stage 0
C0854770|Stage 0 Esophageal Squamous Cell Carcinoma AJCC v7
C0854770|Stage 0 Esophageal Squamous Cell Carcinoma
C0854770|Oesophageal squamous cell carcinoma in situ
C0854770|Esophageal squamous cell carcinoma in situ
C0854770|Esophageal squamous cell carcinoma stage 0
C0854770|Esophagus Squamous Cell Carcinoma in situ
C0854770|Squamous Cell Carcinoma in situ of the Esophagus
C0854770|Stage 0 Esophagus Squamous Cell Carcinoma
C0854770|Stage 0 Squamous Cell Carcinoma of Esophagus
C0854770|Stage 0 Squamous Cell Carcinoma of the Esophagus
C0854771|Oesophageal squamous cell carcinoma stage I
C0854771|Stage I Esophageal Squamous Cell Carcinoma AJCC v7
C0854771|Stage I Esophageal Squamous Cell Carcinoma
C0854771|Esophageal squamous cell carcinoma site unspecified stage I
C0854771|Esophageal squamous cell carcinoma stage I
C0854771|Oesophageal squamous cell carcinoma site unspecified stage I
C0854771|Stage I Esophagus Squamous Cell Carcinoma
C0854771|Stage I Squamous Cell Carcinoma of Esophagus
C0854771|Stage I Squamous Cell Carcinoma of the Esophagus
C0854772|Oesophageal squamous cell carcinoma stage II
C0854772|Stage II Esophageal Squamous Cell Carcinoma AJCC v7
C0854772|Stage II Esophageal Squamous Cell Carcinoma
C0854772|Esophageal squamous cell carcinoma site unspecified stage II
C0854772|Oesophageal squamous cell carcinoma site unspecified stage II
C0854772|Esophageal squamous cell carcinoma stage II
C0854772|Stage II Esophagus Squamous Cell Carcinoma
C0854772|Stage II Squamous Cell Carcinoma of Esophagus
C0854772|Stage II Squamous Cell Carcinoma of the Esophagus
C0854773|Oesophageal squamous cell carcinoma stage III
C0854773|Stage III Esophageal Squamous Cell Carcinoma AJCC v7
C0854773|Stage III Esophageal Squamous Cell Carcinoma
C0854773|Esophageal squamous cell carcinoma stage III
C0854773|Stage III Esophagus Squamous Cell Carcinoma
C0854773|Stage III Squamous Cell Carcinoma of Esophagus
C0854773|Stage III Squamous Cell Carcinoma of the Esophagus
C1142025|Oesophageal squamous cell carcinoma stage IV
C1142025|Stage IV Esophageal Squamous Cell Carcinoma AJCC v7
C1142025|Stage IV Esophageal Squamous Cell Carcinoma
C1142025|Oesophageal squamous cell carcinoma metastatic
C1142025|Oesophageal squamous cell carcinoma site unspecified stage IV
C1142025|Esophageal squamous cell carcinoma metastatic
C1142025|Esophageal squamous cell carcinoma site unspecified stage IV
C1142025|Esophageal squamous cell carcinoma stage IV
C1142025|Metastatic Esophageal Squamous Cell Carcinoma
C1142025|Metastatic Esophagus Squamous Cell Carcinoma
C1142025|Metastatic Squamous Cell Carcinoma of Esophagus
C1142025|Metastatic Squamous Cell Carcinoma of the Esophagus
C1142025|Stage IV Esophagus Squamous Cell Carcinoma
C1142025|Stage IV Squamous Cell Carcinoma of Esophagus
C1142025|Stage IV Squamous Cell Carcinoma of the Esophagus
C0278562|Stage IV Esophageal Cancer AJCC v7
C0278562|Stage IV Esophageal Cancer
C0278562|Oesophageal cancer metastatic
C0278562|Oesophageal neoplasm metastatic
C0278562|Esophageal neoplasm metastatic
C0278562|Esophageal cancer metastatic
C0278562|esophageal cancer, metastatic
C0278562|esophageal cancer, stage IV
C0278562|esophagus cancer, metastatic
C0278562|esophagus cancer, stage IV
C0278562|metastatic esophageal cancer
C0279626|Squamous cell carcinoma of esophagus
C0279626|squamous cell carcinoma of esophagus (diagnosis)
C0279626|ESCC
C0279626|Esophageal Squamous Cell Carcinoma
C0279626|Squamous cell car. - esophagus
C0279626|Squamous cell carcinoma of the esophagus
C0279626|Oesophageal squamous cell carcinoma stage unspecified
C0279626|Squamous cell carcinoma of oesophagus
C0279626|Esophageal squamous cell carcinoma stage unspecified
C0279626|Oesophageal squamous cell carcinoma NOS
C0279626|Esophageal squamous cell carcinoma NOS
C0279626|Squamous cell carcinoma of esophagus NOS
C0279626|Oesophageal epidermoid carcinoma NOS
C0279626|Oesophageal squamous cell carcinoma
C0279626|Esophageal epidermoid carcinoma NOS
C0279626|SCC - Squamous cell carcinoma of esophagus
C0279626|SCC - Squamous cell carcinoma of oesophagus
C0279626|Squamous cell carcinoma of esophagus (disorder)
C0279626|esophageal cancer, squamous cell
C0279626|esophagus cancer, squamous cell
C0279626|squamous cell esophageal cancer
C0279626|squamous cell esophagus cancer
C0279626|Esophageal Epidermoid Carcinoma
C0279626|Esophageal SCC
C0279626|Esophagus SCC
C0279626|Esophagus Squamous Cell Carcinoma
C0279626|SCC of Esophagus
C0279626|SCC of the Esophagus
C2204789|malignant small cell neoplasm of esophagus (diagnosis)
C2204789|malignant small cell neoplasm of esophagus
C2011363|giant cell type neoplasm of esophagus
C2011363|giant cell type neoplasm of esophagus (diagnosis)
C2018647|spindle cell type neoplasm of esophagus (diagnosis)
C2018647|spindle cell type neoplasm of esophagus
C2075606|clear cell type neoplasm of esophagus (diagnosis)
C2075606|clear cell type neoplasm of esophagus
C2204810|myosarcoma of esophagus
C2204810|myosarcoma of esophagus (diagnosis)
C2204823|malignant plasmacytoma of esophagus (diagnosis)
C2204823|malignant plasmacytoma of esophagus
C2204825|malignant mastocytosis of esophagus
C2204825|malignant mastocytosis of esophagus (diagnosis)
C1333466|sarcoma of esophagus (diagnosis)
C1333466|sarcoma of esophagus
C1333466|Esophageal Sarcoma
C1333466|Esophagus Sarcoma
C1333466|Sarcoma of the Esophagus
C1333466|Sarcoma, Esophagus
C2216771|malignant neoplasm of esophagus staging (diagnosis)
C2216771|malignant neoplasm of esophagus staging
C2216771|malignant esophageal neoplasm staging
C2216771|malignant tumor of esophagus staging
C2216771|esophageal cancer staging
C2062505|malignant lymphoma of esophagus (diagnosis)
C2062505|malignant lymphoma of esophagus
C1333453|Esophageal Kaposi Sarcoma
C1333453|Esophageal Kaposi's Sarcoma
C1333453|Kaposi's sarcoma of esophagus (diagnosis)
C1333453|Kaposi's sarcoma of esophagus
C1333453|Esophagus Kaposi's Sarcoma
C1333453|Kaposi's Sarcoma of the Esophagus
C1333463|neurofibroma of esophagus
C1333463|neurofibroma of esophagus (diagnosis)
C1333463|esophageal neurofibroma
C1333463|Esophagus Neurofibroma
C1333463|Neurofibroma of the Esophagus
C2007067|carcinosarcoma of esophagus (diagnosis)
C2007067|carcinosarcoma of esophagus
C1333444|malignant carcinoid tumor of esophagus (diagnosis)
C1333444|malignant carcinoid tumor of esophagus
C1333444|Esophageal Neuroendocrine Tumor G1
C1333444|Esophageal NET G1 (Carcinoid)
C1333444|Esophageal Carcinoid Tumor
C1333444|Esophageal Neuroendocrine Tumor G1 (Carcinoid)
C1333444|Esophageal NET G1
C1333444|Carcinoid Tumor of Esophagus
C1333444|Carcinoid Tumor of the Esophagus
C2204829|balloon cell melanoma of esophagus (diagnosis)
C2204829|balloon cell melanoma of esophagus
C2063891|melanoma of skin of esophagus
C2063891|melanoma of skin of esophagus (diagnosis)
C2984901|Malignant Esophageal Peripheral Nerve Sheath Tumor
C2216772|malignant neoplasm of esophagus TNM staging
C2216772|malignant neoplasm of esophagus TNM staging (diagnosis)
C2216772|esophageal cancer TNM staging
C2216772|malignant tumor of esophagus TNM staging
C2216783|malignant neoplasm of esophagus TNM staging regional lymph nodes (N) (diagnosis)
C2216783|malignant neoplasm of esophagus TNM staging regional lymph nodes (N)
C2216783|malignant esophageal neoplasm TNM staging of regional lymph nodes (N)
C2216783|esophageal cancer TNM staging regional lymph nodes (N)
C2216783|malignant tumor of esophagus TNM staging regional lymph nodes (N)
C2216784|malignant neoplasm of esophagus TNM staging regional lymph nodes (N) N0 (diagnosis)
C2216784|malignant neoplasm of esophagus TNM staging regional lymph nodes (N) N0
C2216784|malignant esophageal neoplasm N0
C2216784|esophageal cancer TNM staging regional lymph nodes (N) N0
C2216784|malignant tumor of esophagus TNM staging regional lymph nodes (N) N0
C2216785|malignant neoplasm of esophagus TNM staging regional lymph nodes (N) N1 (diagnosis)
C2216785|malignant neoplasm of esophagus TNM staging regional lymph nodes (N) N1
C2216785|malignant esophageal neoplasm N1
C2216785|malignant tumor of esophagus TNM staging regional lymph nodes (N) N1
C2216785|esophageal cancer TNM staging regional lymph nodes (N) N1
C2216776|malignant neoplasm of esophagus TNM staging distant metastasis (M) (diagnosis)
C2216776|malignant neoplasm of esophagus TNM staging distant metastasis (M)
C2216776|malignant esophageal neoplasm TNM staging of distant metastasis (M)
C2216776|malignant tumor of esophagus TNM staging distant metastasis (M)
C2216776|esophageal cancer TNM staging distant metastasis (M)
C2216775|malignant neoplasm of esophagus TNM staging distal metastasis (M) M1b
C2216775|malignant neoplasm of esophagus TNM staging distal metastasis (M) M1b (diagnosis)
C2216775|malignant esophageal neoplasm M1b
C2216775|malignant tumor of esophagus TNM staging distal metastasis (M) M1b
C2216775|esophageal cancer TNM staging distal metastasis (M) M1b
C2216773|malignant neoplasm of esophagus TNM staging distal metastasis (M) M0 (diagnosis)
C2216773|malignant neoplasm of esophagus TNM staging distal metastasis (M) M0
C2216773|malignant esophageal neoplasm M0
C2216773|malignant tumor of esophagus TNM staging distal metastasis (M) M0
C2216773|esophageal cancer TNM staging distal metastasis (M) M0
C2216774|malignant neoplasm of esophagus TNM staging distal metastasis (M) M1a
C2216774|malignant neoplasm of esophagus TNM staging distal metastasis (M) M1a (diagnosis)
C2216774|malignant esophageal neoplasm M1a
C2216774|esophageal cancer TNM staging distal metastasis (M) M1a
C2216774|malignant tumor of esophagus TNM staging distal metastasis (M) M1a
C3165092|Leiomyosarcoma of lower esophagus
C3165092|Leiomyosarcoma of lower esophagus (disorder)
C3165092|Leiomyosarcoma of lower oesophagus
C3165092|malignant neoplasm myosarcoma leiomyosarcoma lower esophagus
C3165092|Leiomyosarcoma of lower esophagus (diagnosis)
C3165036|Lymphoma of lower esophagus (disorder)
C3165036|Lymphoma of lower esophagus
C3165036|Lymphoma of lower oesophagus
C3165036|esophageal malignant lymphoma of lower esophagus
C3165036|Lymphoma of lower esophagus (diagnosis)
C2111603|large cell carcinoma of esophagus (diagnosis)
C2111603|large cell carcinoma of esophagus
C2111715|large cell neuroendocrine carcinoma of esophagus
C2111715|large cell neuroendocrine carcinoma of esophagus (diagnosis)
C2111604|large cell carcinoma of esophagus with rhabdoid phenotype (diagnosis)
C2111604|large cell carcinoma of esophagus with rhabdoid phenotype
C2012076|glassy cell carcinoma of esophagus (diagnosis)
C2012076|glassy cell carcinoma of esophagus
C2188058|undifferentiated carcinoma of esophagus (diagnosis)
C2188058|undifferentiated carcinoma of esophagus
C2188058|Esophageal Undifferentiated Carcinoma
C2009877|fusiform type small cell carcinoma of esophagus (diagnosis)
C2009877|fusiform type small cell carcinoma of esophagus
C2037374|superficial spreading melanoma of esophagus
C2037374|superficial spreading melanoma of esophagus (diagnosis)
C2204836|mixed epithelioid and spindle cell melanoma of esophagus (diagnosis)
C2204836|mixed epithelioid and spindle cell melanoma of esophagus
C2063886|adenosquamous carcinoma of esophagus
C2063886|adenosquamous carcinoma of esophagus (diagnosis)
C2063886|Esophageal Adenosquamous Carcinoma
C1333441|adenoid cystic carcinoma of esophagus
C1333441|adenoid cystic carcinoma of esophagus (diagnosis)
C1333441|Esophageal Adenoid Cystic Carcinoma
C1333441|Esophagus Adenoid Cystic Carcinoma
C1333441|Adenoid Cystic Carcinoma of the Esophagus
C1333441|Adenoid Cystic Carcinoma, Esophagus
C1333441|Adenoid Cystic Esophagus Carcinoma
C1333461|mucoepidermoid carcinoma of esophagus
C1333461|mucoepidermoid carcinoma of esophagus (diagnosis)
C1333461|Esophageal Mucoepidermoid Carcinoma
C1333461|Mucoepidermoid Carcinoma of the Esophagus
C1333461|Mucoepidermoid Esophageal Carcinoma
C1333461|Mucoepidermoid Esophagus Carcinoma
C2237936|X-ray UGI Ba swallow- esophageal mass malignant neoplasm ___
C2237936|barium swallow: malignant neoplasm of esophagus
C2237936|barium swallow: malignant neoplasm of esophagus (procedure)
C2204790|malignant epithelioma of esophagus (diagnosis)
C2204790|malignant epithelioma of esophagus
C2204834|epithelioid cell melanoma of esophagus (diagnosis)
C2204834|epithelioid cell melanoma of esophagus
C1282473|local recurrence of malignant neoplasm of esophagus
C1282473|esophageal malignant neoplasm, local recurrence
C1282473|local recurrence of malignant neoplasm of esophagus (diagnosis)
C1282473|Local recurrence of malignant tumor of esophagus (disorder)
C1282473|Local recurrence of malignant tumor of esophagus
C1282473|Local recurrence of malignant tumour of oesophagus
C0349048|Malignant neoplasm, overlapping lesion of esophagus
C0349048|Malignant neoplasm, overlapping lesion of oesophagus
C0349048|Malignant neoplasm, overlapping lesion of esophagus (disorder)
C0349048|Overlapping malignant neoplasm of esophagus (disorder)
C0349048|Overlapping malignant neoplasm of esophagus
C0349048|Overlapping malignant neoplasm of oesophagus
C0346619|Malignant neoplasm of cardioesophageal junction of stomach
C0346619|Malignant neoplasm of gastro-esophageal junction
C0346619|malignant neoplasm of cardioesophageal junction of stomach (diagnosis)
C0346619|esophageal neoplasm malignant cardioesophageal junction of stomach
C0346619|Malignant neoplasm of cardio-esophageal junction of stomach
C0346619|Malignant neoplasm of cardio-oesophageal junction of stomach
C0346619|Malignant neoplasm of gastro-oesophageal junction
C0346619|Malignant neoplasm of cardioesophageal junction of stomach (disorder)
C1300083|Primary malignant neoplasm of oesophagus
C1300083|Primary malignant neoplasm of esophagus (disorder)
C1300083|Primary malignant neoplasm of esophagus
C1300083|Primary malignant neoplasm of esophagus (diagnosis)
C1300083|esophageal malignant neoplasm primary
C0686055|Metastatic Neoplasm to the Esophagus
C0686055|Metastases to oesophagus
C0686055|esophageal malignant neoplasm secondary
C0686055|Secondary malignant neoplasm of esophagus
C0686055|Secondary malignant neoplasm of esophagus (diagnosis)
C0686055|Metastatic Malignant Neoplasm to the Esophagus
C0686055|Metastatic Malignant Neoplasm in the Esophagus
C0686055|Cancer metastatic to esophagus
C0686055|Metastases to esophagus
C0686055|Metastatic malignant neoplasm to esophagus
C0686055|Secondary malignant neoplasm of esophagus (disorder)
C0686055|Secondary malignant neoplasm of oesophagus
C0686055|Metastatic malignant neoplasm to oesophagus
C0686055|Metastatic malignant neoplasm to esophagus, NOS
C0686055|Secondary malignant neoplasm of esophagus, NOS
C0686055|Esophageal Metastasis
C0686055|Metastases to the Esophagus
C0686055|Metastasis to Esophagus
C0686055|Metastasis to the Esophagus
C0686055|Metastatic Tumor to the Esophagus
C4065138|esophagoscopy mass malignant neoplasm
C4065138|esophagoscopy mass malignant neoplasm (procedure)
C0346618|malignant neoplasm of esophagus, stomach, and duodenum
C0346618|digestive neoplasm malignant of esophagus, stomach, and duodenum
C0346618|malignant neoplasm of esophagus, stomach, and duodenum (diagnosis)
C0346618|Malignant tumor of esophagus, stomach and duodenum
C0346618|Malignant tumour of oesophagus, stomach and duodenum
C0346618|Malignant tumor of esophagus, stomach and duodenum (disorder)
C0279865|cellular diagnosis, esophageal cancer
C0279865|esophageal cancer, cellular diagnosis
C0279865|esophagus cancer cellular diagnosis
C0280257|stage, esophageal cancer
C0280257|esophageal cancer, stage
C1333459|Primary Esophageal Lymphoma
C1333459|Esophageal Lymphoma
C1333459|Esophagus Lymphoma
C1333459|Lymphoma of Esophagus
C1333459|Lymphoma of the Esophagus
C1334579|Malignant Esophageal Neoplasm by Topographic Region
C1333460|Esophageal Melanoma
C1333460|Esophagus Melanoma
C1333460|Melanoma of Esophagus
C1333460|Melanoma of the Esophagus
C1334578|Malignant Esophageal Neoplasm by Anatomic Region
C0585126|Perforated carcinoma of esophagus (diagnosis)
C0585126|esophageal neoplasm malignant carcinoma, perforated
C0585126|Perforated carcinoma of esophagus
C0585126|Perforated carcinoma of oesophagus
C0585126|Perforated carcinoma of esophagus (disorder)
C1276562|T3: Esophageal tumor invades adventitia (finding)
C1276562|T3: Esophageal tumor invades adventitia
C1276562|T3: Oesophageal tumour invades adventitia
C1276562|T3: Esophageal tumor invades adventitia (tumor staging)
C2204817|angioimmunoblastic T-cell lymphoma of esophagus
C2204817|angioimmunoblastic T-cell lymphoma of esophagus (diagnosis)
C2204817|angioimmunoblastic lymphadenopathy with dysproteinemia (AILD) of esophagus
C2204821|NK/T-cell lymphoma of esophagus
C2204821|NK/T-cell lymphoma of esophagus (diagnosis)
C2113687|precursor cell lymphoblastic lymphoma of esophagus (diagnosis)
C2113687|precursor cell lymphoblastic lymphoma of esophagus
C2204826|mast cell sarcoma of esophagus (diagnosis)
C2204826|mast cell sarcoma of esophagus
C2113618|precursor B-cell lymphoblastic lymphoma of esophagus
C2113618|precursor B-cell lymphoblastic lymphoma of esophagus (diagnosis)
C2204822|malignant histiocytosis of esophagus
C2204822|malignant histiocytosis of esophagus (diagnosis)
C2204837|Sezary syndrome of esophagus
C2204837|Sezary syndrome of esophagus (diagnosis)
C2204815|marginal zone B-cell lymphoma of esophagus
C2204815|marginal zone B-cell lymphoma of esophagus (diagnosis)
C2113758|precursor T-cell lymphoblastic lymphoma of esophagus (diagnosis)
C2113758|precursor T-cell lymphoblastic lymphoma of esophagus
C2204816|mature T-cell lymphoma of esophagus
C2204816|mature T-cell lymphoma of esophagus (diagnosis)
C0345819|gastric malignant carcinoma lesser curve
C0345819|Carcinoma of lesser curve of stomach (diagnosis)
C0345819|Carcinoma of lesser curve of stomach
C0345819|Carcinoma of lesser curve of stomach (disorder)
C0153423|Malignant neoplasm of greater curvature of stomach, unspecified
C0153423|Greater curvature of stomach, unspecified
C0153423|Malignant neoplasm of greater curvature of stomach
C0153423|malignant neoplasm of greater curvature of stomach (diagnosis)
C0153423|malignant tumor of greater curvature of stomach
C0153423|Mal neo stom great curv
C0153423|Malignant neoplasm of greater curvature of stomach, unsp
C0153423|Ca greater curvature - stomach
C0153423|Malignant neoplasm of greater curve of stomach unspecified
C0153423|Ca greater curvature - stomach (disorder)
C0153423|Malignant neoplasm of greater curve of stomach unspecified (disorder)
C0153423|Malignant tumor of greater curve of stomach
C0153423|Malignant tumour of greater curve of stomach
C0153423|Malignant tumor of greater curve of stomach (disorder)
C0153423|Malignant neoplasm of greater curvature of stomach, NOS
C0699791|Cancer of stomach
C0699791|carcinoma of stomach (diagnosis)
C0699791|carcinoma of stomach
C0699791|Gastric carcinoma
C0699791|Carcinoma;stomach
C0699791|GASTRIC CANCER
C0699791|Stomach Cancer
C0699791|Carcinoma of stomach (disorder)
C0699791|Gastric cancer, NOS
C0699791|Carcinoma gastric
C0699791|Carcinoma stomach
C0699791|Stomach carcinoma
C0699791|Stomach (gastric) cancer
C0699791|Cancer of the Stomach
C0699791|Carcinoma of the Stomach
C2204845|malignant epithelioma of stomach (diagnosis)
C2204845|malignant epithelioma of stomach
C2111678|large cell carcinoma of stomach (diagnosis)
C2111678|large cell carcinoma of stomach
C2012116|glassy cell carcinoma of stomach (diagnosis)
C2012116|glassy cell carcinoma of stomach
C1336858|undifferentiated carcinoma of stomach
C1336858|anaplastic carcinoma of stomach (diagnosis)
C1336858|undifferentiated carcinoma of stomach (diagnosis)
C1336858|anaplastic carcinoma of stomach
C1336858|undifferentiated gastric carcinoma
C1336858|Anaplastic Carcinoma of the Stomach
C1336858|Anaplastic Gastric Carcinoma
C1336858|Undifferentiated Carcinoma of the Stomach
C2082464|pleomorphic carcinoma of stomach
C2082464|pleomorphic carcinoma of stomach (diagnosis)
C2011266|giant cell carcinoma of stomach (diagnosis)
C2011266|giant cell carcinoma of stomach
C2018406|spindle cell carcinoma of stomach (diagnosis)
C2018406|spindle cell carcinoma of stomach
C2011231|giant cell and spindle cell carcinoma of stomach
C2011231|giant cell and spindle cell carcinoma of stomach (diagnosis)
C2142936|pseudosarcomatous carcinoma of stomach
C2142936|pseudosarcomatous carcinoma of stomach (diagnosis)
C2111818|polygonal cell carcinoma of stomach
C2111818|polygonal cell carcinoma of stomach (diagnosis)
C2010505|carcinoma of stomach with osteoclast-like giant cells
C2010505|carcinoma of stomach with osteoclast-like giant cells (diagnosis)
C2010505|gastric carcinoma with osteoclast-like giant cells
C2033236|papillary carcinoma of stomach (diagnosis)
C2033236|papillary carcinoma of stomach
C2189366|verrucous carcinoma of stomach
C2189366|verrucous carcinoma of stomach (diagnosis)
C2010501|diffuse carcinoma of stomach (diagnosis)
C2010501|diffuse carcinoma of stomach
C2010503|parietal cell carcinoma of stomach (diagnosis)
C2010503|parietal cell carcinoma of stomach
C2017458|solid carcinoma of stomach
C2017458|solid carcinoma of stomach (diagnosis)
C2010504|carcinoma simplex of stomach (diagnosis)
C2010504|carcinoma simplex of stomach
C2010502|neuroendocrine carcinoma of stomach (diagnosis)
C2010502|neuroendocrine carcinoma of stomach
C2204850|medullary carcinoma of stomach
C2204850|medullary carcinoma of stomach (diagnosis)
C2204851|epithelial-myoepithelial carcinoma of stomach (diagnosis)
C2204851|epithelial-myoepithelial carcinoma of stomach
C2064167|signet ring cell carcinoma of stomach
C2064167|signet ring cell carcinoma of stomach (diagnosis)
C2064167|gastric signet ring cell carcinoma
C1333761|adenosquamous carcinoma of stomach (diagnosis)
C1333761|adenosquamous carcinoma of stomach
C1333761|gastric adenosquamous carcinoma
C1333761|Adenosquamous Carcinoma of the Stomach
C1333789|squamous cell carcinoma of stomach (diagnosis)
C1333789|squamous cell carcinoma of stomach
C1333789|Gastric Squamous Cell Carcinoma
C1333789|Squamous Cell Carcinoma of the Stomach
C1333788|small cell carcinoma of stomach (diagnosis)
C1333788|small cell carcinoma of stomach
C1333788|gastric small cell carcinoma
C1333788|Gastric Small Cell Neuroendocrine Carcinoma
C1333788|Oat Cell Carcinoma of Stomach
C1333788|Gastric Oat Cell Carcinoma
C1333788|Oat Cell Carcinoma of the Stomach
C1333788|Small Cell Carcinoma of the Stomach
C2983703|Gastric Carcinoma by AJCC v6 Stage
C2984086|Gastric Carcinoma by AJCC v7 Stage
C3272409|Gastric Neuroendocrine Carcinoma
C3272409|Gastric NEC
C3272411|Gastric Mixed Adenoneuroendocrine Carcinoma
C3272411|Gastric MANEC
C0345804|gastric malignant carcinoma body
C0345804|Carcinoma of body of stomach (diagnosis)
C0345804|Carcinoma of body of stomach
C0345804|Carcinoma of body of stomach (disorder)
C0345804|Gastric Body Cancer
C0345804|Gastric Body Carcinoma
C0345804|Cancer of Body of Stomach
C0345804|Cancer of Gastric Body
C0345804|Cancer of the Body of the Stomach
C0345804|Cancer of the Gastric Body
C0345804|Carcinoma of Gastric Body
C0345804|Carcinoma of the Body of the Stomach
C0345804|Carcinoma of the Gastric Body
C0345814|gastric malignant carcinoma pylorus
C0345814|Carcinoma of pylorus (diagnosis)
C0345814|Carcinoma of pylorus
C0345814|Pyloric carcinoma
C0345814|Carcinoma of pylorus (disorder)
C0345809|gastric malignant carcinoma pyloric antrum
C0345809|Carcinoma of pyloric antrum
C0345809|Carcinoma of pyloric antrum (diagnosis)
C0345809|Carcinoma of pyloric antrum (disorder)
C0345794|gastric malignant carcinoma cardia
C0345794|Carcinoma of cardia
C0345794|Carcinoma of cardia (diagnosis)
C0345794|Carcinoma of cardia (disorder)
C0345799|Carcinoma of fundus of stomach
C0345799|Carcinoma of fundus of stomach (diagnosis)
C0345799|gastric malignant carcinoma fundus
C0345799|Carcinoma of fundus of stomach (disorder)
C0345799|Gastric Fundus Cancer
C0345799|Gastric Fundus Carcinoma
C0345799|Cancer of Fundus of Stomach
C0345799|Cancer of Gastric Fundus
C0345799|Cancer of the Fundus of the Stomach
C0345799|Cancer of the Gastric Fundus
C0345799|Carcinoma of Gastric Fundus
C0345799|Carcinoma of the Fundus of the Stomach
C0345799|Carcinoma of the Gastric Fundus
C0740488|gastric malignant carcinoma greater curve
C0740488|Carcinoma of greater curve of stomach (diagnosis)
C0740488|Carcinoma of greater curve of stomach
C0740488|Carcinoma of greater curve of stomach (disorder)
C0349530|Early gastric cancer
C0349530|gastric neoplasm malignant early cancer
C0349530|Early gastric cancer (diagnosis)
C0349530|EGC - Early gastric cancer
C0349530|Early gastric cancer (disorder)
C0349530|EGC
C0349530|Microinvasive Gastric Cancer
C0349530|Superficial Gastric Cancer
C0349530|Superficial Spreading Gastric Cancer
C0349530|Surface Gastric Cancer
C0349531|Late gastric cancer (diagnosis)
C0349531|Late gastric cancer
C0349531|gastric neoplasm malignant late cancer
C0349531|LGC - Late gastric cancer
C0349531|Late gastric cancer (disorder)
C3899661|Childhood Gastric Carcinoma
C0280253|stage, gastric cancer
C0280253|gastric cancer stage
C0280253|stomach cancer stage
C0279889|cellular diagnosis, gastric cancer
C0279889|gastric cancer cellular diagnosis
C0279889|stomach cancer cellular diagnosis
C1333763|Gastric Cardia Cancer
C1333763|Gastric Cardia Carcinoma
C1333763|Cancer of Gastric Cardia
C1333763|Cancer of the Gastric Cardia
C1333763|Carcinoma of Cardia of Stomach
C1333763|Carcinoma of Gastric Cardia
C1333763|Carcinoma of the Cardia of the Stomach
C1333763|Carcinoma of the Gastric Cardia
C0278502|Gastric cancer recurrent
C0278502|Recurrent Gastric Carcinoma
C0278502|Recurrent Gastric Cancer
C0278502|Stomach cancer recurrent
C0278502|Gastric carcinoma recurrent
C0278502|Stomach carcinoma recurrent
C0278502|gastric cancer, recurrent
C0278502|stomach cancer, recurrent
C0278502|Gastric Carcinoma, Recurrent
C0278502|Recurrent Cancer of Stomach
C0278502|Recurrent Cancer of the Stomach
C0278502|Recurrent Carcinoma of Stomach
C0278502|Recurrent Carcinoma of the Stomach
C0278502|Recurrent Stomach Cancer
C0278502|Recurrent Stomach Carcinoma
C1333787|Gastric Pylorus Cancer
C1333787|Gastric Pylorus Carcinoma
C1333787|Cancer of Gastric Pylorus
C1333787|Cancer of Pylorus of Stomach
C1333787|Cancer of the Gastric Pylorus
C1333787|Cancer of the Pylorus of the Stomach
C1333787|Carcinoma of Gastric Pylorus
C1333787|Carcinoma of Pylorus of Stomach
C1333787|Carcinoma of the Gastric Pylorus
C1333787|Carcinoma of the Pylorus of the Stomach
C0278701|Gastric adenocarcinoma
C0278701|adenocarcinoma of stomach
C0278701|adenocarcinoma of stomach (diagnosis)
C0278701|Adenocarcinoma gastric
C0278701|Adenocarcinoma - stomach
C0278701|Adenocarcinoma of the stomach
C0278701|Cancer of stomach, adenocarcinoma
C0278701|Adenocarcinoma of stomach (disorder)
C0278701|gastric cancer, adenocarcinoma
C0278701|stomach cancer, adenocarcinoma
C0278701|stomach, adenocarcinoma of the
C0278701|Stomach Adenocarcinoma
C0809960|Cancer of rectum and anus
C0809962|Cancer of other GI organs; peritoneum
