# tui|tui|txt
C0013862||PAGE|
C0013862||page|
C0013862||page Polyacrylamide Gel Electrophoresis|
C0065374||Lysinopril|medication
# C3536832||Air|physical_exam # JIRA/BIOMED-377
C1321899||paste|
C0001975||Alcohol|social
C0020517||ALLERGIES|
C0013227||General drug type|
C0010294||creatinine|lab
C0032825||Potassium Chloride|lab
C0012634||Disease|
C0039082||Syndrome|
C0001457||ADA|
C3811629||ADA|
C0201931||pCO2|lab
C0202155||pO2|lab
C0032952||Prednisone|medication
# C0065374||lisinopril| # JIRA/BIOMED-265
C0032821||Potassium|lab
C0596019||chloride|lab
C0373675||Magnesium|
C3811652||April|
C0022885||Test|
C1266240||pg|
C1442775||if|
C1441488||Auto|
C0406810||NAME|
C0009905||pill|
C0489531||Allergies|
C3539909||Allergies|
C0449416||Source|
C2825142||Results|
C1873497||Normal|
C1413137||CAST|
C1868670||Other|
C0518766||Vital Signs|
C0311392||Sign|
C0277814||Sitting|
C3714536||Social History|
C2004062||History|
C0270724||Plan|
C1273518||Responsible|
# C0006675||Calcium|lab # JIRA/BIOMED-373
C0311392||signed|
C0421451||DOB|
C3812881||Author|
C3160715||Mixed|
C1301526||Clare|
C2919019||severe|
C1272751||does|
C0424101||innattention|
C1299585||does not|
C1299586||difficulty|
C1416798||large|
C0449255||context|
C3541994||dressed|
CN235300||delayed|
C0178539||cellular|
C2700258||volume|
C1441613||ID|
C0037813||ms|
C1880121||color|
C2827757||resistant|
C0947630||study|
C3272888||clarity|
C1979963||profile|
C2362103||computer assisted|
C4049938||activity|
C0085672||MICRO|
C0002778||ANALYSIS|
C1328856||CHIP|
C4050322||MAP|
C2827755||intermediate|
C1299487||Patient name|
C0455458||Past medical history|
C2676739||glass|
C1254351||drugs|
C1299586||difficulty|
C2826292||scan|
C1416798||large|
C0460139||pressure|
C0442739||unchange|
C2699517||ABSENT|
C3542022||SOFT|
C0039225||Tablet|
C0006935||Capsule|
C0994475||Pill|
C0041942||Urea|lab
C0028158||Nitrogen|lab
# C0017725||Glucose|lab # JIRA/BIOMED-372
# C0024467||Magnesium|  # JIRA/BIOMED-378
C2931488||not provided|
C0442726||Detected|