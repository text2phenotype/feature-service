C0854086|Social alcohol drinker
C1531491|Alcohol consumption counseling
C0085762|Alcohol abuse
C0551570|History of alcohol use:Finding:Point in time:^Patient:Narrative:Reported
C0560219|Alcohol intake above recommended sensible limits
0679277|alcohol use disorder classification
C0687132|heavy drinking
C0740870|ALCOHOL USE FOR SLEEP
C0740872|social drinking
C1387092|alcohol; harmful use
C1545431|Patient drug or alcohol use
C1976670|Use of alcohol at least weekly
C2136082|alcohol use interfering with school
C2136085|alcohol use causing hazard
C2215686|alcohol use during pregnancy
C2215687|alcohol use interfering with work
C3837075|intervention for alcohol use
C3838370|brief intervention for alcohol use
C3841867|Patient admits to alcohol use
C0001948|Alcohol consumption
C0552479|Alcohol use history
C0038586|Substance Use Disorders
C0001948|Alcohol consumption (SNOMED:160573003)
C0687725|Alcoholics
C0556297|Current drinker
C0337678|Alcoholic beverage heavy drinker
C0552479|Alcohol use history
C0085762|Alcohol abuse
C2215684|alcohol consumption history (history)
C0001956|Alcohol Use Disorder
C0001969|Alcoholic Intoxication
C0001973|Alcoholic Intoxication, Chronic
C0683991|Ex-alcoholic
C0237123|Alcohol or Other Drugs use
C0854086|Social alcohol drinker
C2366975|counseling about risk of alcohol consumption
C2366975|counseling about risk of alcohol consumption (treatment)
C2366975|education performed about risk of alcohol consumption
C1531492|Alcohol counselling by other agencies (procedure)
C1531492|Counselling about alcohol by other agencies
C1531492|Counseling about alcohol by other agencies (procedure)
C1531492|Alcohol counseling by other agencies
C1531492|Alcohol counselling by other agencies
C1531492|Counseling about alcohol by other agencies
C1531492|Alcohol counselling by other agencies (regime/therapy)
C3494740|Alcohol brief intervention
C3494740|Alcohol brief intervention (procedure)
C3165324|Counseling About Alcohol Use
C3165324|Counselling About Alcohol Use
C0418859|Advice on alcohol consumption
C0418859|Advice relating to alcohol consumption
C0418859|Education about alcohol consumption
C0418859|Education about alcohol consumption (procedure)
C0418859|Advice relating to alcohol consumption (procedure)
C0418859|Advice on alcohol consumption (procedure)
C0418859|Advice on alcohol consumption (regime/therapy)
C0085762|Abuse, Alcohol
C0085762|Alcohol abuse
C0085762|alcohol abuse (diagnosis)
C0085762|ethanol abuse
C0085762|ETOH abuse
C0085762|Alcohol abuse-unspec
C0085762|rndx alcohol abuse
C0085762|rndx alcohol abuse (diagnosis)
C0085762|Alcohol abuse, unspecified
C0085762|Alcohol abuse, unspecified drinking behavior
C0085762|Ethanol abuse (finding)
C0085762|Alcohol abuse, unspecified drinking behaviour
C0085762|AA - Alcohol abuse
C0085762|Alcohol abuse (disorder)
C0085762|abuse; alcohol
C0085762|alcohol; abuse
C0085762|problem; alcohol use
C0085762|alcohol; use, problem
C0085762|Problem Drinking
C2874370|Alcohol abuse, uncomplicated
C2874370|alcohol abuse - uncomplicated
C2874370|alcohol abuse - uncomplicated (diagnosis)
C2874371|Alcohol abuse with intoxication
C2874371|Alcohol abuse with intoxication, unspecified
C2874371|alcohol abuse with intoxication (diagnosis)
C2874377|Alcohol abuse with alcohol-induced mood disorder
C2874377|Alcohol abuse with alcohol-induced psychotic disorder, unspecified
C2874377|Alcohol abuse with alcohol-induced psychotic disorder
C2874377|Alcohol abuse with alcohol-induced psychotic disorder, unsp
C2874377|alcohol abuse with alcohol-induced mood disorder (diagnosis)
C2874377|alcohol abuse with alcohol-induced psychotic disorder (diagnosis)
C2874381|Alcohol abuse with other alcohol-induced disorders
C2874381|Alcohol abuse with other alcohol-induced disorder
C2874382|Alcohol abuse with unspecified alcohol-induced disorder
C1812624|Alcohol abuse, continuous drinking behavior
C1812624|continuous alcohol abuse (diagnosis)
C1812624|continuous alcohol abuse
C1812624|continuous ETOH abuse
C1812624|continuous ethanol abuse
C1812624|Alcohol abuse-continuous
C1812624|Alcohol abuse, continuous
C0154515|episodic alcohol abuse
C0154515|episodic alcohol abuse (diagnosis)
C0154515|Alcohol abuse, episodic drinking behavior
C0154515|episodic ethanol abuse
C0154515|episodic ETOH abuse
C0154515|Alcohol abuse-episodic
C0154515|Alcohol abuse, episodic
C0154515|Alcohol abuse, episodic drinking behaviour
C0154516|alcohol abuse in remission
C0154516|alcohol abuse in remission (diagnosis)
C0154516|Alcohol abuse, in remission
C0154516|ETOH abuse in remission
C0154516|ethanol abuse in remission
C0154516|Alcohol abuse-in remiss
C2874372|Alcohol abuse with intoxication, uncomplicated
C2874372|alcohol abuse with intoxication - uncomplicated
C2874372|alcohol abuse with intoxication - uncomplicated (diagnosis)
C2874373|Alcohol abuse with intoxication delirium
C2874373|alcohol abuse with intoxication delirium (diagnosis)
C2874375|Alcohol abuse with alcohol-induced psychotic disorder with delusions
C2874375|Alcohol abuse w alcoh-induce psychotic disorder w delusions
C2874375|alcohol abuse with alcohol-induced psychotic disorder with delusions (diagnosis)
C2874376|Alcohol abuse with alcohol-induced psychotic disorder with hallucinations
C2874376|Alcohol abuse w alcoh-induce psychotic disorder w hallucin
C2874376|alcohol abuse with alcohol-induced psychotic disorder with hallucinations (diagnosis)
C3509160|alcohol abuse with alcohol-induced disorder (diagnosis)
C3509160|alcohol abuse with alcohol-induced disorder
C2874378|Alcohol abuse with alcohol-induced anxiety disorder
C2874378|alcohol abuse with alcohol-induced anxiety disorder (diagnosis)
C2874379|Alcohol abuse with alcohol-induced sexual dysfunction
C2874379|alcohol abuse with alcohol-induced sexual dysfunction (diagnosis)
C2874380|Alcohol abuse with alcohol-induced sleep disorder
C2874380|alcohol abuse with alcohol-induced sleep disorder (diagnosis)
C0338709|Nondependent alcohol abuse
C0338709|Alcohol abuse -non dep.
C0338709|Nondependent alcohol abuse, unspecified (disorder)
C0338709|Nondependent alcohol abuse, unspecified
C0338709|Nondependent alcohol abuse NOS
C0338709|Nondependent alcohol abuse NOS (disorder)
C0338709|Non-dependent abuse of alcohol
C0338709|alcohol abuse nondependent
C0338709|Nondependent alcohol abuse (diagnosis)
C0338709|Nondependent abuse of alcohol
C0338709|Nondependent alcohol abuse (disorder)
C0338709|alcohol; use, harmful (non-dependent)
C0338709|use; alcohol, harmful (non-dependent)
C0001973|Alcoholism
C0001973|Dipsomania
C0001973|Chronic Alcoholic Intoxication
C0001973|Intoxication, Chronic Alcoholic
C0001973|Mental and behavioral disorders due to use of alcohol, dependence syndrome
C0001973|Mental and behavioural disorders due to use of alcohol, dependence syndrome
C0001973|ALCOHOL DEPENDENCE
C0001973|ALCOHOLIC INTOX CHRONIC
C0001973|ETOHism
C0001973|ETOH dependence
C0001973|addicted to alcohol
C0001973|alcohol dependence (diagnosis)
C0001973|Alcoholism [Disease/Finding]
C0001973|Alcoholic Intoxication, Chronic
C0001973|Abuse;alcohol;chronic
C0001973|Addiction;alcohol
C0001973|Intoxication;alcohol;chronic
C0001973|Dependence;alcohol
C0001973|Alcoholism;chronic
C0001973|alcoholism/alcohol abuse
C0001973|Addiction, Alcohol
C0001973|Dependence, Alcohol
C0001973|Unspecified chronic alcoholism (disorder)
C0001973|Alcohol problem drinking
C0001973|[X]Mental and behavioural disorders due to use of alcohol: dependence syndrome
C0001973|Chronic alcoholism (disorder)
C0001973|Alcohol dependence syndrome (& [dipsomania]) (disorder)
C0001973|Chronic alcoholism (& [dipsomania])
C0001973|[X]Mental and behavioral disorders due to use of alcohol: dependence syndrome
C0001973|Chronic alcoholism
C0001973|Alcohol dependence syndrome (& [dipsomania])
C0001973|Alcohol dependence syndrome NOS
C0001973|Chronic alcoholism NOS (disorder)
C0001973|[X]Alcohol addiction
C0001973|Chronic alcoholism NOS
C0001973|[X]Dipsomania
C0001973|(Alcohol dependence syndrome [including alcoholism]) or (alcohol problem drinking) (disorder)
C0001973|Alcohol dependence syndrome
C0001973|Alcohol dependence syndrome NOS (disorder)
C0001973|Chronic alcoholism (& [dipsomania]) (disorder)
C0001973|(Alcohol dependence syndrome [including alcoholism]) or (alcohol problem drinking)
C0001973|Unspecified chronic alcoholism
C0001973|Dipsomania (finding)
C0001973|[X]Mental and behavioral disorders due to use of alcohol: dependence syndrome (disorder)
C0001973|[X]Chronic alcoholism
C0001973|alcohol abuse - persistent
C0001973|alcohol abuse - persistent (diagnosis)
C0001973|Alcohol Addiction
C0001973|Alcohol dependency
C0001973|Alcoholism and Alcohol Abuse
C0001973|Alcohol abuse chronic
C0001973|Alcohol abuse, continuous drinking behaviour
C0001973|Alcohol abuse, continuous drinking behavior
C0001973|Chronic alcohol abuse
C0001973|Persistent alcohol abuse
C0001973|Alcohol dependence (disorder)
C0001973|Alcoholism (disorder)
C0001973|Persistent alcohol abuse (disorder)
C0001973|chronic; drunkenness
C0001973|dependence; alcohol
C0001973|drunkenness; chronic
C0001973|addiction; alcohol
C0001973|alcohol; addiction
C0001973|alcohol; dependence
C0001973|Alcoholism, NOS
C0001973|Chronic alcoholism [Ambiguous]
C0001973|dependence; ethyl alcohol
C0001973|ethyl alcohol; dependence
C0001973|chronic alcohol intoxication
C0349269|Abuse of non-dependence-producing substances
C0349269|[X]Abuse of non-dependence-producing substances
C0349269|Abuse of non-dependence-producing substances (disorder)
C0582513|Methanol abuse
C0582513|Methanol abuse (diagnosis)
C0582513|unspecified psych substance abuse methanol
C0582513|Methanol abuse (disorder)
C0238265|Central demyelination of corpus callosum
C0238265|Marchiafava-Bignami disease
C0238265|Marchiafava Bignami disease
C0238265|Marchiafava Bignami Syndrome
C0238265|central demyelination of corpus callosum (diagnosis)
C0238265|Marchiafava-Bignami disease (diagnosis)
C0238265|Marchiafava-Bignami Syndrome
C0238265|Marchiafava-Bignami Disease [Disease/Finding]
C0238265|Marchiafava disease
C0238265|Marchiafava-Bignami disease (disorder)
C0238265|Central demyelination of corpus callosum (disorder)
C0238265|Marchiafava
C0238265|corpus callosum; demyelination
C0238265|demyelination; corpus callosum
C0238265|encephalopathy; demyelinating callosal
C0556330|Drinks in morning to get rid of hangover
C0556330|Drinks in morning to get rid of hangover (finding)
C0556343|Drinking bout
C0556343|Drinking bout (finding)
C0556383|Feels drinking is out of control
C0556383|Feels drinking is out of control (finding)
C0522172|Feeling drunk
C0522172|Drunkenness feeling of
C0522172|Feeling groggy
C0522172|Feeling intoxicated
C0522172|Feeling intoxicated (finding)
C0556364|Unable to stop drinking before intoxication
C0556364|Unable to stop drinking before intoxication (finding)
C0560219|Excessive alcohol use
C0560219|Alcohol intake above recommended sensible limits
C0560219|Alcohol intake above recommended sensible limits (finding)
C0560219|Excessive alcohol consumption
C0560219|XS - Excessive alcohol consumption
C0560219|XS - Excessive ethanol consumption
C0560219|Excessive ethanol consumption
C0560219|Excessive drinking of alcohol NOS
C0556337|Alcoholic binges exceeding safe amounts
C0556337|Alcoholic binges exceeding safe amounts (finding)
C0556336|Alcoholic binges exceeding sensible amounts
C0556336|Alcoholic binges exceeding sensible amounts (finding)
C0556346|Binge drinking
C0556346|Drinking, Binge
C0556346|Binge Drinking [Disease/Finding]
C0556346|Alcohol binge
C0556346|Drinking binge
C0556346|Drinking binge (finding)
C0556335|Binge drinker
C0556335|Bout drinker
C0556335|Episodic drinker
C0556335|Binge drinker (finding)
C0556363|Unable to control spontaneous drinking bouts
C0556363|Unable to control spontaneous drinking bouts (finding)
C2106524|combined drug and alcohol abuse (diagnosis)
C2106524|combined drug and alcohol abuse
C0551570|History of alcohol use:Finding:Point in time:^Patient:Narrative:Reported
C0551570|History of alcohol use:Find:Pt:^Patient:Nar:Reported
C0551570|Alcohol use Hx Reported
C0551570|History of alcohol use Narrative
C2181572|a breathalyzer for blood alcohol content showed an excessive blood alcohol level
C2181572|breathalyzer for blood alcohol content excessive blood alcohol level
C2181572|breathalyzer for blood alcohol content: excessive blood alcohol level (lab test)
C2181572|breathalyzer for blood alcohol content: excessive blood alcohol level
C1387092|harmful; use, alcohol
C1387092|alcohol; harmful use
C2136086|alcohol use causing hazard at work (history)
C2136086|alcohol use causing hazard at work
C2136087|alcohol use causing hazard while driving
C2136087|alcohol use causing hazard while driving (history)
C1959897|Alcohol consumption during pregnancy
C1959897|Alcohol consumption during pregnancy (finding)
C3838370|brief intervention for alcohol use (treatment)
C3838370|brief intervention for alcohol use
C3838370|intervention for alcohol use brief
C0001948|ALCOHOL USE
C0001948|Alcohol Drinking
C0001948|Consumption, Alcohol
C0001948|alcoholic beverage consumption
C0001948|Alcohol consumption
C0001948|drinking alcohol
C0001948|Alcohol product use
C0001948|Drinking
C0001948|alcohol use (diagnosis)
C0001948|Alcohol consumption NOS
C0001948|Alcohol intake (observable entity)
C0001948|Alcohol consumption NOS (observable entity)
C0001948|Alcohol intake
C0001948|Alcohol consumption NOS (finding)
C0001948|Drinking, Alcohol
C0001948|AI - Alcohol intake
C0001948|ETOH - Alcohol intake
C0001948|Alcoholic drink intake
C0001948|Ethanol intake
C0001948|alcohol; use
C0001948|use; alcohol
C0001948|Drinking (Alcohol)
C0854087|Abstains from alcohol
C0687725|Alcoholic
C0687725|Alcoholics
C0687725|Boozer
C0687725|Dependent drinker
C0687725|Problem drinker
C0687725|Problem drinker (finding)
C0687725|Problem drinker (life style)
C1698582|Maternal alcohol use
C0683991|Ex-alcoholic
C0001962|Alcohol
C0001962|Ethanol
C0001962|Ethyl Alcohol
C0001962|Alcohol, Grain
C0001962|ETOH
C0001962|Absolute Ethanol
C0001962|Methylcarbinol
C0001962|ALCOHOL,ETHYL
C0001962|Alcohol, Ethyl
C0001962|Grain Alcohol
C0001962|Ethanol [Chemical/Ingredient]
C0001962|EtOH - Alcohol
C0001962|Ethyl alcohol (substance)
C0001962|Drinking alcohol
C0001962|EtOH - Ethanol
C0001962|Ethyl alcohol (product)
C0001962|Alcohol (Grain)
C0556297|Current drinker of alcohol
C0556297|Alcoholic beverage drinker
C0556297|Current drinker
C0556297|Alcohol user
C0556297|Drinks alcohol
C0556297|Current drinker of alcohol (finding)
C0556297|Alcoholic beverage drinker, NOS
C0556297|Current drinker (life style)
C3650363|alcohol use with alcohol-induced disorder (diagnosis)
C3650363|alcohol use with alcohol-induced disorder
C4042862|Drinking, College
C4042862|Alcohol Drinking in College
C4042862|Student Drinking, College
C4042862|Student Drinking, University
C4042862|Alcohol Drinking, College Students
C4042862|College Drinking
C4042862|College Student Drinking
C4042862|University Student Drinking
C0684314|Teenage Drinking
C0684314|Underage Drinking
C0684314|Drinking, Teen
C0684314|Alcohol Consumption, Adolescent
C0684314|Alcohol Consumption, Youth
C0684314|Drinking, Teenage
C0684314|Drinking, Adolescent
C0684314|Alcohol Use, Underage
C0684314|Alcohol Use, Adolescent
C0684314|Drinking, Underage
C0684314|Drinking, Youth
C0684314|Alcohol Consumption, Underage
C0684314|Underage Alcohol Use
C0684314|Adolescent Alcohol Use
C0684314|Youth Alcohol Consumption
C0684314|Youth Drinking
C0684314|Underage Alcohol Consumption
C0684314|Adolescent Drinking
C0684314|Teen Drinking
C0684314|Adolescent Alcohol Consumption
C0559430|Beer intake
C0559430|Beer intake (observable entity)
C0559433|Spirits intake (observable entity)
C0559433|Hard liquor intake (observable entity)
C0559433|hard liquor consumption (history)
C0559433|hard liquor consumption
C0559433|Spirits intake
C0559433|Hard liquor intake
C0559432|Wine intake
C0559432|Wine intake (observable entity)
C2114426|previous attempts to decrease alcohol consumption (history)
C2114426|previous attempts to decrease alcohol consumption
C2030272|heavy alcohol consumption
C2030272|heavy alcohol consumption (history)
C2133669|alcohol consumption within last 12 hours (history)
C2133669|alcohol consumption within last 12 hours
C2133669|alcohol consumption within the last 12 hours
C2136008|drinking in moderation (two drinks/day or fewer) (history)
C2136008|drinking in moderation (two drinks/day or fewer)
C2136008|drinking in moderation (2 drinks / day or fewer)
C2136008|drinking in moderation (2 drinks/day or fewer)
C2048467|inability to further reduce amount of alcohol (history)
C2048467|inability to further reduce amount of alcohol
C2048467|inability to further reduce amount of alcohol consumed
C2048484|inability to quit drinking alcohol (history)
C2048484|inability to quit drinking alcohol
C2136082|alcohol use interfering with school
C2136082|alcohol use interfering with school (history)
C2136083|alcohol use disrupting home environment
C2136083|alcohol use disrupting home environment (history)
C2136084|alcohol use causing legal problems
C2136084|alcohol use causing legal problems (history)
C2136085|alcohol use causing hazard (history)
C2136085|alcohol use causing hazard
C2136088|alcohol use consumes much time (history)
C2136088|alcohol use consumes much time
C2136092|alcohol use results in reduced important activities (history)
C2136092|alcohol use results in reduced important activities
C2136111|drinking more and for longer periods than intended
C2136111|drinking alcohol more and for longer periods than intended (history)
C2136111|drinking alcohol more and for longer periods than intended
C2136112|alcohol use continues despite knowledge of harmful effects
C2136112|alcohol use continues despite knowledge of harmful effects (history)
C2163372|current drinking being denied but suspected (history)
C2163372|current drinking being denied but suspected
C2163372|suspected covert drinking
C2215685|alcohol use affecting relationships with others (history)
C2215685|alcohol use affecting relationships with others
C2215687|alcohol use interfering with work (history)
C2215687|alcohol use interfering with work
C2199079|drinking more alcohol than friends or associates (history)
C2199079|drinking more alcohol than friends or associates
C2029398|having drink of alcohol in morning to get going
C2029398|having drink of alcohol in morning to get going (history)
C2199076|drinking alcohol frequently before age 18
C2199076|drinking alcohol frequently before age 18 (history)
C2199076|drinking alcohol frequently before the age of 18
C2107808|beer consumption (history)
C2107808|beer consumption
C2107808|consumption of beer (history)
C2107808|consumption of beer
C2203276|wine consumption (history)
C2203276|wine consumption
C2220425|History of being a social drinker
C2220425|social drinker (history)
C2220425|social drinker
C2220425|being a social drinker
C2220425|a social drinker
C2048464|inability to control amount of alcohol consumed
C2048464|inability to control amount of alcohol consumed (history)
C2107728|considered quitting drinking alcohol (history)
C2107728|considered quitting drinking alcohol
C2107728|having considered quitting drinking
C2011202|getting angry when talked to about drinking
C2011202|getting angry when talked to about drinking (history)
C2199077|drinking alcohol regularly and feeling guilty about it (history)
C2199077|drinking alcohol regularly, feeling guilty about it
C2199077|drinking alcohol regularly and feeling guilty about it
C2165493|denying that drinking is causing problems
C2165493|denying that drinking is causing problems (history)
C2220520|behavior changes after small amounts of alcohol (history)
C2220520|behavior changes after small amounts of alcohol
C2215683|alcohol consumption cut within last 48 hours (history)
C2215683|alcohol consumption cut within last 48 hours
C2215683|alcohol consumption was cut within the last 48 hours
C2169567|recent increase in alcohol consumption (history)
C2169567|recent increase in alcohol consumption
C2169538|recent decrease in alcohol consumption
C2169538|recent decrease in alcohol consumption (history)
C0038587|Substance Withdrawal Syndrome
C0038587|Substance Withdrawal Syndromes
C0038587|Syndrome, Substance Withdrawal
C0038587|Syndromes, Substance Withdrawal
C0038587|Withdrawal Syndrome, Substance
C0038587|Withdrawal Syndromes, Substance
C0038587|Withdrawal syndrome
C0038587|Substance Withdrawal Syndrome [Disease/Finding]
C0038587|Drug Withdrawal
C0038587|Syndrome withdrawal
C1510472|Dependence, Drug
C1510472|DRUG DEPENDENCE
C1510472|Drug Dependency
C1510472|drug addiction
C1510472|drug dependence (diagnosis)
C1510472|Addiction, Drug
C1510472|Addiction any drug
C1510472|Abuse;drug(s);dependent
C1510472|Addiction;drug(s)
C1510472|Dependence;drug(s)
C1510472|Drug dependence NOS
C1510472|Dependence syndrome (disorder)
C1510472|Drug dependence NOS (disorder)
C1510472|[X]Drug addiction NOS
C1510472|Dependence syndrome
C1510472|substance abuse drug dependent
C1510472|Dependent drug abuse
C1510472|Dependent drug abuse (diagnosis)
C1510472|Unspecified drug dependence
C1510472|Drug dependence, unspecified
C1510472|Addiction to drugs
C1510472|Dependence drug (NOS)
C1510472|Dependent drug abuse (disorder)
C1510472|Drug dependence (disorder)
C1510472|Psychoactive substance dependence (disorder)
C1510472|Psychoactive substance dependence
C1510472|dependence; drugs
C1510472|dependence; drug
C1510472|dependence; substance
C1510472|drug; dependence
C1510472|drugs; dependence
C1510472|Psychoactive substance dependence, NOS
C1510472|Drug dependence, NOS
C1510472|Dependency (Drug)
C1510472|Chemical Dependence
C1510472|Drug addiction NOS
C1510472|drug abuse and dependency
C0679272|polydrug abuse
C0679272|multidrug abuse
C0700319|Mentally ill chemical abuse
C0700319|MICA
C0013222|Disorder, Drug Use
C0013222|Drug Use Disorder
C0013222|DRUG USE DIS
C0013222|drug use disorders (diagnosis)
C0013222|drug use disorders
C0017782|Glue Sniffing (inhalant abuse)
C0017782|Abuses, Glue
C0017782|Glue Abuses
C0017782|Abuse, Glue
C0017782|Glue Sniffing
C0017782|Glue Sniffings
C0017782|Abuse;drug(s);glue
C0017782|Glue Abuse
C0017782|glue; sniffing
C0017782|sniffing; glue
C0033882|Psychoactive substance use disorder (disorder)
C0033882|Psychoactive substance use disorder
C0033882|Psychoactive substance use disorder, NOS
C2919052|Alcohol or other drugs dependence
C3665355|drug-induced disorder
C3665355|drug-induced disorder (diagnosis)
C0236664|Alcohol Related Disorders
C0236664|Alcohol-Related Disorder
C0236664|Alcohol-Related Disorders
C0236664|Disorder, Alcohol-Related
C0236664|Disorders, Alcohol-Related
C0236664|ALCOHOL RELATED DIS
C0236664|Alcohol-Related Disorders [Disease/Finding]
C0236664|alcohol-related disorders (diagnosis)
C0236664|alcohol disorders
C0236664|Alcohol-induced organic mental disorder (disorder)
C0236664|Alcohol-induced organic mental disorder
C0236664|Alcohol-induced organic mental disorder, NOS
C0236664|Alcohol-related disorder, NOS
C0236664|Alcohol-related disorder NOS
C0236734|caffeine-related disorders
C0236734|caffeine-related disorders (diagnosis)
C0236734|Caffeine-related disorder (disorder)
C0236734|Caffeine-related disorder
C0236734|Caffeine-related disorder, NOS
C0236738|inhalant-related disorders (diagnosis)
C0236738|inhalant-related disorders
C0236738|Inhalant related disorders
C0236738|Inhalant induced mental disorder
C0236738|Inhalant-induced organic mental disorder (disorder)
C0236738|Inhalant-induced organic mental disorder
C0236738|Inhalant-related disorder
C0236738|Inhalant-induced organic mental disorder, NOS
C0236738|Inhalant-related disorder, NOS
C0376384|Disorder, Nicotine Use
C0376384|Nicotine Use Disorders
C0376384|Use Disorder, Nicotine
C0376384|NICOTINE USE DIS
C0376384|nicotine-related disorders (diagnosis)
C0376384|nicotine-related disorders
C0376384|Nicotine induced mental disorder
C0376384|Nicotine-induced organic mental disorder (disorder)
C0376384|Nicotine-induced organic mental disorder
C0376384|Nicotine-related disorder
C0376384|Nicotine-induced organic mental disorder, NOS
C0376384|Nicotine-related disorder, NOS
C0376384|Nicotine Use Disorder
C2063802|unspecified substance disorders (diagnosis)
C2063802|unspecified substance disorders
C0038586|SUBSTANCE USE DISORDER
C0038586|Disorder, Substance Use
C0038586|SUBSTANCE USE DIS
C0038586|substance use disorders (diagnosis)
C0038586|substance use disorders
C0740858|Abuse, Substance
C0740858|Abuses, Substance
C0740858|Substance abuse
C0740858|Substance Abuses
C0740858|Substance abuse problem
C0740858|rndx substance abuse
C0740858|rndx substance abuse (diagnosis)
C0740858|Substance Abuse Problems
C0740858|substance abuse (diagnosis)
C0740858|Harmful substance use (disorder)
C0740858|Harmful substance use
C0740858|Nondependent abuse of substance
C0740858|Substance abuse (disorder)
C0740858|disorder, substance abuse
C0740858|substance abuse disorder
C0037263|Alcoholic, Skid Row
C0037263|Alcoholics, Skid Row
C0037263|Skid Row Alcoholics
C0037263|Skid Row Alcoholic
C2960643|Drinks alcoholic cider
C2960643|Drinks alcoholic cider (finding)
C0552479|alcohol use (history)
C0552479|ETOH use
C0552479|alcohol use
C0552479|Alcohol Use History
C0552479|History of alcohol use
C0425331|Drinks beer and hard liquor (finding)
C0425331|Drinks beer and spirits (finding)
C0425331|Drinks beer and spirits
C0425331|Drinks beer and spirits (life style)
C0425331|Drinks beer and hard liquor
C4065069|first alcohol use (history)
C4065069|first alcohol use
C0337678|Alcoholic beverage heavy drinker
C0337678|Heavy drinker (finding)
C0337678|Heavy drinker
C0337678|Drunk
C0337678|Drinks heavily
C0337678|Heavy drinker (life style)
C0337677|Alcoholic beverage moderate drinker
C0337677|Moderate drinker (finding)
C0337677|Moderate drinker
C0337677|Moderate drinker (life style)
C0337676|Alcoholic beverage mild drinker
C0337676|Social drinker
C0337676|Social drinker (finding)
C0337676|Social drinker (life style)
C0425330|Beer drinker (finding)
C0425330|Beer drinker
C0425330|Beer drinker (life style)
C0425332|Drinks wine (finding)
C0425332|Drinks wine
C0425332|Drinks wine (life style)
C0425329|Spirit drinker (finding)
C0425329|Drinker of hard liquor (finding)
C0425329|Spirit drinker
C0425329|Spirit drinker (life style)
C0425329|Drinker of hard liquor
C0556300|Fairly heavy drinker
C0556300|Fairly heavy drinker (finding)
C0556300|Fairly heavy drinker (life style)
C0556301|Very heavy drinker
C0556301|Very heavy drinker (finding)
C0556301|Very heavy drinker (life style)
C0556299|Light drinker (finding)
C0556299|Light drinker
C0556299|Light drinker (life style)
C0556298|Drinks occasionally
C0556298|Drinks on special occasions
C0556298|Occasional drinker
C0556298|Occasional drinker (finding)
C0556298|Occasional drinker (life style)
C0425319|Heavy drinker - 7-9u/day
C0425319|Heavy drinker - 7-9u/day (finding)
C0425319|Heavy drinker - 7-9u/day (life style)
C2242867|recovering alcoholic
C2242867|recovering alcoholic (history)
C2136009|never drank alcohol
C2136009|never drank alcohol (history)
C0425321|stopped drinking alcohol
C0425321|stopped drinking alcohol (history)
C0425321|having stopped drinking alcohol
C0425321|Stopped drinking alcohol (finding)
C0425321|Stopped drinking alcohol (life style)
C3249902|audit alcohol use disorders identification test ___(0-40)
C3249902|audit alcohol use disorders identification test ___(0-40) (history)
C3249903|raps rapid alcohol problems screen ___(0-4)
C3249903|raps rapid alcohol problems screen ___(0-4) (history)
C3249904|ciwa-ar clinical institute withdrawal of alcohol scale ___(0-42) (history)
C3249904|ciwa-ar clinical institute withdrawal of alcohol scale ___(0-42)
C3249901|cage screening test for alcohol dependence ___(0-4)
C3249901|cage screening test for alcohol dependence ___(0-4) (history)
C0496556|Mild alcohol intoxication
C0496557|Moderate alcohol intoxication
C0496558|Severe alcohol intoxication
C0496559|Very severe alcohol intoxication
C0812429|Acute alcoholic intoxication in alcoholism
C0812429|Ac alcohol intox-unspec
C0812429|Acute drunkenness (in alcoholism)
C0812429|Acute alcoholic intoxication in alcoholism, unspecified
C0812429|Acute alcoholic intoxication in alcoholism, unspecified drinking behavior
C0812429|Acute alcoholic intoxication, unspecified, in alcoholism
C0812429|Acute alcoholic intoxication, unspecified, in alcoholism (disorder)
C0812429|Acute alcoholic intoxication in alcoholism NOS
C0812429|Acute alcoholic intoxication in alcoholism NOS (disorder)
C0812429|acute alcohol intoxication in alcoholism
C0812429|alcohol intoxication - acute in alcoholism
C0812429|acute alcohol intoxication in alcoholism (diagnosis)
C0812429|Acute alcoholic intoxication in alcoholism, unspecified drinking behaviour
C0812429|Alcohol dependence with acute alcoholic intoxication
C0812429|Acute alcoholic intoxication in alcoholism (disorder)
C0812429|drunkenness; acute in alcoholism
C0812429|acute; drunkenness in alcoholism
C0812429|Acute alcoholic intoxication, unspecified drinking behavior
C0812429|Acute drunkenness in alcoholism
C0394996|Acute alcoholic intoxication
C0394996|Mental and behavioral disorders due to use of alcohol, acute intoxication
C0394996|Mental and behavioural disorders due to use of alcohol, acute intoxication
C0394996|Intoxication;alcohol;acute
C0394996|[X]Mental and behavioural disorders due to use of alcohol: acute intoxication
C0394996|[X]Mental and behavioral disorders due to use of alcohol: acute intoxication (disorder)
C0394996|[X]Mental and behavioral disorders due to use of alcohol: acute intoxication
C0394996|Alcohol intoxication acute
C0394996|Alcohol intoxication, acute
C0394996|Acute alcohol intoxication
C0001950|Idiosyncratic alcohol intoxication
C0001950|alcohol idiosyncratic intoxication (diagnosis)
C0001950|alcohol idiosyncratic intoxication
C0001950|Pathologic alcohol intox
C0001950|alcohol intoxication - pathological (diagnosis)
C0001950|alcohol intoxication - pathological
C0001950|Pathological alcohol intoxication
C0001950|Pathological drunkenness
C0001950|Pathological intoxication
C0001950|Extreme sensitivity to alcohol syndrome
C0001950|Idiosyncratic intoxication
C0001950|Drunkenness - pathological
C0001950|Idiosyncratic intoxication (disorder)
C0001950|Pathological alcohol intoxication (disorder)
C0001950|drunkenness; pathological
C0001950|intoxication; alcohol, idiosyncratic
C0001950|intoxication; alcohol, pathological
C0001950|intoxication; pathologic
C0001950|pathologic; intoxication
C0001950|pathological; drunkenness
C0001950|alcohol; intoxication, idiosyncratic
C0001950|alcohol; intoxication, pathological
C0001950|Pathologic alcohol intoxication
C0001950|Pathologic drunkenness
C0001969|Alcoholic Intoxication
C0001969|Alcohol Intoxication
C0001969|Drunk
C0001969|INTOX ALCOHOLIC
C0001969|ALCOHOLIC INTOX
C0001969|alcohol intoxication (diagnosis)
C0001969|Drunkennesses
C0001969|Intoxication, Alcoholic
C0001969|Alcoholic Intoxication [Disease/Finding]
C0001969|Drunkenness
C0001969|Abuse;alcohol;acute
C0001969|Intoxication - alcohol
C0001969|Drunkenness NOS
C0001969|Inebriety NOS
C0001969|Inebriety NOS (disorder)
C0001969|Drunkenness NOS (disorder)
C0001969|Alcohol intoxication (disorder)
C0001969|inebriety
C0001969|intoxication; alcohol
C0001969|alcohol; intoxication
C0001969|Intoxication (Alcohol)
C0001969|Addiction;alcohol;acute
C2104528|continuous alcohol intoxication (diagnosis)
C2104528|continuous alcohol intoxication
C2104529|episodic alcohol intoxication
C2104529|episodic alcohol intoxication (diagnosis)
C2104530|alcohol intoxication in remission (diagnosis)
C2104530|alcohol intoxication in remission
C3650362|alcohol intoxication - uncomplicated
C3650362|alcohol use with intoxication - uncomplicated (diagnosis)
C3650362|alcohol use with intoxication - uncomplicated
C0236654|alcohol intoxication delirium
C0236654|alcohol intoxication delirium (diagnosis)
C0236654|Alcohol intoxication delirium (disorder)
C0236654|intoxication; alcohol, delirium
C0236654|alcohol; delirium, intoxication
C0236654|alcohol; intoxication, delirium
C0393756|Hangover from alcohol
C0393756|Alcoholic hangover
C0393756|Hangover (alcohol)
C0393756|Hangover alcoholic
C0393756|Hangover
C0393756|Hangover effect
C0393756|Hangover (finding)
C0393756|Hangover, alcohol
C0033936|Psychoses, Alcoholic
C0033936|Alcoholic psychoses
C0033936|alcoholic psychosis
C0033936|Mental and behavioral disorders due to use of alcohol, psychotic disorder
C0033936|Mental and behavioural disorders due to use of alcohol, psychotic disorder
C0033936|alcohol-induced psychotic disorder
C0033936|alcohol-induced psychotic disorder (diagnosis)
C0033936|Alcohol mental disor NOS
C0033936|Psychoses, Alcoholic [Disease/Finding]
C0033936|Psychosis;alcoholic
C0033936|Alcohol induced psychosis
C0033936|[X]Alcoholic psychosis NOS
C0033936|Alcoholic psychoses (disorder)
C0033936|[X]Mental and behavioral disorders due to use of alcohol: psychotic disorder
C0033936|[X]Mental and behavioural disorders due to use of alcohol: psychotic disorder
C0033936|Alcoholic psychosis NOS
C0033936|Alcoholic psychosis NOS (disorder)
C0033936|[X]Mental and behavioral disorders due to use of alcohol: psychotic disorder (disorder)
C0033936|Alcoholic psychosis, unspecified
C0033936|Unspecified alcoholic psychosis
C0033936|Psychosis alcoholic
C0033936|Alcohol-induced psychosis (disorder)
C0033936|Alcohol-induced psychosis
C0033936|disorder; psychotic, alcohol (due to), alcoholic
C0033936|alcoholism; psychosis
C0033936|psychosis; alcoholic
C0033936|psychotic; disorder, alcohol (due to), alcoholic
C0033936|Alcohol-induced psychosis, NOS
C0033936|Alcoholic psychosis, NOS
C0033936|Alcoholism with psychosis
C0033936|Unspecified alcohol-induced mental disorders
C0392621|methanol poisoning
C0392621|poisoning by methyl alcohol
C0392621|poisoning by methyl alcohol (diagnosis)
C0392621|Methyl alcohol poisoning
C0556374|alcohol influenced driving
C0556374|drunk driving
C0556374|driving while intoxicated
C0556374|Drink driving
C0556374|Drunk driving (finding)
C0556374|Drink driving (finding)
C0338785|alcohol dependence with continuous drinking behavior
C0338785|alcohol dependence with continuous drinking behavior (diagnosis)
C0338785|Continuous chronic alcoholism
C0338785|Continuous chronic alcoholism (disorder)
C2874383|Alcohol dependence, uncomplicated
C2874383|alcohol dependence uncomplicated (diagnosis)
C2874383|alcohol dependence uncomplicated
C2197979|alcohol dependence in remission (diagnosis)
C2197979|alcohol dependence in remission
C2197979|Alcohol dependence, in remission
C2874387|Alcohol dependence with intoxication
C2874387|Alcohol dependence with intoxication, unspecified
C2874387|alcohol dependence with intoxication (diagnosis)
C2874392|Alcohol dependence with withdrawal
C2874392|Alcohol dependence with withdrawal, unspecified
C2874392|alcohol dependence with withdrawal (diagnosis)
C2874393|Alcohol dependence with alcohol-induced mood disorder
C2874393|alcohol dependence with alcohol-induced mood disorder (diagnosis)
C2874397|Alcohol dependence with alcohol-induced psychotic disorder
C2874397|Alcohol dependence with alcohol-induced psychotic disorder, unspecified
C2874397|Alcohol dependence w alcoh-induce psychotic disorder, unsp
C2874397|alcohol dependence with alcohol-induced psychotic disorder (diagnosis)
C2874398|Alcohol dependence with alcohol-induced persisting amnestic disorder
C2874398|Alcohol depend w alcoh-induce persisting amnestic disorder
C2874399|Alcohol dependence with alcohol-induced persisting dementia
C2874403|Alcohol dependence with other alcohol-induced disorder
C2874403|Alcohol dependence with other alcohol-induced disorders
C2874404|Alcohol dependence with unspecified alcohol-induced disorder
C0338784|alcohol dependence with episodic drinking behavior
C0338784|alcohol dependence with episodic drinking behavior (diagnosis)
C0338784|Episodic chronic alcoholism
C0338784|Episodic chronic alcoholism (disorder)
C0236656|alcohol-induced persistent dementia (diagnosis)
C0236656|alcohol-induced persistent dementia
C0236656|alcohol dependence with dementia (diagnosis)
C0236656|alcohol dependence with dementia
C0236656|Alcohol induced persisting dementia
C0236656|Alcohol persist dementia
C0236656|Dementia;alcoholic
C0236656|Alcoholic dementia NOS
C0236656|[X]Alcoholic dementia NOS
C0236656|[X]Chronic alcoholic brain syndrome
C0236656|Alcoholic dementia NOS (disorder)
C0236656|chronic organic mental disorder alcoholic brain syndrome
C0236656|Chronic alcoholic brain syndrome
C0236656|Chronic alcoholic brain syndrome (diagnosis)
C0236656|Dementia associated with alcoholism
C0236656|Alcohol-induced persisting dementia
C0236656|Alcoholic dementia
C0236656|Chronic alcoholic brain syndrome (disorder)
C0236656|Dementia associated with alcoholism (disorder)
C0236656|brain; syndrome, alcoholic (chronic)
C0236656|dementia; alcoholic
C0236656|dementia; alcohol
C0236656|alcohol; dementia
C0236656|syndrome; brain, alcoholic (chronic)
C0236656|Alcoholism associated with dementia NOS
C2874389|Alcohol dependence with withdrawal, uncomplicated
C2874389|alcohol dependence with withdrawal - uncomplicated (diagnosis)
C2874389|alcohol dependence with withdrawal - uncomplicated
C2874390|Alcohol dependence with withdrawal delirium
C2874390|alcohol dependence with withdrawal delirium (diagnosis)
C2874391|Alcohol dependence with withdrawal with perceptual disturbance
C2874391|Alcohol dependence w withdrawal with perceptual disturbance
C2874391|alcohol dependence with withdrawal with perceptual disturbance (diagnosis)
C2874395|Alcohol dependence with alcohol-induced psychotic disorder with delusions
C2874395|Alcohol depend w alcoh-induce psychotic disorder w delusions
C2874395|alcohol dependence with alcohol-induced psychotic disorder with delusions (diagnosis)
C2874396|Alcohol dependence with alcohol-induced psychotic disorder with hallucinations
C2874396|Alcohol depend w alcoh-induce psychotic disorder w hallucin
C2874396|alcohol dependence with alcohol-induced psychotic disorder with hallucinations (diagnosis)
C3509162|alcohol dependence with alcohol-induced persistng amnestic disorder
C3509162|alcohol dependence with alcohol-induced persistng amnestic disorder (diagnosis)
C3509163|alcohol dependence with alcohol-induced persistng dementia
C3509163|alcohol dependence with alcohol-induced persistng dementia (diagnosis)
C3509161|alcohol dependence with alcohol-induced disorder
C3509161|alcohol dependence with alcohol-induced disorder (diagnosis)
C2874400|Alcohol dependence with alcohol-induced anxiety disorder
C2874400|alcohol dependence with alcohol-induced anxiety disorder (diagnosis)
C2874401|Alcohol dependence with alcohol-induced sexual dysfunction
C2874401|alcohol dependence with alcohol-induced sexual dysfunction (diagnosis)
C2874402|Alcohol dependence with alcohol-induced sleep disorder
C2874402|alcohol dependence with alcohol-induced sleep disorder (diagnosis)
C2874386|Alcohol dependence with intoxication delirium
C2874386|alcohol dependence with intoxication delirium (diagnosis)
C0023896|Liver Disease, Alcoholic
C0023896|Liver Diseases, Alcoholic
C0023896|Alcoholic Liver Disease
C0023896|Alcoholic liver disease, unspecified
C0023896|LIVER DIS ALCOHOLIC
C0023896|ALCOHOLIC LIVER DIS
C0023896|alcohol induced liver disorder
C0023896|Liver Diseases, Alcoholic [Disease/Finding]
C0023896|Alcoholic Liver Diseases
C0023896|alcoholic liver disease (diagnosis)
C0023896|Alcoholic liver disease NOS
C0023896|Hepatopathy alcoholic
C0023896|ALD - Alcoholic liver disease
C0023896|disease (or disorder); liver, alcoholic
C0023896|liver; alcohol
C0023896|liver; disease, alcoholic
C0023896|alcohol; liver
C0023896|Alcoholic liver disease, NOS
C0272023|Non megaloblastic anemia due to alcoholism
C0272023|Non megaloblastic anaemia due to alcoholism
C0272023|Non megaloblastic anemia due to alcoholism (disorder)
C3839769|Alcohol dependence in childbirth (disorder)
C3839769|Alcohol dependence in childbirth
C1411379|Alcohol dependence in pregnancy (disorder)
C1411379|Alcohol dependence in pregnancy
C1411379|pregnancy; alcohol dependence
C4075901|Mild alcohol dependence (disorder)
C4075901|Mild alcohol dependence
C4075720|Severe alcohol dependence (disorder)
C4075720|Severe alcohol dependence
C4075073|Moderate alcohol dependence (disorder)
C4075073|Moderate alcohol dependence
C4076151|Thrombocytopaenia co-occurrent and due to alcoholism
C4076151|Thrombocytopenia co-occurrent and due to alcoholism
C4076151|Thrombocytopenia co-occurrent and due to alcoholism (disorder)
C0338783|Chronic alcoholism in remission
C0338783|Chronic alcoholism in remission (disorder)
C1442981|ALCOHOLIC LIVER DAMAGE
C1442981|alcoholic liver damage (diagnosis)
C1442981|Alcohol liver damage NOS
C1442981|Alcoholic liver damage unspecified (disorder)
C1442981|Alcoholic liver damage NOS (disorder)
C1442981|Alcoholic liver damage NOS
C1442981|Alcoholic liver damage unspecified
C1442981|Alcoholic liver damage, unspecified
C1442981|Alcoholic liver damage (disorder)
C1442981|damage; liver, alcoholic
C1442981|liver; damage, alcoholic
C1442981|Alcoholic liver damage, NOS
C1386568|dependence; methylated spirit
C1386568|methylated spirit; dependence
C1386585|dependence; methyl alcohol
C1386585|methyl alcohol; dependence
C1387095|poisoning; alcohol, with dependence
C1387095|alcohol; poisoning, with dependence
C1395804|drinking; excess, habit (continual)
C1395804|drinking; excessive, habit (continual)
C1395804|excess; drinking, habit (continual)
C1395804|excessive; drinking, habit (continual)
C1395805|drinking; habitual
C1395805|habitual; drinking
C0014984|ethanolism
C0392620|Alcohol poisoning
C0392620|poisoning by ethyl alcohol (diagnosis)
C0392620|poisoning by alcohol
C0392620|poisoning by alcohol (diagnosis)
C0392620|poisoning by ethyl alcohol
C0392620|Ethanol poisoning
C0392620|Ethyl alcohol poisoning
C0392620|ethylism
C0392620|poisoning; alcohol
C0392620|alcohol; poisoning
C0338787|Continuous acute alcoholic intoxication in alcoholism
C0338787|Continuous acute alcoholic intoxication in alcoholism (disorder)
C0338788|Episodic acute alcoholic intoxication in alcoholism
C0338788|Episodic acute alcoholic intoxication in alcoholism (disorder)
C0856321|Alcoholism (excluding psychosis)
C0856321|Alcoholism (excl psychosis)
C0848500|Drinks too much
C0349464|Korsakoff Syndrome
C0349464|Psychosis, Korsakoff
C0349464|Syndrome, Korsakoff
C0349464|Wernicke Korsakoff syndrome
C0349464|Korsakoff's psychosis
C0349464|Wernicke-Korsakoff syndrome
C0349464|Syndrome, Wernicke-Korsakoff
C0349464|Korsakoff's syndrome
C0349464|Wernicke Encephalopathy
C0349464|Korsakoff Psychosis
C0349464|Korsakoff Syndrome [Disease/Finding]
C0349464|Korsakoff Psychoses
C0349464|Psychoses, Korsakoff
C0349464|Syndromes, Wernicke-Korsakoff
C0349464|Wernicke-Korsakoff Syndromes
C0349464|Korsakov's psychosis
C0349464|Korsakov psychosis
C0349464|Wernicke-Korsakov syndrome (disorder)
C0349464|Wernicke-Korsakov syndrome
C0349464|Korsakov psychosis (disorder)
C0349464|Korsakoff's psychosis (diagnosis)
C0349464|ALCOHOL-INDUCED ENCEPHALOPATHY
C0349464|Korsakoff's disease
C0349464|Korsakov's syndrome
C0349464|Korsakoff's psychosis (disorder)
C0349464|Korsakov; psychosis
C0349464|Korsakov
C0349464|Korsakoffs Psychosis
C0349464|Korsakoff's psychosis, alcoholic
C0001940|Alcohol Amnestic Disorder
C0001940|Alcohol Amnestic Disorders
C0001940|Amnestic Disorder, Alcohol
C0001940|Amnestic Disorders, Alcohol
C0001940|Mental and behavioral disorders due to use of alcohol, amnesic syndrome
C0001940|Mental and behavioural disorders due to use of alcohol, amnesic syndrome
C0001940|ALCOHOL AMNESTIC DIS
C0001940|ALCOHOL IND AMNESTIC SYNDROME
C0001940|ALCOHOL IND DYSMNESIC SYNDROME
C0001940|ALCOHOL IND KORSAKOFF SYNDROME
C0001940|ALCOHOL IND PERSISTING AMNESTIC DIS
C0001940|AMNESTIC PSYCHOSIS ALCOHOL IND
C0001940|ALCOHOL IND AMNESTIC PSYCHOSIS
C0001940|ALCOHOL IND DYSMNESIC PSYCHOSIS
C0001940|alcohol-induced persisting amnestic disorder (diagnosis)
C0001940|alcohol-induced persisting amnestic disorder
C0001940|Alcohol Induced Amnestic Psychosis
C0001940|Alcohol-Induced Amnestic Psychoses
C0001940|Amnestic Psychoses, Alcohol-Induced
C0001940|Amnestic Psychosis, Alcohol Induced
C0001940|Psychoses, Alcohol-Induced Amnestic
C0001940|Psychosis, Alcohol-Induced Amnestic
C0001940|Alcohol Induced Amnestic Syndrome
C0001940|Alcohol-Induced Amnestic Syndromes
C0001940|Amnestic Syndrome, Alcohol-Induced
C0001940|Amnestic Syndromes, Alcohol-Induced
C0001940|Syndrome, Alcohol-Induced Amnestic
C0001940|Syndromes, Alcohol-Induced Amnestic
C0001940|Alcohol Amnestic Syndromes
C0001940|Amnestic Syndrome, Alcohol
C0001940|Amnestic Syndromes, Alcohol
C0001940|Syndrome, Alcohol Amnestic
C0001940|Syndromes, Alcohol Amnestic
C0001940|Alcohol Induced Dysmnesic Psychosis
C0001940|Alcohol-Induced Dysmnesic Psychoses
C0001940|Dysmnesic Psychoses, Alcohol-Induced
C0001940|Dysmnesic Psychosis, Alcohol-Induced
C0001940|Psychoses, Alcohol-Induced Dysmnesic
C0001940|Psychosis, Alcohol-Induced Dysmnesic
C0001940|Alcohol Induced Dysmnesic Syndrome
C0001940|Alcohol-Induced Dysmnesic Syndromes
C0001940|Dysmnesic Syndrome, Alcohol-Induced
C0001940|Dysmnesic Syndromes, Alcohol-Induced
C0001940|Syndrome, Alcohol-Induced Dysmnesic
C0001940|Syndromes, Alcohol-Induced Dysmnesic
C0001940|Alcohol Induced Korsakoff Syndrome
C0001940|Alcohol-Induced Korsakoff Syndromes
C0001940|Korsakoff Syndrome, Alcohol-Induced
C0001940|Korsakoff Syndromes, Alcohol-Induced
C0001940|Syndrome, Alcohol-Induced Korsakoff
C0001940|Syndromes, Alcohol-Induced Korsakoff
C0001940|Korsakoff Syndrome, Alcoholic
C0001940|Syndrome, Alcoholic Korsakoff
C0001940|Alcohol amnestic disordr
C0001940|Alcohol Amnestic Syndrome
C0001940|Alcohol-Induced Dysmnesic Syndrome
C0001940|Alcoholic Korsakoff Syndrome
C0001940|Alcohol-Induced Dysmnesic Psychosis
C0001940|Alcohol-Induced Amnestic Psychosis
C0001940|Alcohol-Induced Amnestic Syndrome
C0001940|Amnestic Psychosis, Alcohol-Induced
C0001940|Alcohol Amnestic Disorder [Disease/Finding]
C0001940|Alcohol-Induced Korsakoff Syndrome
C0001940|Korsakoffs psychosis;alcoholic
C0001940|Alcohol Induced Persisting Amnestic Disorder
C0001940|Alcoholic Korsakoff Syndromes
C0001940|Korsakoff Syndromes, Alcoholic
C0001940|Syndromes, Alcoholic Korsakoff
C0001940|Korsakoff's psychosis (alcoholic)
C0001940|[X]Korsakov's psychosis, alcohol-induced
C0001940|[X]Mental and behavioural disorders due to use of alcohol: amnesic syndrome
C0001940|[X]Mental and behavioral disorders due to use of alcohol: amnesic syndrome
C0001940|Alcohol amnestic syndrome NOS (disorder)
C0001940|[X]Mental and behavioral disorders due to use of alcohol: amnesic syndrome (disorder)
C0001940|Alcohol amnestic syndrome NOS
C0001940|Korsakoff's psychosis alcoholic
C0001940|Korsakov's psychosis, alcoholic
C0001940|Alcoholic amnestic syndrome
C0001940|Amnesic syndrome due to alcohol
C0001940|Korsakov alcoholic psychosis
C0001940|Korsakov syndrome - alcoholic
C0001940|Alcohol amnestic disorder (disorder)
C0001940|Korsakov; alcoholism
C0001940|alcohol; amnestic syndrome
C0001940|alcoholism; Korsakov
C0001940|psychosis; Korsakov, alcohol
C0001940|psychosis; alcoholic, Korsakov
C0001940|psychosis; alcoholic, polyneuritic
C0001940|amnestic; syndrome, alcohol-induced
C0001940|syndrome; amnestic, alcohol-induced
C0001940|syndrome; amnestic, alcohol
C0001940|Alcoholic Korsakoff's Psychosis
C0001940|Korsakoffs alcoholic psychosis
C0154474|Other and unspecified alcohol dependence
C0154474|Other and unspecified alcohol dependence, unspecified drinking behavior
C0154474|Alcoh dep NEC/NOS-unspec
C0154474|Other and unspecified alcohol dependence, unspecified
C0242510|Drug use
C0242510|Drug usage
C0237123|Alcohol or Other Drugs use
C0237123|Substance use
C0237123|Alcohol - drug use
