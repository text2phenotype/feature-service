C0524909|Hepatitis B, Chronic
C0744831|Chronic active hepatitis B
C0276612|Chronic active type B viral hepatitis
C0276613|Chronic persistent type B viral hepatitis
C0744833|HEPATITIS B CHRONIC PERSISTENT INFECTION
C1827079|Hepatic coma due to chronic hepatitis B
C2074982|chronic viral hepatitis delta infection with hepatitis B (diagnosis)
C2118427|acute hepatitis D infection with chronic hepatitis B
C2074977|chronic hepatitis B infection with fulminant hepatic failure
C2074978|chronic hepatitis B infection with hepatic coma
C4075603|Occult chronic type B viral hepatitis
C0375002|Chronic viral hepatitis B with hepatic coma without hepatitis delta
C0375003|Chronic viral hepatitis B with hepatic coma with hepatitis delta
C0375007|Chronic viral hepatitis B without mention of hepatic coma with hepatitis delta
C0276612|chronic active type hepatitis B virus (diagnosis)
C0276612|chronic active type hepatitis B virus
C0276612|hepatitis b virus - chronic active
C0276612|Chronic active type B viral hepatitis
C0276612|Chronic active type B viral hepatitis (disorder)
C0276613|Chronic persistent type B viral hepatitis (diagnosis)
C0276613|Chronic persistent type B viral hepatitis
C0276613|hepatitis b virus - chronic persistent
C0276613|Chronic immune tolerant hepatitis B
C0276613|Chronic persistent type B viral hepatitis (disorder)
C0276614|chronic aggressive type B viral hepatitis (diagnosis)
C0276614|chronic aggressive type B viral hepatitis
C0276614|hepatitis b virus - chronic aggressive type
C0276614|Chronic aggressive type B viral hepatitis (disorder)
C0276610|Chronic viral hepatitis B without delta-agent
C0276610|Chronic viral hepatitis B without delta-agent (disorder)
C0524909|Hepatitis B, Chronic
C0524909|chronic viral hepatitis B infection
C0524909|chronic hepatitis B infection (diagnosis)
C0524909|chronic hepatitis B infection
C0524909|chronic hepatitis, B virus
C0524909|Chronic (viral) hepatitis B
C0524909|Chronic Hepatitis B
C0524909|Hepatitis B, Chronic [Disease/Finding]
C0524909|Chronic type B viral hepatitis
C0524909|Chronic viral hepatitis B
C0524909|Chronic type B viral hepatitis (disorder)
C0524909|hepatitis; virus, chronic, type B
C0400918|Chronic viral hepatitis B with delta-agent
C0400918|chronic viral hepatitis B infection with hepatitis delta
C0400918|chronic hepatitis B infection with hepatitis delta
C0400918|chronic hepatitis, B virus with hepatitis delta
C0400918|chronic hepatitis B infection with hepatitis delta (diagnosis)
C0400918|Chronic viral hepatitis B with hepatitis D
C0400918|Chronic viral hepatitis B with hepatitis D (disorder)
C0400918|hepatitis; virus, chronic, type B, with delta-agent
C2074978|chronic hepatitis, B virus with hepatic coma
C2074978|chronic viral hepatitis B infection with hepatic coma
C2074978|chronic hepatitis B infection with hepatic coma
C2074978|chronic hepatitis B infection with hepatic coma (diagnosis)
C2074976|chronic hepatitis B infection with coma with hepatitis delta (diagnosis)
C2074976|chronic hepatitis B infection with coma with hepatitis delta
C2074976|chronic hepatitis, B virus coma with hepatitis delta
C2074976|chronic viral hepatitis B infection with coma with hepatitis delta
C2074977|chronic viral hepatitis B infection with fulminant hepatic failure
C2074977|chronic hepatitis B infection with fulminant hepatic failure (diagnosis)
C2074977|chronic hepatitis B infection with fulminant hepatic failure
C2074977|chronic hepatitis, B virus with fulminant hepatic failure
C3838179|hepatitis, b virus - chronic without hepatitis delta
C3838179|chronic hepatitis, B virus without hepatitis delta (diagnosis)
C3838179|chronic hepatitis, B virus without hepatitis delta
C4075603|Occult chronic type B viral hepatitis (disorder)
C4075603|Occult chronic type B viral hepatitis
C4075603|Occult hepatitis B infection
C1827079|Chronic viral hepatitis B with hepatic coma
C1827079|Hepatic coma due to chronic hepatitis B (disorder)
C1827079|Chronic hepatitis B with hepatic coma
C1827079|Hepatic coma due to chronic hepatitis B
C1827079|Chronic hepatitis B with hepatic coma (disorder)
C0494789|Chronic active hepatitis, not elsewhere classified
C0494787|Chronic persistent hepatitis, not elsewhere classified
C4041189|Hepatic coma due to chronic hepatitis B with delta agent (disorder)
C4041189|Hepatic coma due to chronic hepatitis B with delta agent
C2074981|chronic hepatitis D infection with chronic hepatitis B (diagnosis)
C2074981|chronic hepatitis, delta virus with chronic Hepatitis B
C2074981|chronic hepatitis D infection with chronic hepatitis B
C2074983|chronic hepatitis D infection with hepatitis B carrier state (diagnosis)
C2074983|chronic hepatitis, delta virus with carrier state Hepatitis B
C2074983|chronic hepatitis D infection with hepatitis B carrier state
C0375002|Hpt B chrn coma wo dlta
C0375002|Chronic viral hepatitis B with hepatic coma without hepatitis delta
C0375002|Viral hepatitis B with hepatic coma, chronic, without mention of hepatitis delta
C0375003|Hpt B chrn coma w dlta
C0375003|Chronic viral hepatitis B with hepatic coma with hepatitis delta
C0375007|Hpt B chrn wo cm w dlta
C0375007|Chronic viral hepatitis B without mention of hepatic coma with hepatitis delta
