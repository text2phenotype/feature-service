General|attraction||phil||attraction
General|attraction||philia||attraction
General|auto|auto|||
General|base|bas||basolateral|base
General|base|basi||basicranial|base
General|base|basio||basioccipital|base
General|base|baso||basophil|base
General|bio|bio||biology|life
General|break||clast||to break
General|chem|chem||chemistry|chemistry, drug
General|chem|pharma||pharmacology|
General|de|de|||dephosphated (noise?)
General|enzyme||ase||enzyme
General|fake|pseud/o||pseudoephedrine|denotes something false or fake
General|flow||flux|reflux|to flow, flow, flowing
General|flow||rrhea|diarrhea|discharge, flow
General|genetics|hered|||inheritance
General|healthy|eu||euthymia|healthy, normal
General|healthy|bene||beneficial|good
General|water|hydr/o||hydrocele|hydrogen, water
General|study||logy|biology|study of
General|study||gnosis|diagnosis|knowledge
General|meta|meta||metastasis|beyond
General|new|neo|||new
General|post|post||postmastectomy|after, behind
General|pro|pro|||
General|production||plasia|dysplasia|formation, development
General|production||trophy|hypertrophy|development, process of nourishment
General|production||poiesis|Thrombopoiesis|formation, production
General|production||genesis|spermatogenesis|production, origin
General|production||gen||producing, produced by
General|protection||phylaxis|prophylaxis|protection
General |protein|albumin||albuminuria|protein
General|re|re|||regurgitation (noise?)
General|specialist||ician|physician|specialist
General|specialist||logist|oncologist|
General|specialist||ist|radiologist|specialist
General|split||fida||to split, splitting
General|stasis||stasis|hemostasis|stopping, controlling
General|syn|syn|||
General|anti|contra||contralateral|opposite, against
General|anti|anti||antibacterial|against
General|different|allo|||other, different
General|different|hetero||heterozygous|other, different
General|same|homo||homogenous|same
General|same|homeo||homeostasis|
General|non|non||nonbacterial|not
General|non|non-||non-hodgkin's|not
