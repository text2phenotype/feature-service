Condition|abnormal|dys||dysplastic|abnormal, bad, painful, difficult
Condition|abnormal|mal||malnutrition|poor, bad
Condition|abnormal|para||parakeratosis|abnormal, near, beside
Condition|abnormal||osis|keratosis|abnormal condition
Condition|abnormal||pathy|nephrapathy|disease process
Condition|abnormal||plakia|leukoplakia|condition of patches
Condition|bone||malacia|osteomalacia|condition of softening
Condition|cancer|carcin||carcinogen|cancer
Condition|cancer||sarcoma|osteosarcoma|connective tissue cancer
Condition|cancer||carcinoma|choriocarcinoma|cancer of epithelial origin
Condition|cancer||oma||tumor, mass
Condition|cancer||plasm|neoplasm|condition of formation
Condition|cancer||cytoma|astrocytoma|cell tumor
Condition|cells||cytosis|lymphocytosis|abnormal increase of cells
Condition|cells||emia|anemia|blood condition
Condition|colorectal||chezia|hematochezia|condition of stools
Condition|death|necr||necrosis|death (especially tissue)
Condition|digestive||dipsia|polydipsia|diet, condition of thirst
Condition|digestive||orexia|anorexia|diet, appetite condition
Condition|digestive||pepsia|dyspepsia|digestion condition
Condition|digestive||phagia|dysphagia|condition of swallowing, eating
Condition|digestive||chalasia|achalasia|condition of relaxation (throat/digestive)
Condition|displacement||ptosis|blepharoptosis|drooping, prolapse, falling
Condition|displacement||lapse|prolapse|to fall, to slide, to sag
Condition|displacement||listhesis|spondylolisthesis|slippage
Condition|drome||drome||to run, running
Condition|enlargement||megaly|cardiomegaly|enlargement
Condition|enlargement||ectasis|bronchiectasis|dilation
Condition|eye||opia|hyperopia|vision condition
Condition|eye||opsia|bradyopsia|vision condition
Condition|fast|tachy||tachypnea|rapid, fast
Condition|fast|oxy|||rapid
Condition|hardening|isch||ischemia|restriction, constricted (blood)
Condition|hardening|scler/o||sclerosis|hard; hardened; hardening
Condition|hardening||sclerosis|atherosclerosis|abnormal hardening of tissue
Condition|hardening||stenosis|arteriostenosis|abnormal condition of narrowing
Condition|heart||cardia|tachycardia|condition of the heart
Condition|heart||cardial|myocardial|condition of the heart
Condition|hyper|hyper||hyperextension|excessive, above
Condition|hypo|hypo||hypodermic|deficient, below, under, decreased
Condition|hypo||penia|thrombocytopenia|deficiency
Condition|infection||virus|parvovirus|pertaining to virus
Condition|infection|bacteri||bacterial|pertaining to bacteria
Condition|inflammation||itis|tracheobronchitis|infammation
Condition|itch|psor||psoriasis|
Condition|lung||pnea|apnea|breathing
Condition|psych||phrenia|schizophrenia|denoting something "split" or "double-sided"
Condition|psych||phobia|acrophobia|condition of fear, extreme sensitivity
Condition|psych||mania|trichotillomania|condition of madness
Condition|psych||thymia|dysthymia|condition, state of mind
Condition|movement||paresis|hemiparesis|slight paralysis
Condition|movement||plegia|paraplegia|paralysis
Condition|movement|scoli/o||scoliosis|curved, bent
Condition|movement||sthenia|myasthenia|condition of strength
Condition|pain||algia|cephalalgia|pain
Condition|pain||dynia|pharyngodynia|pain
Condition|PertainingTo||ism|hypersplenism|condition, state of
Condition|PertainingTo||ia|dysphoria|condition
Condition|PertainingTo||iasis|cholelithiasis|condition, process of
Condition|PertainingTo||lysis|onycholysis|loosening, breaking down, freeing from adhesions, separation
Condition|rupture||rrhage|hemorrhage|bursting forth, rupture
Condition|rupture||rrhexis|angiorrhexis|rupture
Condition|rupture||spadias|hypospadias|tear
Condition|rupture|herni||hernia|protrusion, rupture
Condition|seizure||lepsy||seizure
Condition|skin|ichthy/o|||skin condition
Condition|slow|brady||bradycardia|slow
Condition|spasm||ismus||spasm, contraction
Condition|spasm||spasm||sudden, involuntary contraction
Condition|spine|spondyl/o||spondylolisthesis|change in vertebrae
Condition|swelling||edema|lymphedema|swelling
Condition|swelling||cele|hydrocele|herniation, protrusion
Condition|tension||tension||pressure, process of stretching
Condition|thromb|thromb||thrombosis|blood clot; coagulation; thrombin
Condition|toxin|tox||toxoplasmosis|toxin, poison
Condition|urinary||uria|hematuria|urinary condition
Condition|vomit||emesis|hematemesis|vomiting
Condition|vomit||ptysis|hemoptysis|spitting
