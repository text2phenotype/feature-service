C0007634|T025|cells|
C0005767|T024|blood|
C3668946|T033|activity|
C0007634|T025|cell|
C0087111|T061|treatment|
C0449201|T029|per|
C0012634|T047|disease|
C0392148|T061|presence|
C0086045|T041|concentration|
C0040300|T024|tissue|
C0440102|T130|various|
C0033684|T123|protein|
C0033684|T116|protein|
C3714514|T046|infection|
C0086045|T041|concentrations|
C1272883|T122|injection|
C1533685|T061|injection|
C0445223|T033|related|
C0023884|T023|liver|
C0002778|T059|analysis|
C0456984|T033|test|
C0221198|T033|lesions|
C0001554|T057|administration|
C1533734|T061|administration|
C0014442|T109|enzyme|
C0014442|T126|enzyme|
C0011900|T033|diagnosis|
C0040300|T024|tissues|
C0456984|T033|Tests|
C0043047|T197|water|
C0043047|T121|water|
C0460139|T033|pressure|
C1764827|T123|isolated|
C0439631|T061|primary|
C0087111|T061|therapy|
C1444656|T033|indicated|
C1304686|T034|pH|lab,
C0456984|T033|tested|
C0080194|T037|strain|
C0080194|T037|strains|
C0225810|T029|basis|
C0003241|T129|antibody|
C0003241|T116|antibody|
C0021469|T044|inhibition|
C0441610|T061|reduction|
C2242979|T059|culture|
C2242979|T059|cultures|
C1123023|T022|skin|
C1689985|T190|absence|
C1292856|T061|stimulation|
C0026845|T024|muscle|
C0037473|T123|Sodium|
C0037473|T196|Sodium|
C0018787|T023|heart|
C0013227|T121|drug|
C0003320|T129|antigen|
C0225810|T029|based|
C0006104|T023|brain|
C0442726|T033|detected|
C0033684|T123|proteins|
C0033684|T116|proteins|
C0184661|T061|procedure|
C0001721|T041|affected|
C0003241|T129|antibodies|
C0003241|T116|antibodies|
C0027651|T191|tumor|
C0332575|T033|red|
C0022646|T023|renal|
C4082130|T033|prepared|
C0274281|T037|exposure|
C0332293|T061|treated with|
C0043227|T057|work|
C1306577|T033|Death|
C0022646|T023|Kidney|
C0018563|T023|hand|
C0025344|T040|periods|
C0027740|T024|nerve|
C0262950|T023|bone|
C0025519|T040|metabolism|
C0017725|T123|glucose|lab,
C0017725|T109|glucose|lab,
C0017725|T121|glucose|lab,
C0557351|T033|employed|social,
C0013227|T121|drugs|
C0024109|T023|lung|
C0030054|T196|Oxygen|treatment,
C0030054|T121|Oxygen|treatment,
C1272883|T122|injections|
C1533685|T061|injections|
C0042196|T061|inoculation|
C0012854|T123|DNA|
C0012854|T114|DNA|
C0233324|T040|term|
C3714514|T046|infections|
C0427965|T033|sensitivity|
C0221198|T033|lesion|
C3668946|T033|activities|
C0015252|T061|removal|
C0027651|T191|tumors|
C0012634|T047|diseases|
C1963578|T061|release|
C1299583|T033|independent|
C0184661|T061|procedures|
C0039082|T047|syndrome|
C0033213|T033|problems|
C0033213|T033|problem|
C0087111|T061|therapeutic|
C0014442|T109|enzymes|
C0014442|T126|enzymes|
C3263723|T037|injury|
C0037993|T023|spleen|
C0019932|T125|hormone|
C0003320|T129|antigens|
C0006675|T123|calcium|lab,
C0006675|T123|calcium|lab,medication,
C0006675|T196|calcium|lab,
C0006675|T196|calcium|lab,medication,
C0006675|T121|calcium|lab,
C0006675|T121|calcium|lab,medication,
C0226896|T030|oral|
C0344211|T061|support|
C0005847|T023|vascular|
C0577559|T033|mass|
# C0006826|T191|cancer| JIRA/SANDS-173
C0311392|T033|signs|
C0007097|T191|carcinoma|
C0004083|T041|association|
# C0028158|T196|nitrogen| JIRA/BIOMED-375
C0026018|T059|microscopy|lab,
C0027769|T184|nervous|
C0233324|T040|terms|
C0022023|T196|ion|
C0009498|T116|complement|
C0009498|T129|complement|
C0031603|T121|phosphate|lab,
C0031603|T197|phosphate|lab,
C0024264|T025|lymphocytes|lab,
C2752151|T122|extracts|
C0162867|T024|media|
C0596019|T196|chloride|lab,
C0009566|T046|complications|
C0010957|T037|damage|
C0001924|T123|albumin|lab,
C0001924|T116|albumin|lab,
C0086972|T033|separated|
C0032961|T040|pregnancy|diagnosis,
C0032961|T040|pregnancy|diagnosis,problem,
C0449416|T033|source|
C1510438|T059|assay|
C0005847|T023|vessels|
# C0032821|T196|potassium|lab,
# C0032821|T196|potassium|lab,medication, JIRA/BIOMED-376
C0017243|T122|gel|
C0003842|T023|artery|
C0262926|T033|history|
C1299581|T033|able|
C0015967|T033|fever|
C0449381|T033|parameters|
C0021853|T023|intestinal|
C0085639|T033|fall|
C3536832|T121|air|
C3536832|T197|air|
C1546956|T033|died|
C0022023|T196|ions|
C0010834|T026|cytoplasm|
C0597357|T192|receptor|
C0597357|T116|receptor|
C0023175|T196|leads|
C0023175|T131|leads|
C0013842|T059|electron microscopy|lab,
C0014609|T024|epithelium|
C1261381|T061|destruction|
C2752151|T122|extract|
C0007610|T026|nuclei|
C0004268|T041|attention|
C0023175|T196|led|
C0023175|T131|led|
C0185023|T061|fixation|
C0024109|T023|lungs|
C1314687|T033|sex|
C0007009|T196|carbon|
C0228174|T023|cerebral|
C0005823|T040|blood pressure|lab,
C0014792|T025|erythrocytes|
C0013879|T196|elements|
C0007610|T026|nucleus|
C0225810|T029|base|
C0597357|T192|receptors|
C0597357|T116|receptors|
C0014653|T040|equilibrium|
C0030193|T184|pain|problem,
C0029974|T025|egg|
C0019046|T123|hemoglobin|lab,
C0019046|T116|hemoglobin|lab,
C0518015|T059|hemoglobin|lab,
C0027763|T022|nervous system|
C0021400|T047|influenza|immunization,
C0021400|T047|influenza|immunization,lab,
C0021400|T047|influenza|immunization,lab,diagnosis,
C0021400|T047|influenza|immunization,lab,diagnosis,problem,
C0205054|T029|hepatic|
C0026237|T026|mitochondria|
C0038720|T197|sulfate|
C1522449|T061|radiation|
C0005528|T043|transport|
C0038960|T122|suspensions|
C0225326|T121|fibers|
C0005615|T040|birth|
C0020275|T196|hydrogen|
C0013855|T059|electrophoresis|
C0574032|T061|infusion|
C0011570|T048|depression|diagnosis,
C0011570|T048|depression|diagnosis,problem,
C0600688|T037|Toxicity|
C0012634|T047|disorders|
C0035668|T114|RNA|
C0015677|T109|fat|
C0015677|T121|fat|
C0023779|T109|lipid|
C0334094|T046|proliferation|
C0026845|T024|Muscles|
C0030011|T044|oxidation|
C1306645|T060|x-ray|lab,
C0442739|T033|unchanged|
C0001975|T121|alcohol|social,
C0001975|T109|alcohol|social,
C0027540|T042|necrosis|
C0038960|T122|suspension|
C0015392|T023|eye|
C0008377|T123|cholesterol|lab,
C0008377|T109|cholesterol|lab,
C0020538|T047|hypertension|diagnosis,
C0020538|T047|hypertension|diagnosis,problem,
C0079240|T059|dilution|
C0005953|T024|bone marrow|
C0032285|T047|pneumonia|diagnosis,
C0032285|T047|pneumonia|diagnosis,problem,
C3853573|T122|granules|
C0017649|T123|globulin|lab,
C0017649|T116|globulin|lab,
C0028778|T046|obstruction|
C0042210|T121|vaccine|
C0042210|T129|vaccine|
C0449416|T033|sources|
C0022646|T023|kidneys|
C0021641|T121|insulin|medication,
C0021641|T116|insulin|medication,
C0021641|T125|insulin|medication,
C0007004|T109|carbohydrate|
C0002520|T116|amino acids|
C0002520|T123|amino acids|
C0002520|T121|amino acids|
C0040132|T023|thyroid|
C2752151|T122|extracted|
C0011164|T046|degeneration|
C1697794|T122|liquid|
C0000726|T029|abdominal|
C0032005|T023|pituitary|
C0042890|T127|Vitamin|
C0042890|T109|Vitamin|
C0042890|T121|Vitamin|
C0233494|T048|tension|
C0020971|T061|immunization|
C0002520|T116|amino acid|
C0002520|T123|amino acid|
C0002520|T121|amino acid|
C0021853|T023|intestine|
C0020960|T121|antiserum|
C0020960|T129|antiserum|
C0020960|T116|antiserum|
C0002871|T047|anemia|diagnosis,
C0002871|T047|anemia|diagnosis,problem,
C0185115|T061|Extraction|
C0032932|T044|precipitation|
C0041236|T116|trypsin|lab,
C0041236|T126|trypsin|lab,
C0041236|T121|trypsin|lab,
C0026649|T040|movement|
C0302583|T123|iron|lab,
C0302583|T123|iron|lab,medication,
C0302583|T196|iron|lab,
C0302583|T196|iron|lab,medication,
C0302583|T121|iron|lab,
C0302583|T121|iron|lab,medication,
C0699748|T046|pathogenesis|
C0038435|T033|stress|problem,
C0344315|T033|depressed|
C0029974|T025|eggs|
C0221423|T184|illness|
C0001801|T044|agglutination|
C0027740|T024|nerves|
C0005558|T060|biopsy|lab,
C0005558|T060|biopsy|lab,procedure,
C0023175|T196|Lead|lab,
C0023175|T196|Lead|lab,social,
C0023175|T131|Lead|lab,
C0023175|T131|Lead|lab,social,
C0018670|T029|head|
C0549206|T033|pregnant|
C0030016|T116|dehydrogenase|
C0030016|T126|dehydrogenase|
C2242979|T059|cultured|
C1510420|T190|cavity|
C0683278|T048|suffering|
C0589120|T033|follow-up|
C0024264|T025|lymphocyte|lab,
C0041296|T047|tuberculosis|diagnosis,
C0041296|T047|tuberculosis|diagnosis,problem,
C0037494|T121|NaCl|medication,
C0037494|T123|NaCl|medication,
C0037494|T197|NaCl|medication,
C1510411|T046|transformation|
C0003842|T023|arteries|
C0035295|T023|reticulum|
C0521119|T026|extracellular|
C0000975|T109|acetate|
C0000975|T121|acetate|
C0023516|T025|leucocytes|lab,
C0002778|T059|analyses|
C0038351|T023|stomach|
C0035253|T056|resting|
C0027651|T191|tumour|
C3714787|T022|central nervous system|
C1140999|T046|contraction|
C0036974|T046|shock|diagnosis,
C0036974|T046|shock|diagnosis,problem,
C1963578|T061|released|
C0021368|T046|inflammation|
C0020960|T121|antisera|
C0020960|T129|antisera|
C0020960|T116|antisera|
C0030274|T023|pancreatic|
C0038128|T130|stained|
C0199176|T061|prevention|
C0152060|T061|division|
C0001771|T121|agar|
C0001771|T130|agar|
C0001771|T109|agar|
C0036679|T046|separation|
C0019932|T125|hormones|
C0442034|T029|peritoneal|
C0035253|T056|rest|
C1306577|T033|deaths|
C0031678|T116|phosphatase|
C0031678|T126|phosphatase|
C0042449|T023|vein|
C0027882|T025|neurons|
C0009780|T024|connective tissue|
C0013604|T033|edema|problem,
C0005773|T025|blood cells|
C0019080|T046|bleeding|
C0038636|T123|sucrose|medication,
C0038636|T121|sucrose|medication,
C0038636|T109|sucrose|medication,
C0439775|T061|elevation|
C0023175|T196|leading|
C0023175|T131|leading|
C0028778|T046|block|
C0008633|T026|chromosome|
C0006901|T023|capillary|
C3714660|T037|trauma|problem,
C0185117|T061|expression|
C0006901|T023|capillaries|
C0003232|T195|antibiotic|
C0006141|T023|breast|
C0038999|T033|swelling|
C0016030|T025|fibroblasts|
C0439857|T048|dependence|
C2239178|T033|newborn|
C0232338|T040|blood flow|
C0024432|T025|macrophages|
C0024204|T023|lymph nodes|
C0020852|T116|IgG|lab,
C0020852|T129|IgG|lab,
C0020852|T121|IgG|lab,
C0442811|T033|very low|
C0728940|T061|resection|
C0030274|T023|pancreas|
C0022417|T030|joint|
C0040549|T123|toxin|
C0040549|T131|toxin|
C0032594|T121|polysaccharide|
C0032594|T109|polysaccharide|
C0013343|T130|dye|
C0035139|T061|replacement|
C0041942|T121|urea|lab,
C0041942|T123|urea|lab,
C0041942|T109|urea|lab,
C0019080|T046|hemorrhage|
C1299586|T033|difficulties|
C0222045|T023|scale|
C0014792|T025|erythrocyte|lab,
C1378566|T122|solid|
C0007703|T059|centrifugation|
C0233660|T048|blocking|
C0524637|T041|recognition|
C0023418|T191|leukemia|diagnosis,
C0023418|T191|leukemia|diagnosis,problem,
C0014653|T040|balance|
C0003232|T195|antibiotics|
C0001721|T041|affecting|
C0031001|T061|perfusion|
C0242209|T109|sugar|
C0242209|T121|sugar|
C0699900|T040|degradation|
C0009443|T047|cold|
C0037925|T023|spinal cord|
C0344211|T061|supported|
C0031308|T043|phagocytosis|
C1184740|T023|tubercle|
C0301625|T040|suppression|
C0557061|T061|DISCUSSION|
C3665472|T061|chemotherapy|procedure,
C0456909|T033|blind|
C0817096|T029|chest|
C0332293|T061|treated by|
C0040113|T023|thymus|
C0684321|T041|regression|
C0019588|T109|histamine|lab,
C0019588|T123|histamine|lab,
C0162340|T041|understanding|
C0004398|T060|autopsy|procedure,
C0003483|T023|aortic|
C0034929|T042|reflex|
C0005682|T023|bladder|
C0024348|T046|lysis|
C0028778|T046|occlusion|
C0026649|T040|movements|
C0014597|T025|epithelial cells|
C0687028|T023|duct|
C0012634|T047|disorder|
C0007332|T116|casein|
C0007332|T121|casein|
C1299582|T033|unable|
C0424927|T033|education|
C0002903|T061|anesthesia|procedure,
C0017237|T121|gelatin|
C0017237|T116|gelatin|
C0017237|T122|gelatin|
C0374711|T061|repair|
C1947940|T122|oil|
C0038317|T109|steroid|medication,
C1444775|T033|sharp|
C0460139|T033|pressures|
C0071499|T122|polyacrylamide|
C0071499|T109|polyacrylamide|
C0034963|T042|regeneration|
C0560175|T033|carrier|
C0042196|T061|vaccination|
C0030956|T116|peptide|
C0442739|T033|no change|
C1627358|T061|enhancement|
C0014239|T026|endoplasmic reticulum|
C1304680|T033|attack|
C0600138|T033|plays|
C1510438|T059|assays|
C0000925|T037|cut|
C1261473|T191|sarcoma|diagnosis,
C1261473|T191|sarcoma|diagnosis,problem,
C0220892|T195|penicillin|allergy,
C0220892|T195|penicillin|allergy,medication,
C0220892|T109|penicillin|allergy,
C0220892|T109|penicillin|allergy,medication,
C0684336|T046|impairment|
C0015259|T056|exercise|social,
C0032961|T040|gestation|
C0085639|T033|fell|
C0009566|T046|complication|
C0085672|T059|micro|
C0425245|T033|mobility|
C0017547|T047|giant|
C0009325|T116|collagen|
C0031705|T196|phosphorus|lab,
C0242417|T116|oxidase|
C0242417|T126|oxidase|
C0225326|T121|fibres|
C0014994|T121|ether|medication,
C0014994|T109|ether|medication,
C0027651|T191|TUMOURS|
C0596012|T033|reaches|
C0028429|T023|nasal|
C0013227|T121|medicine|
C0033308|T121|progesterone|lab,
C0033308|T121|progesterone|lab,medication,
C0033308|T125|progesterone|lab,
C0033308|T125|progesterone|lab,medication,
C0033308|T109|progesterone|lab,
C0033308|T109|progesterone|lab,medication,
C0332448|T046|infiltration|
C0702249|T061|infiltration|
C0015684|T109|fatty acids|
C0002611|T197|ammonium|
C0020507|T046|hyperplasia|
C1299586|T033|difficulty|
C0011209|T061|delivery|
C0311392|T033|sign|
C0033727|T196|hydrogen ion|
C1283786|T023|blood vessels|
C0034580|T059|radioimmunoassay|lab,
C0001443|T123|adenosine|medication,
C0001443|T114|adenosine|medication,
C0001443|T121|adenosine|medication,
C0015392|T023|eyes|
C0008633|T026|chromosomes|
C0005821|T025|platelet|lab,
C0005821|T025|platelet|lab,treatment,
C0003864|T047|arthritis|diagnosis,
C0003864|T047|arthritis|diagnosis,problem,
C0014792|T025|red blood cells|lab,
C1277078|T121|red blood cells|lab,
C0557854|T057|service|
C0021308|T046|infarction|
C0445356|T033|unrelated|
C0040077|T123|thymidine|lab,
C0040077|T114|thymidine|lab,
C0020564|T046|hypertrophy|
C0181074|T122|graft|
C0001041|T121|acetylcholine|medication,
C0001041|T109|acetylcholine|medication,
C0001041|T123|acetylcholine|medication,
C0043227|T057|working|
C0522224|T033|paralysis|diagnosis,
C0522224|T033|paralysis|diagnosis,problem,
C0232217|T042|conduction|
C0230445|T029|calf|
C0523465|T059|serum albumin|lab,
C0564405|T033|relief|
C0376261|T109|lactate|lab,
C0376261|T121|lactate|lab,
C1295697|T034|axis|
C0004457|T023|axis|
C0333641|T046|atrophy|
C0817096|T029|thoracic|
C0039601|T121|testosterone|lab,
C0039601|T121|testosterone|lab,medication,
C0039601|T125|testosterone|lab,
C0039601|T125|testosterone|lab,medication,
C0039601|T109|testosterone|lab,
C0039601|T109|testosterone|lab,medication,
C1325847|T040|sensitization|
C0027530|T029|neck|
C0040732|T061|transplantation|
C0022663|T023|glomerular|
C1444648|T033|offered|
C0024467|T196|magnesium|lab,
C0024467|T196|magnesium|lab,medication,
C0043240|T040|healing|
C0557854|T057|services|
C0226896|T030|mouth|
C0017911|T123|glycogen|
C0017911|T109|glycogen|
C0225326|T121|fiber|
C0003483|T023|aorta|
C0035298|T023|retinal|
C0035331|T121|retinal|
C0035331|T127|retinal|
C0035331|T109|retinal|
C0442737|T033|not found|
C0009368|T023|colon|
C0007012|T123|carbon dioxide|lab,
C0007012|T197|carbon dioxide|lab,
C0011946|T061|dialysis|procedure,
C0021027|T121|immunoglobulin|
C0021027|T116|immunoglobulin|
C0021027|T129|immunoglobulin|
C0728940|T061|excision|
C0001465|T121|AMP|
C0001465|T123|AMP|
C0001465|T114|AMP|
C0023607|T125|LH|lab,
C0023607|T116|LH|lab,
C0023607|T121|LH|lab,
C3263723|T037|Injuries|
C0018827|T023|ventricle|
C0589507|T041|initiation|
C0020517|T046|hypersensitivity|
C0085639|T033|falls|
C0020564|T046|enlargement|
C1293134|T061|enlargement|
C2711450|T190|enlargement|
C0013030|T121|dopamine|medication,
C0013030|T109|dopamine|medication,
C0013030|T123|dopamine|medication,
C0001804|T129|agglutinins|
C0087111|T061|treatments|
C0303920|T130|fluorescent|
C0303920|T109|fluorescent|
C0042149|T023|uterus|
C0023516|T025|leukocytes|lab,
C2937287|T043|hemolysis|diagnosis,
C2937287|T043|hemolysis|diagnosis,problem,
C1720436|T033|anesthetized|
C1546956|T033|dead|
C0442804|T033|very high|
C2939419|T191|metastases|diagnosis,
C2939419|T191|metastases|diagnosis,problem,
C0004461|T026|axons|
C1510438|T059|assayed|
C0002055|T197|alkali|
C1261287|T046|stenosis|
C0043250|T037|wound|
C0023884|T023|livers|
C0560175|T033|carriers|
C0041485|T123|tyrosine|lab,
C0041485|T123|tyrosine|lab,medication,
C0041485|T116|tyrosine|lab,
C0041485|T116|tyrosine|lab,medication,
C0041485|T121|tyrosine|lab,
C0041485|T121|tyrosine|lab,medication,
C0020861|T116|IgM|lab,
C0020861|T129|IgM|lab,
C0013443|T023|ear|
C0205039|T023|bronchial|
C0728899|T033|intoxication|
C0029266|T041|orientation|
C0025552|T197|metal|
C0229889|T023|lymphatic|
C0010454|T130|culture medium|
C0004259|T121|atropine|medication,
C0004259|T109|atropine|medication,
C0014912|T121|estradiol|lab,
C0014912|T121|estradiol|lab,medication,
C0014912|T125|estradiol|lab,
C0014912|T125|estradiol|lab,medication,
C0014912|T109|estradiol|lab,
C0014912|T109|estradiol|lab,medication,
C0013832|T197|electrolytes|
C0013832|T121|electrolytes|
C0041466|T047|typhoid|diagnosis,
C0041466|T047|typhoid|diagnosis,problem,
C0041296|T047|tuberculous|diagnosis,
C0041296|T047|tuberculous|diagnosis,problem,
C0023779|T109|lipids|
C0019158|T047|hepatitis|diagnosis,
C0019158|T047|hepatitis|diagnosis,problem,
C0016006|T121|fibrinogen|lab,
C0016006|T123|fibrinogen|lab,
C0016006|T116|fibrinogen|lab,
C0431085|T025|tumor cells|
C0028630|T114|nucleotide|
C0013832|T197|electrolyte|
C0013832|T121|electrolyte|
C0005847|T023|vessel|
C0030471|T030|sinus|
C0014939|T121|estrogen|lab,
C0014939|T121|estrogen|lab,medication,
C0014939|T125|estrogen|lab,
C0014939|T125|estrogen|lab,medication,
C0014939|T109|estrogen|lab,
C0014939|T109|estrogen|lab,medication,
C0011906|T060|differential diagnosis|
C0007301|T024|cartilage|
C0040284|T059|tissue culture|
C0015982|T121|fibrin|
C0015982|T123|fibrin|
C0015982|T116|fibrin|
C0015663|T033|fasting|
C0013303|T023|duodenal|
C0007603|T026|cell membrane|
C0042449|T023|veins|
C0005821|T025|platelets|lab,
C0577559|T033|masses|
C0038317|T109|steroids|
C0544452|T033|remission|
C1282864|T030|lumen|
C0079603|T059|immunofluorescence|
C0017861|T121|glycerol|
C0017861|T123|glycerol|
C0017861|T109|glycerol|
C0013103|T061|drainage|
C0016059|T046|fibrosis|
C0014038|T047|encephalitis|diagnosis,
C0014038|T047|encephalitis|diagnosis,problem,
C0007097|T191|carcinomas|
C0005558|T060|biopsies|procedure,
C0003765|T123|arginine|medication,
C0003765|T116|arginine|medication,
C0003765|T121|arginine|medication,
C0032961|T040|pregnancies|
C0007603|T026|plasma membrane|
C0008238|T131|chloroform|medication,
C0008238|T130|chloroform|medication,
C0008238|T109|chloroform|medication,
C1267092|T024|smooth muscle|
C0151526|T033|premature|
C0205054|T029|portal|
C1305923|T116|polypeptide|
C0181074|T122|grafts|
C1258666|T047|ganglia|
C0079240|T059|dilutions|
C0024337|T121|lysine|medication,
C0024337|T123|lysine|medication,
C0024337|T116|lysine|medication,
C0002978|T060|angiography|procedure,
C0040053|T046|thrombosis|
C0033371|T125|prolactin|lab,
C0033371|T116|prolactin|lab,
C0033371|T121|prolactin|lab,
C0008546|T116|chromatin|
C0041582|T047|ulcer|problem,
C0042232|T023|vaginal|
C0027051|T047|myocardial infarction|diagnosis,
C0027051|T047|myocardial infarction|diagnosis,problem,
C0020663|T023|hypothalamus|
C0018799|T047|heart disease|problem,
C0009968|T123|copper|lab,
C0009968|T196|copper|lab,
C0009968|T121|copper|lab,
C0344211|T061|supports|
C0037868|T025|Sperm|
C1964256|T060|illumination|
C0332835|T024|transplanted|
C0040732|T061|transplanted|
C0030909|T121|pepsin|medication,
C0030909|T116|pepsin|medication,
C0014257|T024|endothelium|
C0009356|T121|collodion|medication,
C0009356|T109|collodion|medication,
C0021852|T023|small intestine|
C0332837|T037|implanted|
C1704229|T122|implanted|
C0021107|T061|implantation|
C1704608|T122|films|
C0028778|T046|blocked|
C1304680|T033|attacks|
C0041289|T116|tuberculin|medication,
C0041289|T130|tuberculin|medication,
C0041289|T129|tuberculin|medication,
C0039128|T047|syphilis|diagnosis,
C0039128|T047|syphilis|diagnosis,problem,
C0025646|T121|methionine|medication,
C0025646|T123|methionine|medication,
C0025646|T116|methionine|medication,
C0021968|T121|iodine|medication,
C0021968|T196|iodine|medication,
C0019134|T109|heparin|medication,
C0019134|T121|heparin|medication,
C0019134|T123|heparin|medication,
C0001962|T121|ethanol|lab,
C0001962|T121|ethanol|lab,social,
C0001962|T109|ethanol|lab,
C0001962|T109|ethanol|lab,social,
C0028778|T046|blocking|
C3203359|T037|rupture|
C0035298|T023|retina|
C0202165|T059|hydrogen ion concentration|
C0012359|T046|dilatation|
C0037494|T121|sodium chloride|medication,
C0037494|T123|sodium chloride|medication,
C0037494|T197|sodium chloride|medication,
C0849912|T033|emotional|
C1140999|T046|contractions|
C0007648|T123|cellulose|
C0007648|T109|cellulose|
C0001916|T019|albino|
C0001721|T041|affects|
C0023401|T123|leucine|medication,
C0023401|T116|leucine|medication,
C0023401|T121|leucine|medication,
C1704608|T122|film|
C0332128|T033|examined for|
C0001655|T125|ACTH|lab,
C0001655|T116|ACTH|lab,
C0001655|T121|ACTH|lab,
C0032343|T037|poisoning|
C1320226|T033|incubation period|
C1258666|T047|ganglion|
C1293131|T061|fusion|
C0008405|T123|choline|medication,
C0008405|T109|choline|medication,
C0008405|T121|choline|medication,
C0231221|T033|asymptomatic|
C0030956|T116|peptides|
C0017890|T123|glycine|medication,
C0017890|T116|glycine|medication,
C0017890|T121|glycine|medication,
C0006935|T122|capsule|
C0229665|T024|arterial blood|
C0001551|T121|Adjuvant|
C0001551|T129|Adjuvant|
C0042789|T040|vision|
C0790233|T197|distilled water|
C0790233|T121|distilled water|
C0301911|T044|complement fixation|lab,
C0035094|T116|renin|lab,
C0035094|T126|renin|lab,
C0028259|T020|nodules|
C0027697|T047|nephritis|diagnosis,
C0027697|T047|nephritis|diagnosis,problem,
C0015684|T109|fatty acid|
C0021853|T023|bowel|
C0024299|T191|lymphoma|diagnosis,
C0024299|T191|lymphoma|diagnosis,problem,
C0024204|T023|lymph node|
C0031727|T116|kinase|
C0031727|T126|kinase|
C0042196|T061|inoculations|
C0225336|T025|endothelial cells|
C0014136|T022|endocrine|
C0010137|T121|cortisone|medication,
C0010137|T125|cortisone|medication,
C0010137|T109|cortisone|medication,
C1623038|T047|cirrhosis|diagnosis,
C1623038|T047|cirrhosis|diagnosis,problem,
C0156543|T033|abortion|procedure,
C0014070|T047|encephalomyelitis|diagnosis,
C0014070|T047|encephalomyelitis|diagnosis,problem,
C1442959|T040|nutrition|
C0028351|T121|noradrenaline|lab,
C0028351|T121|noradrenaline|lab,medication,
C0028351|T109|noradrenaline|lab,
C0028351|T109|noradrenaline|lab,medication,
C0028351|T125|noradrenaline|lab,
C0028351|T125|noradrenaline|lab,medication,
C0524466|T029|intracranial|
C0012546|T047|diphtheria|immunization,
C0012546|T047|diphtheria|immunization,diagnosis,
C0012546|T047|diphtheria|immunization,diagnosis,problem,
C0565514|T061|compression|
C0023820|T116|lipoprotein|
C0023820|T123|lipoprotein|
C0020885|T023|ileum|
C0014898|T109|ester|
C0009637|T040|conception|
C0002059|T116|alkaline phosphatase|lab,
C0002059|T126|alkaline phosphatase|lab,
C0242692|T024|skeletal muscle|
C0546816|T041|persistence|
C0030054|T196|O2|lab,
C0030054|T196|O2|lab,treatment,
C0030054|T121|O2|lab,
C0030054|T121|O2|lab,treatment,
# C0006826|T191|malignancy|problem, JIRA/SANDS-173
C0013343|T130|dyes|
C0376259|T109|citrate|
C0376259|T121|citrate|
C0004461|T026|axon|
C0042210|T121|vaccines|
C0042210|T129|vaccines|
C0244104|T123|pyruvate|lab,
C0244104|T109|pyruvate|lab,
C0027021|T116|peroxidase|
C0027021|T126|peroxidase|
C0028606|T114|nucleic acid|
C0028606|T123|nucleic acid|
C0027061|T024|myocardium|
C0018494|T023|hair|
C0016169|T190|fistula|
C0015811|T023|femoral|
C0301642|T044|denaturation|
C0443985|T129|HCl|medication,
C0684271|T040|drinking|
C0032074|T041|planning|
C0027651|T191|neoplasms|
C0022116|T046|ischemia|
C0015450|T029|face|
C0687028|T023|ducts|
C0010709|T047|cysts|
C0205042|T023|coronary artery|
C0262950|T023|bones|
C0038435|T033|stressed|
C0332461|T033|plaque|
C0020835|T116|IgA|lab,
C0020835|T129|IgA|lab,
C0013879|T196|element|
C0282335|T023|respiratory tract|
C0023690|T061|ligation|
C0014520|T024|epidermis|
C0004096|T047|asthma|diagnosis,
C0004096|T047|asthma|diagnosis,problem,
C0344211|T061|supporting|
C0035078|T047|renal failure|diagnosis,
C0035078|T047|renal failure|diagnosis,problem,
C0028351|T121|norepinephrine|lab,
C0028351|T121|norepinephrine|lab,medication,
C0028351|T109|norepinephrine|lab,
C0028351|T109|norepinephrine|lab,medication,
C0028351|T125|norepinephrine|lab,
C0028351|T125|norepinephrine|lab,medication,
C0025289|T047|meningitis|diagnosis,
C0025289|T047|meningitis|diagnosis,problem,
C0015385|T023|limb|
C0022346|T046|jaundice|diagnosis,
C0022346|T046|jaundice|diagnosis,problem,
C0301872|T042|immune response|
C0016658|T037|fracture|diagnosis,
C0016658|T037|fracture|diagnosis,problem,
C0016504|T023|foot|
C0001473|T116|ATPase|
C0001473|T126|ATPase|
C0030946|T116|protease|
C0030946|T126|protease|
C0030946|T121|protease|
C0024530|T047|malaria|diagnosis,
C0024530|T047|malaria|diagnosis,problem,
C0039597|T023|testis|
C0004048|T040|Inhalation|
C0231239|T184|Fluctuations|
C0010654|T123|cysteine|medication,
C0010654|T116|cysteine|medication,
C0278134|T184|anaesthesia|procedure,
C0042963|T184|vomiting|problem,
C0700042|T029|ocular|
C1269575|T023|medulla|
C0024432|T025|macrophage|
C1140621|T029|leg|
C0014264|T131|endotoxin|
C0014264|T109|endotoxin|
C0013303|T023|duodenum|
C0040405|T060|CT|lab,
C0040405|T060|CT|lab,procedure,
C0003075|T196|anion|
C0026473|T025|monocytes|lab,
C0021493|T061|intraperitoneal injection|procedure,
C0018905|T059|hemagglutination|lab,
C0011991|T184|diarrhea|problem,
#C0006826|T191|cancers| JIRA/BIOMED-374
C0232804|T042|renal function|
C1314687|T033|sexes|
C0003873|T047|rheumatoid arthritis|diagnosis,
C0003873|T047|rheumatoid arthritis|diagnosis,problem,
C1961028|T033|oriented|
C0026724|T024|mucosal|
C0013227|T121|medication|
C0242184|T046|hypoxia|diagnosis,
C0242184|T046|hypoxia|diagnosis,problem,
C0016658|T037|fractures|
C0225328|T026|fibrils|
C0010294|T123|creatinine|lab,
C0010294|T109|creatinine|lab,
C0086881|T030|canal|
C0000833|T047|abscess|problem,
C0031208|T041|personality|
C0023317|T023|lens|
C0259862|T122|emulsion|
C0001455|T121|cyclic AMP|
C0001455|T123|cyclic AMP|
C0001455|T114|cyclic AMP|
C0332447|T190|anomalies|
C0037125|T196|silver|
C1963578|T061|releasing|
C0030125|T121|pass|
C0030125|T109|pass|
C0024090|T029|lumbar|
C0443235|T061|impulses|
C0185003|T061|closure|
C0225810|T029|bases|
C0162340|T041|understood|
C0456984|T033|testing|
C0441621|T060|sampling|
C0028630|T114|nucleotides|
C1510470|T040|motility|
C0022417|T030|joints|
C1265875|T020|disintegration|
C0070570|T121|phenol|medication,
C0070570|T109|phenol|medication,
C0017189|T022|gastrointestinal tract|
C0733758|T125|FSH|lab,
C0733758|T116|FSH|lab,
C0733758|T121|FSH|lab,
C0003962|T033|ascites|diagnosis,
C0003962|T033|ascites|diagnosis,problem,
C0002607|T121|ammonia|lab,
C0002607|T197|ammonia|lab,
C0032120|T123|plasma proteins|
C0032120|T116|plasma proteins|
C0030797|T023|pelvic|
C0020268|T121|cortisol|lab,
C0020268|T125|cortisol|lab,
C0020268|T109|cortisol|lab,
C0007004|T109|carbohydrates|
C0001804|T129|Agglutinin|
C0001418|T191|adenocarcinoma|diagnosis,
C0001418|T191|adenocarcinoma|diagnosis,problem,
C0037313|T040|sleep|
C0036429|T046|sclerosis|
C0524865|T061|reconstruction|
C0032120|T123|plasma protein|
C0032120|T116|plasma protein|
C0015967|T033|febrile|
C0012632|T041|discrimination|
C0231170|T033|disability|
C0010505|T197|cyanide|lab,
C0039259|T023|tail|
C0038179|T121|starch|
C0038179|T123|starch|
C0038179|T109|starch|
C0033497|T121|propranolol|medication,
C0033497|T109|propranolol|medication,
C0031715|T044|phosphorylation|
C0029939|T023|ovary|
C0027540|T042|necrotic|
C0018787|T023|hearts|
C0011980|T023|diaphragm|
C0005367|T197|bicarbonate|lab,
C0005367|T121|bicarbonate|lab,
C1140618|T023|arm|
C0000726|T029|abdomen|
C0041582|T047|ulcers|
C1879316|T061|transfusion|procedure,
C0443640|T116|specific antibody|
C0443640|T129|specific antibody|
C0013862|T059|polyacrylamide gel electrophoresis|
C0026549|T121|morphine|allergy,
C0026549|T121|morphine|allergy,medication,
C0026549|T109|morphine|allergy,
C0026549|T109|morphine|allergy,medication,
C0005778|T042|clotting|
C0005790|T059|clotting|
C0020517|T046|allergy|
C2584946|T033|alive|
C0001898|T123|alanine|medication,
C0001898|T116|alanine|medication,
C0001109|T116|acid phosphatase|lab,
C0001109|T126|acid phosphatase|lab,
C1704247|T030|peritoneal cavity|
C0030518|T023|Parathyroid|
C0017243|T122|gels|
C0949307|T121|formalin|
C0949307|T109|formalin|
C0949307|T131|formalin|
C0274281|T037|exposures|social,
C0001721|T041|affect|
C0036751|T109|5-hydroxytryptamine|lab,
C0036751|T123|5-hydroxytryptamine|lab,
C0036572|T184|seizures|problem,
C0026882|T045|mutation|
C0023516|T025|leucocyte|lab,
C0022742|T023|knee|
C0013819|T060|EEG|lab,
C0013819|T060|EEG|lab,procedure,
C0006104|T023|brains|
C0185023|T061|attachment|
C0014563|T109|adrenaline|lab,
C0014563|T109|adrenaline|lab,medication,
C0014563|T125|adrenaline|lab,
C0014563|T125|adrenaline|lab,medication,
C0014563|T121|adrenaline|lab,
C0014563|T121|adrenaline|lab,medication,
C0038128|T130|stain|
C1522449|T061|radiotherapy|treatment,
C0017649|T123|globulins|
C0017649|T116|globulins|
C0014898|T109|Esters|
C0013618|T121|EDTA|
C0013618|T109|EDTA|
C0003445|T121|antitoxin|
C0003445|T129|antitoxin|
C0033572|T023|prostate|
C0001002|T109|acetone|
C0001002|T121|acetone|
C0443343|T033|unstable|
C0087130|T033|uncertain|
C0036751|T109|serotonin|lab,
C0036751|T123|serotonin|lab,
C0032594|T121|polysaccharides|
C0032594|T109|polysaccharides|
C0026162|T197|mineral|
C0025474|T029|mesenteric|
C0000768|T019|malformations|
C0017817|T123|glutathione|medication,
C0017817|T116|glutathione|medication,
C0332853|T020|anastomosis|
C0677554|T061|anastomosis|
C0042214|T047|vaccinia|
C0332154|T033|Treated for|
C0040018|T121|thrombin|medication,
C0040018|T116|thrombin|medication,
C0040018|T126|thrombin|medication,
C0233324|T040|termed|
C0037638|T130|solvent|
C0031676|T123|phospholipid|
C0031676|T109|phospholipid|
C0026018|T059|Microscopic examination|
C0010709|T047|cyst|
C0010031|T023|cornea|
C0001407|T114|adenine|
C0001407|T123|adenine|
C3714552|T184|weakness|problem,
C0202231|T059|Thyroxine|lab,
C0202231|T059|Thyroxine|lab,medication,
C0040165|T121|thyroxine|lab,
C0040165|T121|thyroxine|lab,medication,
C0040165|T125|thyroxine|lab,
C0040165|T125|thyroxine|lab,medication,
C0040165|T116|thyroxine|lab,
C0040165|T116|thyroxine|lab,medication,
C0023689|T116|synthetase|
C0023689|T126|synthetase|
C0227952|T023|sheath|
C0015385|T023|extremities|
C0086140|T121|dextran|medication,
C0086140|T109|dextran|medication,
C0042027|T023|urinary tract|
C0038454|T047|stroke|diagnosis,
C0038454|T047|stroke|diagnosis,problem,
C3845714|T033|several days|
C0229992|T041|mind|
C0430389|T059|light microscopy|lab,
C0016945|T123|galactose|lab,
C0016945|T109|galactose|lab,
C1444662|T033|discontinued|
C1533591|T042|calcification|
C0004799|T024|basement membrane|
C0043250|T037|wounds|
C0450093|T033|very large|
C0038425|T195|streptomycin|medication,
C0038425|T109|streptomycin|medication,
C0030016|T116|reductase|
C0030016|T126|reductase|
C0017651|T023|pallidum|
C0026969|T024|myelin|
C2939419|T191|metastasis|
C0022864|T040|labor|
C0021368|T046|inflammatory reaction|problem,
C0018183|T025|granulocytes|lab,
C0017687|T121|glucagon|lab,
C0017687|T121|glucagon|lab,medication,
C0017687|T125|glucagon|lab,
C0017687|T125|glucagon|lab,medication,
C0017687|T116|glucagon|lab,
C0017687|T116|glucagon|lab,medication,
C0000983|T121|acetic acid|medication,
C0000983|T130|acetic acid|medication,
C0000983|T109|acetic acid|medication,
C0037995|T061|splenectomy|procedure,
C0031676|T123|phospholipids|
C0031676|T109|phospholipids|
C0235169|T184|excitability|
C0001122|T046|acidosis|problem,
C0041249|T121|tryptophan|medication,
C0041249|T123|tryptophan|medication,
C0041249|T116|tryptophan|medication,
C0441636|T061|shortening|
C0027651|T191|neoplasm|
C0023516|T025|leukocyte|lab,
C0031617|T123|lecithin|lab,
C0031617|T123|lecithin|lab,medication,
C0031617|T109|lecithin|lab,
C0031617|T109|lecithin|lab,medication,
C0031617|T121|lecithin|lab,
C0031617|T121|lecithin|lab,medication,
C0014563|T109|epinephrine|lab,
C0014563|T109|epinephrine|lab,medication,
C0014563|T125|epinephrine|lab,
C0014563|T125|epinephrine|lab,medication,
C0014563|T121|epinephrine|lab,
C0014563|T121|epinephrine|lab,medication,
C0010583|T121|cyclophosphamide|medication,
C0010583|T109|cyclophosphamide|medication,
C0007874|T023|cervix|
C0002792|T046|anaphylaxis|diagnosis,
C0002792|T046|anaphylaxis|diagnosis,problem,
C0041618|T060|ultrasound|procedure,
C0038774|T196|sulfur|
C0038774|T121|sulfur|
C0037868|T025|spermatozoa|
C0027749|T026|nerve fibers|
C0026255|T043|mitosis|
C0025202|T191|melanoma|diagnosis,
C0025202|T191|melanoma|diagnosis,problem,
C0225326|T121|fibre|
C0333288|T046|dissection|
C0012737|T061|dissection|
C0741847|T061|bypass|
C0043481|T196|zinc|lab,
C0043481|T196|zinc|lab,medication,
C0043481|T121|zinc|lab,
C0043481|T121|zinc|lab,medication,
C0039597|T023|testes|
C0199176|T061|prophylaxis|
C0030305|T047|pancreatitis|diagnosis,
C0030305|T047|pancreatitis|diagnosis,problem,
C0022262|T196|isotope|
C0021400|T047|influenzae|
C0344441|T059|histology|lab,
C0344441|T059|histology|lab,procedure,
C0019602|T123|histidine|medication,
C0019602|T116|histidine|medication,
C0019602|T121|histidine|medication,
C0016327|T197|fluoride|medication,
C0016327|T121|fluoride|medication,
C0003018|T121|angiotensin|
C0003018|T123|angiotensin|
C0003018|T116|angiotensin|
C0002932|T121|anesthetic|
C0229667|T024|venous blood|
C0243026|T047|septicemia|diagnosis,
C0243026|T047|septicemia|diagnosis,problem,
C0441610|T061|reductions|
C0443235|T061|impulse|
C0008354|T047|cholera|diagnosis,
C0008354|T047|cholera|diagnosis,problem,
C0230445|T029|calves|
C0003467|T048|anxiety|diagnosis,
C0003467|T048|anxiety|diagnosis,problem,
C0042760|T026|virus particles|
C0443640|T116|Specific antibodies|
C0443640|T129|Specific antibodies|
C0033572|T023|prostatic|
C0031180|T197|peroxide|
C0409974|T047|Lupus|diagnosis,
C0409974|T047|Lupus|diagnosis,problem,
C0032300|T047|lobar pneumonia|diagnosis,
C0032300|T047|lobar pneumonia|diagnosis,problem,
C0574032|T061|infusions|
C0040426|T023|teeth|
C0028429|T023|nose|
C0027950|T025|neutrophils|lab,
C0023764|T116|lipase|lab,
C0023764|T126|lipase|lab,
C0023764|T121|lipase|lab,
C0015385|T023|limbs|
C0019721|T116|HLA|
C0019721|T129|HLA|
C1290905|T033|discrepancy|
C0201682|T059|chemistry|
C1510420|T190|cavities|problem,
C0003075|T196|anions|
C0002620|T130|ammonium sulfate|
C0002620|T197|ammonium sulfate|
C0002508|T109|amines|
C0001459|T123|ADP|
C0001459|T114|ADP|
C0040284|T059|tissue cultures|
C0205400|T033|thickening|
C0037638|T130|solvents|
C0027950|T025|polymorphonuclear leucocytes|lab,
C0023185|T041|learning|
C0019080|T046|hemorrhages|
C0017725|T123|Dextrose|medication,
C0017725|T109|Dextrose|medication,
C0017725|T121|Dextrose|medication,
C0277786|T033|complaints|
C0003968|T121|Ascorbic acid|medication,
C0003968|T127|Ascorbic acid|medication,
C0003968|T109|Ascorbic acid|medication,
C0425382|T033|adopted|
C0001430|T191|adenoma|diagnosis,
C1444777|T033|splitting|
C0037506|T121|sodium dodecyl sulfate|
C0037506|T109|sodium dodecyl sulfate|
C0037506|T122|sodium dodecyl sulfate|
C0475463|T116|neutralizing antibodies|
C0475463|T129|neutralizing antibodies|
C0023820|T116|lipoproteins|
C0023820|T123|lipoproteins|
C0220839|T123|glutamate|medication,
C0220839|T116|glutamate|medication,
C0016030|T025|fibroblast|
C0002508|T109|amine|
C0458827|T023|airway|
C0039614|T047|tetanus|immunization,
C0039614|T047|tetanus|immunization,diagnosis,
C0039614|T047|tetanus|immunization,diagnosis,problem,
C0040165|T121|T4|lab,
C0040165|T125|T4|lab,
C0040165|T116|T4|lab,
C0228243|T030|T4|lab,
C0475371|T033|T4|lab,
C0075429|T121|succinate|
C0075429|T109|succinate|
C0035542|T116|ribonuclease|
C0035542|T126|ribonuclease|
C0025424|T131|mercury|lab,
C0025424|T196|mercury|lab,
C0019080|T046|haemorrhage|
C0011041|T131|DDT|
C0011041|T109|DDT|
C1261287|T046|constriction|
C0008260|T123|chlorophyll|
C0008260|T109|chlorophyll|
C0007585|T059|cell cultures|
C0007430|T061|catheterization|
C0004153|T047|atherosclerosis|diagnosis,
C0004153|T047|atherosclerosis|diagnosis,problem,
C0002940|T047|aneurysm|diagnosis,
C0002940|T047|aneurysm|diagnosis,problem,
C1273517|T033|used by|
C0041471|T047|typhus|diagnosis,
C0041471|T047|typhus|diagnosis,problem,
C0034991|T061|rehabilitation|treatment,
C1444783|T033|instability|
C0262926|T033|histories|
C0019552|T023|hip|
C0017968|T116|glycoprotein|
C0017968|T123|glycoprotein|
C0022663|T023|glomeruli|
C0014894|T116|esterase|
C0014894|T126|esterase|
C0013443|T023|ears|
C0440049|T130|spores|
C0034052|T023|pulmonary artery|
C0694756|T030|intrauterine|
C0020364|T116|hydroxylase|
C0020364|T126|hydroxylase|
C0018801|T047|heart failure|diagnosis,
C0018801|T047|heart failure|diagnosis,problem,
C0060520|T130|fluorescein|
C0060520|T109|fluorescein|
C0015852|T044|fermentation|
C0001617|T121|corticosteroids|
C0001617|T125|corticosteroids|
C0001617|T109|corticosteroids|
C0006142|T191|breast cancer|diagnosis,
C0006142|T191|breast cancer|diagnosis,problem,
C0005773|T025|blood cell|
C0005437|T109|bilirubin|lab,
C0005437|T123|bilirubin|lab,
C0279516|T195|antibacterial|
C0000924|T037|accident|
C0042890|T127|vitamins|
C0042890|T109|vitamins|
C0042890|T121|vitamins|
C1268443|T025|normal cells|
C0229889|T023|lymphatics|
C0184898|T061|Incision|
C0991568|T122|drops|
C0441513|T061|construction|
C0004372|T046|autolysis|
C0000833|T047|abscesses|
C0036825|T123|serum proteins|
C0036825|T116|serum proteins|
C0026837|T184|rigid|
C0220903|T109|purine|
C0032861|T122|powder|
C0031453|T123|phenylalanine|medication,
C0031453|T116|phenylalanine|medication,
C0031453|T121|phenylalanine|medication,
C0031307|T025|phagocytes|
C0549099|T033|perforation|
C0029219|T026|organelles|
C0026882|T045|mutations|
C0021107|T061|insertion|
C0232197|T047|fibrillation|
C0231800|T042|expiratory|
C0011164|T046|degenerative changes|diagnosis,
C0011164|T046|degenerative changes|diagnosis,problem,
C1265875|T020|decay|
C0008168|T195|chloramphenicol|medication,
C0008168|T109|chloramphenicol|medication,
C0007412|T123|catecholamines|lab,
C0007412|T121|catecholamines|lab,
C0028778|T046|blocks|
C0042839|T109|vitamin A|lab,
C0042839|T109|vitamin A|lab,medication,
C0042839|T127|vitamin A|lab,
C0042839|T127|vitamin A|lab,medication,
C0042839|T121|vitamin A|lab,
C0042839|T121|vitamin A|lab,medication,
C0040549|T123|toxins|
C0040549|T131|toxins|
C0032346|T131|poison|
C0233174|T033|parallelism|
C0023038|T061|laparotomy|procedure,
C0021966|T197|iodide|
C0020746|T197|ice|
C0020268|T121|hydrocortisone|medication,
C0020268|T125|hydrocortisone|medication,
C0020268|T109|hydrocortisone|medication,
C0011603|T047|dermatitis|diagnosis,
C0011603|T047|dermatitis|diagnosis,problem,
C0007603|T026|cell membranes|
C0036720|T123|serine|medication,
C0036720|T116|serine|medication,
C0036720|T121|serine|medication,
C0035953|T056|running|
C0033706|T121|prothrombin|
C0033706|T123|prothrombin|
C0033706|T116|prothrombin|
C1305923|T116|polypeptides|
C0176996|T061|nephrectomy|procedure,
C0035696|T123|mRNA|
C0035696|T114|mRNA|
C0025746|T121|Methylene Blue|
C0025746|T130|Methylene Blue|
C0025746|T109|Methylene Blue|
C0022925|T042|lactation|
C0020259|T130|hydrochloric acid|
C0020259|T197|hydrochloric acid|
C0017007|T116|gamma globulin|lab,
C0017007|T129|gamma globulin|lab,
C0259862|T122|emulsions|
C0231303|T041|distress|
C0700124|T033|dilated|
C0010957|T037|damaged|
C0010682|T123|cystine|medication,
C0010682|T116|cystine|medication,
C0010682|T121|cystine|medication,
C0007765|T023|cerebellum|
C0699900|T040|catabolism|
C0440746|T024|brain tissue|
C0042479|T131|venom|
C0037303|T023|skull|
C0026828|T042|innervation|
C0020944|T061|immobilization|
C0014876|T023|esophagus|
C0009871|T121|contraceptives|
C0007776|T023|cerebral cortex|
C0007412|T123|catecholamine|
C0007412|T121|catecholamine|
C0007367|T116|catalase|
C0007367|T126|catalase|
C0043395|T047|yellow fever|diagnosis,
C0043395|T047|yellow fever|diagnosis,problem,
C1262477|T033|weight loss|problem,
C0041980|T123|uric acid|lab,
C0041980|T109|uric acid|lab,
C0040160|T121|TSH|lab,
C0040160|T125|TSH|lab,
C0040160|T116|TSH|lab,
C0040732|T061|transplants|
C0332835|T024|transplants|
C0040732|T061|transplant|
C0332835|T024|transplant|
C0040329|T121|tobacco|social,
C0040329|T131|tobacco|social,
C0040329|T109|tobacco|social,
C1278878|T023|thyroid gland|
C0039597|T023|testicle|
C0813207|T061|shunt|
C1442858|T033|shunt|
C0035553|T026|ribosomes|
C1304757|T034|protein concentration|
C0007603|T026|plasma membranes|
C0029939|T023|ovaries|
C0027497|T184|nausea|problem,
C0025260|T041|memory|
C0022949|T123|lactose|
C0022949|T109|lactose|
C0061472|T123|glutamic acid|medication,
C0061472|T116|glutamic acid|medication,
C0061472|T121|glutamic acid|medication,
C0017526|T025|giant cells|
C0016564|T131|formaldehyde|
C0016564|T109|formaldehyde|
C0016564|T121|formaldehyde|
C0200069|T060|fertility|
C0015895|T040|fertility|
C0011175|T047|dehydration|problem,
C0010286|T123|creatine|medication,
C0010286|T116|creatine|medication,
C1704638|T122|cone|
C0007465|T033|cause of death|
C0036774|T123|bovine serum albumin|
C0036774|T116|bovine serum albumin|
C0332447|T190|anomaly|
C0001811|T040|aging|
C0043227|T057|worked|
C0041004|T123|triglyceride|
C0041004|T109|triglyceride|
C0040578|T023|trachea|
C0600688|T037|toxic effects|
C0039231|T046|tachycardia|problem,
C0038128|T130|stains|
C1306645|T060|radiographs|
C0429627|T033|oxygen uptake|
C1269830|T033|margin|
C0162429|T047|malnutrition|diagnosis,
C0162429|T047|malnutrition|diagnosis,problem,
C0022378|T023|jejunum|
C0020649|T033|hypotension|diagnosis,
C0020649|T033|hypotension|diagnosis,problem,
C2981153|T033|focusing|
C0014939|T121|estrogens|
C0014939|T125|estrogens|
C0014939|T109|estrogens|
C0202006|T059|estrogens|
C0011900|T033|diagnoses|
C0152060|T061|cutting|
C0700198|T046|aspiration|
C0349707|T061|aspiration|
C0332461|T033|plaques|
C0013604|T033|oedema|problem,
C0736268|T023|liver tissue|
C0013922|T046|embolism|
C0002871|T047|anaemia|diagnosis,
C0002871|T047|anaemia|diagnosis,problem,
C0002006|T121|aldosterone|lab,
C0002006|T125|aldosterone|lab,
C0002006|T109|aldosterone|lab,
C1705480|T121|vasopressin|lab,
C1705480|T121|vasopressin|lab,medication,
C1705480|T116|vasopressin|lab,
C1705480|T116|vasopressin|lab,medication,
C1705480|T125|vasopressin|lab,
C1705480|T125|vasopressin|lab,medication,
C0041609|T059|ultracentrifugation|
C3887532|T046|ulceration|
C0031354|T023|throat|
C0039082|T047|syndromes|
C0037949|T023|spine|