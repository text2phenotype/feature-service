C0031117|Peripheral Neuropathy
C0027868|Neuromuscular Disease
C0027868|Neuromuscular Diseases
C0027868|Myoneural disorders
C0027868|neuromuscular disorder
C0027868|Myoneural disorders, unspecified
C0027868|Myoneural disorder, unspecified
C0027868|NEUROMUSCULAR DIS
C0027868|Combined disorder of muscle AND peripheral nerve
C0027868|myoneural disorder
C0027868|neuromuscular diseases (diagnosis)
C0027868|myoneural disorder (diagnosis)
C0027868|Neuromuscular disorders
C0027868|Myoneural disorders NOS
C0027868|Neuromuscular Diseases [Disease/Finding]
C0027868|Combined disorder of muscle AND peripheral nerve (disorder)
C0027868|Myoneural disorder NOS
C0027868|Myoneural disorder NOS (disorder)
C0027868|Neuromyopathy
C0027868|Neuromuscular disorder NOS
C0027868|Neuromyopathy (disorder)
C0027868|disease (or disorder); myoneural
C0027868|disease (or disorder); neuromuscular system
C0027868|Myoneural disorder, NOS
C0027868|Neuromuscular disease, NOS
C0027868|Neuromyopathy, NOS
C0027868|Combined disorder of muscle AND peripheral nerve [Ambiguous]
C0029132|Lesion, Neural-Optical
C0029132|Lesions, Neural-Optical
C0029132|Neural Optical Lesion
C0029132|Neural-Optical Lesions
C0029132|Optic Nerve Disease
C0029132|Optic Nerve Diseases
C0029132|optic nerve disorder
C0029132|SECOND CRANIAL NERVE DIS
C0029132|OPTIC NERVE DIS
C0029132|CRANIAL NERVE II DIS
C0029132|Disorder of the optic nerve
C0029132|disorder of optic nerve (diagnosis)
C0029132|disorder of optic nerve
C0029132|Neuropathies, Optic
C0029132|Neuropathy, Optic
C0029132|Optic Neuropathies
C0029132|Second Cranial Nerve Disorder
C0029132|Second Cranial Nerve Diseases
C0029132|Cranial Nerve II Disorder
C0029132|Neural-Optical Lesion
C0029132|Optic Nerve Diseases [Disease/Finding]
C0029132|Optic Neuropathy
C0029132|Cranial Nerve II Diseases
C0029132|Disorders of the IInd cranial nerve
C0029132|Disorders of the second nerve
C0029132|Optic nerve disorders
C0029132|Disorder of cranial nerve 2
C0029132|Disorder of second cranial nerve
C0029132|Optic nerve--Diseases
C0029132|Optic nerve disorder NOS
C0029132|Disorder of optic nerve (disorder)
C0029132|cranial nerve; disorder, second (optic)
C0029132|disease (or disorder); cranial nerve, second (optic)
C0029132|disease (or disorder); nerve, optic
C0029132|disease (or disorder); optic nerve
C0029132|n.opticus; disorder
C0029132|optic nerve; disorder
C0029132|Disorder of optic nerve, NOS
C0007286|Carpal Tunnel Syndrome
C0007286|Carpal Tunnel Syndromes
C0007286|Syndromes, Carpal Tunnel
C0007286|Syndrome, Carpal Tunnel
C0007286|CTS1
C0007286|CTS (carpal tunnel syndrome)
C0007286|carpal tunnel syndrome (diagnosis)
C0007286|Compression Neuropathy, Carpal Tunnel
C0007286|Median Neuropathy, Carpal Tunnel
C0007286|Carpal Tunnel Syndrome [Disease/Finding]
C0007286|Entrapment Neuropathy, Carpal Tunnel
C0007286|Carpal tunnel syndrome, unspecified upper limb
C0007286|Amyotrophy, Thenar, Of Carpal Origin
C0007286|Median nerve entrapment
C0007286|Carpal tunnel syndrome (disorder)
C0007286|CTS - Carpal tunnel syndrome
C0007286|CTS
C0007286|Distal median nerve entrapment
C0007286|Distal median nerve compression
C0007286|Median nerve compression
C0007286|Carpal canal
C0007286|Carpal tunnel
C0007286|Median nerve entrapment (disorder)
C0007286|carpal tunnel; syndrome
C0007286|compression; median nerve (in carpal tunnel)
C0007286|entrapment; neuropathic, nerve, median
C0007286|n.medianus; compression (in carpal tunnel)
C0007286|neuropathy; entrapment, nerve, median
C0007286|syndrome; carpal tunnel
C0007286|carpal tunnel median neuropathy
C0007286|Carpel tunnel syndrome
C0007286|Syndrome carpel tunnel
C0011882|Diabetic Neuropathies
C0011882|Neuropathies, Diabetic
C0011882|Diabetes with neurological manifestations
C0011882|Diabetic Neuropathy
C0011882|Neuropathy, Diabetic
C0011882|Diabetic Neuropathies [Disease/Finding]
C0011882|Neuropathy;diabetic
C0011882|Neuropathy - diabetic
C0011882|Diabetes + neuropathy
C0011882|Diabetic neuropathy (disorder)
C0011882|Diabetes mellitus with neuropathy
C0011882|Diabetes mellitus with neurological manifestation
C0011882|Diabetes mellitus NOS with neurological manifestation (disorder)
C0011882|Diabetes mellitus NOS with neurological manifestation
C0011882|neuropathy; diabetes (manifestation)
C0011882|Diabetic neuropathy (disorder) [Ambiguous]
C0015469|Facial Paralysis
C0015469|Paralyses, Facial
C0015469|Paralysis, Facial
C0015469|Facial Palsies
C0015469|Palsies, Facial
C0015469|Palsy, Facial
C0015469|Bell's Palsy
C0015469|Facial palsy
C0015469|Facial Paralysis [Disease/Finding]
C0015469|Palsy;facial
C0015469|Facial nerve paralysis
C0015469|Facial nerve palsy
C0015469|Facial nerve palsy (cranial nerve VII)
C0015469|Seventh nerve palsy
C0015469|VII nerve palsy
C0015469|Seventh nerve paralysis
C0015469|Facial nerve paralysis (disorder)
C0015469|Facial nerve palsies
C0015469|Paralysis Of Facial Nerve
C0015469|Nerve Paralysis, Facial
C0015469|Paralysis facial
C0015469|Facial palsy (disorder)
C0015469|facial; paralysis
C0015469|paralysis; facial nerve
C0015469|paralysis; facial
C0015469|Facial nerve paralysis, NOS
C0015469|VII th nerve palsy
C0015469|Palsy;VII nerve
C0030443|Familial Periodic Paralyses
C0030443|Paralyses, Familial Periodic
C0030443|Paralysis, Familial Periodic
C0030443|Periodic Paralyses, Familial
C0030443|Familial periodic paralysis
C0030443|familial periodic paralysis syndrome (diagnosis)
C0030443|familial periodic paralysis syndrome
C0030443|Paralyses, Familial Periodic [Disease/Finding]
C0030443|Periodic Paralysis, Familial
C0030443|Familial periodic paralysis (disorder)
C0030443|Paralysis periodic
C0030443|Cavarre disease
C0030443|Familial myoplegia
C0030443|Familial recurrent paralysis
C0030443|Myoplegic dystrophy
C0030443|Periodic myotonia
C0030443|paralysis; periodic
C0030443|periodic; paralysis
C0030443|Familial periodic paralysis, NOS
C0030443|Periodic paralysis
C0030443|Familial periodic paralysis (disorder) [Ambiguous]
C0027813|Neuritides
C0027813|Neuritis
C0027813|Neuritis, NOS
C0027813|neuritis (diagnosis)
C0027813|Neuritis -RETIRED-
C0027813|Neuritides, Peripheral
C0027813|Peripheral Neuritides
C0027813|Peripheral Neuritis
C0027813|Neuritis [Disease/Finding]
C0027813|Neuritis, Peripheral
C0027813|Neuritis;peripheral
C0027813|Neuritis (disorder)
C0027813|Neuritis unspecified
C0027813|Neuritis unspecified (disorder)
C0027813|Peripheral neuritis NOS
C0027813|Neuritis NOS
C0027813|Neuritis peripheral
C0027813|Peripheral neuritis (disorder)
C0027813|neuritis; peripheral
C0027813|peripheral; neuritis
C0027813|Peripheral neuritis, NOS
C0036396|Sciatica
C0036396|sciatica (diagnosis)
C0036396|Ischias
C0036396|Neuralgias, Sciatic
C0036396|Sciatic Neuralgias
C0036396|Sciatica, unspecified side
C0036396|Sciatic Neuralgia
C0036396|Sciatica [Disease/Finding]
C0036396|Neuralgia, Sciatic
C0036396|Sciatia
C0036396|Sciatica (disorder)
C0036396|Ischialgia
C0036396|Cotugno's disease
C0036396|Neuralgia-neuritis of sciatic nerve
C0036396|Sciatica neuralgia
C0036396|Neuralgia or neuritis of sciatic nerve
C0039621|Tetanies
C0039621|Tetany
C0039621|[D]Tetany (context-dependent category)
C0039621|[D]Tetany NOS (context-dependent category)
C0039621|tetany (physical finding)
C0039621|fingers and wrists curl up (symptom)
C0039621|fingers and wrists curl up
C0039621|Tetany [Disease/Finding]
C0039621|[D]Tetany (situation)
C0039621|[D]Tetany NOS
C0039621|Tetany (finding)
C0039621|[D]Tetany NOS (situation)
C0039621|[D]Tetany
C0039621|Tetany (disorder)
C0039621|Tetany, NOS
C0039621|Tetany [Ambiguous]
C0040997|Fothergill's neuralgia
C0040997|Neuralgias, Trigeminal
C0040997|Trigeminal Neuralgia
C0040997|Trigeminal Neuralgias
C0040997|Neuralgia, Trigeminal
C0040997|FOTHERGILL DIS
C0040997|tic douloureux
C0040997|trifocal neuralgia
C0040997|Tic doloreux
C0040997|Disease, Fothergill
C0040997|Neuralgia, Epileptiform
C0040997|Epileptiform Neuralgias
C0040997|Neuralgias, Epileptiform
C0040997|Neuralgia, Trifacial
C0040997|Neuralgias, Trifacial
C0040997|Trifacial Neuralgias
C0040997|Fothergill Disease
C0040997|Trifacial Neuralgia
C0040997|Trigeminal Neuralgia [Disease/Finding]
C0040997|Epileptiform Neuralgia
C0040997|TN
C0040997|Tic Douleureux
C0040997|Trigeminal neuralgia NOS
C0040997|Trigeminal neuralgia [no drugs here] (disorder)
C0040997|Trigeminal neuralgia [no drugs here]
C0040997|Trigeminal neuralgia NOS (disorder)
C0040997|Trigeminal neuralgia (disorder)
C0040997|Trigeminal neuralgia (diagnosis)
C0040997|Neuralgia trigeminal
C0040997|TN - Trigeminal neuralgia
C0040997|Fothergill; neuralgia
C0040997|Fothergill; trigeminal neuralgia
C0040997|cranial nerve; neuralgia, fifth or trigeminal
C0040997|douloureux; tic
C0040997|neuralgia; Fothergill
C0040997|neuralgia; cranial nerve, fifth or trigeminal
C0040997|neuralgia; trifacial
C0040997|neuralgia; trigeminal
C0040997|pain; trigeminal
C0040997|tic; douloureux
C0040997|trifacial; neuralgia
C0040997|trigeminal neuralgia; Fothergill
C0040997|trigeminal; neuralgia
C0040997|trigeminal; pain
C0040997|Trigeminal neuralgia, NOS
C0040997|Tic Doloureux
C0596694|hereditary peripheral nervous system disorder
C0151313|Peripheral sensory neuropathy
C0151313|Sensory neuropathy
C0151313|Peripheral neuropathy, sensory
C0151313|Sensory peripheral neuropathies
C0151313|Sensory peripheral neuropathy
C0151313|Sensory neuropathy (disorder)
C0027796|Neuralgias
C0027796|Neuralgia
C0027796|Neuralgia, NOS
C0027796|neuralgia (diagnosis)
C0027796|Neuralgia -RETIRED-
C0027796|Neurodynias
C0027796|Neuralgia [Disease/Finding]
C0027796|Neurodynia
C0027796|Neuropathic Pains
C0027796|Pains, Neuropathic
C0027796|Pain, Neuropathic
C0027796|Neuropathic Pain
C0027796|Neuralgia (disorder)
C0027796|Neuralgia unspecified
C0027796|Neuralgia unspecified (disorder)
C0027796|neuralgia (symptom)
C0027796|Neuralgia NOS
C0235025|Peripheral motor neuropathy
C0235025|Motor neuropathy
C0235025|Motor Neuritides
C0235025|Motor Neuritis
C0235025|Neuritides, Motor
C0235025|Motor peripheral neuropathy
C0235025|Neuritis motor
C0235025|Neuritis, Motor
C0235025|Peripheral motor neuropathy (disorder)
C0085677|Alcoholic polyneuropathy
C0085677|ALCOHOL IND POLYNEUROPATHY
C0085677|ALCOHOL IND PERIPHERAL NEUROPATHY
C0085677|PERIPHERAL NEUROPATHY ALCOHOL IND
C0085677|ALCOHOL RELAT POLYNEUROPATHY
C0085677|ALCOHOL RELAT AUTONOMIC POLYNEUROPATHY
C0085677|Alcohol-induced polyneuropathy -RETIRED-
C0085677|alcoholic polyneuropathy (diagnosis)
C0085677|Polyneuropathy alcoholic
C0085677|Alcohol-Related Autonomic Polyneuropathies
C0085677|Autonomic Polyneuropathies, Alcohol-Related
C0085677|Polyneuropathies, Alcohol-Related Autonomic
C0085677|Alcohol Related Autonomic Polyneuropathy
C0085677|Autonomic Polyneuropathy, Alcohol-Related
C0085677|Polyneuropathy, Alcohol-Related Autonomic
C0085677|Alcohol Induced Peripheral Neuropathy
C0085677|Alcohol-Induced Peripheral Neuropathies
C0085677|Neuropathies, Alcohol-Induced Peripheral
C0085677|Neuropathy, Alcohol-Induced Peripheral
C0085677|Peripheral Neuropathies, Alcohol-Induced
C0085677|Peripheral Neuropathy, Alcohol Induced
C0085677|Alcohol-Induced Polyneuropathies
C0085677|Polyneuropathies, Alcohol-Induced
C0085677|Alcohol Induced Polyneuropathy
C0085677|Polyneuropathy, Alcohol-Induced
C0085677|Alcohol-Related Polyneuropathies
C0085677|Polyneuropathies, Alcohol-Related
C0085677|Alcohol Related Polyneuropathy
C0085677|Polyneuropathy, Alcohol-Related
C0085677|Alcoholic Neuropathies
C0085677|Alcoholic Neuropathy
C0085677|Neuropathies, Alcoholic
C0085677|Alcoholic Polyneuritides
C0085677|Alcoholic Polyneuritis
C0085677|Polyneuritides, Alcoholic
C0085677|Alcoholic Polyneuropathies
C0085677|Polyneuropathies, Alcoholic
C0085677|Neuropathy, Alcoholic
C0085677|Polyneuritis, Alcoholic
C0085677|Polyneuropathy, Alcoholic
C0085677|Alcoholic Neuropathy [Disease/Finding]
C0085677|Alcohol-Induced Peripheral Neuropathy
C0085677|Alcohol-Induced Polyneuropathy
C0085677|Peripheral Neuropathy, Alcohol-Induced
C0085677|Alcohol-Related Autonomic Polyneuropathy
C0085677|Alcohol-Related Polyneuropathy
C0085677|Neuropathy;alcoholic
C0085677|Alcohol-induced polyneuropathy (disorder)
C0085677|Alcohol-related polyneuropathy (disorder)
C0085677|Alcoholic peripheral neuropathy
C0085677|Alcoholic polyneuropathy (disorder)
C0085677|polyneuropathy; alcoholic
C0085677|polyneuropathy; alcohol
C0085677|alcohol; polyneuropathy
C0393842|Polyneuropathy in neoplastic disease
C0393842|malignant neoplasm; polyneuropathy (etiology)
C0393842|malignant neoplasm; polyneuropathy (manifestation)
C0393842|neoplasm; polyneuropathy (manifestation)
C0393842|polyneuropathy; malignant neoplasm (etiology)
C0393842|polyneuropathy; malignant neoplasm (manifestation)
C0393842|polyneuropathy; neoplasm (manifestation)
C0270932|Polyneuropathy in malignant disease
C0270932|PERIPHERAL NEUROPATHY PARANEOPL
C0270932|PARANEOPL POLYNEUROPATHY
C0270932|NEUROPATHY PARANEOPL
C0270932|POLYNEUROPATHY PARANEOPL
C0270932|PARANEOPL PERIPHERAL NEUROPATHY
C0270932|PARANEOPL NEUROPATHY
C0270932|polyneuropathy due to malignant disease (diagnosis)
C0270932|polyneuropathy due to malignant disease
C0270932|Neuropathies, Paraneoplastic
C0270932|Paraneoplastic Neuropathies
C0270932|Neuropathies, Paraneoplastic Peripheral
C0270932|Neuropathy, Paraneoplastic Peripheral
C0270932|Paraneoplastic Peripheral Neuropathies
C0270932|Peripheral Neuropathies, Paraneoplastic
C0270932|Paraneoplastic Polyneuropathies
C0270932|Polyneuropathies, Paraneoplastic
C0270932|Paraneoplastic Polyneuropathy
C0270932|Neuropathy in malig dis
C0270932|Paraneoplastic Neuropathy
C0270932|Neuropathy, Paraneoplastic
C0270932|Paraneoplastic Peripheral Neuropathy
C0270932|Polyneuropathy, Paraneoplastic
C0270932|Paraneoplastic Polyneuropathy [Disease/Finding]
C0270932|Peripheral Neuropathy, Paraneoplastic
C0270932|Paraneoplastic peripheral neuropathy (disorder)
C0270932|Carcinomatous neuropathy
C0270932|Polyneuropathy in malignancy
C0270932|Carcinomatous peripheral neuropathy
C0270932|Paraneoplastic neuropathy (disorder)
C0859672|Other hereditary and idiopathic peripheral neuropathy
C0859672|Hereditary and idiopathic peripheral neuropathy, other
C0859673|Unspecified hereditary and idiopathic peripheral neuropathy
C0859673|Idio periph neurpthy NOS
C0477394|Other specified polyneuropathies
C0477394|[X]Other specified polyneuropathies
C0477394|[X]Other specified polyneuropathies (disorder)
C0494489|Mononeuropathies of lower limb
C0494489|Mononeuropathy of lower limb, unspecified
C0494489|Unspecified mononeuropathy of unspecified lower limb
C0494489|Unspecified mononeuropathy of lower limb
C0494489|Mononeuropathy of lower limb (disorder)
C0494489|Mononeuropathy of lower limb
C0154762|Polyneuropathy due to drugs
C0154762|Drug-induced polyneuropathy
C0154762|drug-induced polyneuropathy (diagnosis)
C0154762|Neuropathy due to drugs
C0154762|Polyneuropathy due to drug (disorder)
C0154762|Polyneuropathy caused by drug (disorder)
C0154762|Polyneuropathy caused by drug
C0154762|Drug-related polyneuropathy
C0154762|Polyneuropathy due to drug
C0154762|Polyneuropathy due to drug, NOS
C0494518|Autonomic neuropathy in endocrine and metabolic diseases
C0494518|neuropathy; peripheral, autonomic, in metabolic disease (manifestation)
C0235023|Neuritis bulbar
C0235026|Neuritides, Sensory
C0235026|Sensory Neuritides
C0235026|Sensory Neuritis
C0235026|Neuritis sensory
C0235026|Neuritis, Sensory
C0235919|Nerve root liaison
C0235919|Nerve root lesion
C0235919|Nerve root lesion NOS
C0238309|Ischaemic neuropathy
C0238309|Ischemic neuropathy
C0238309|Ischaemic peripheral neuropathy
C0238309|Ischemic neuropathy (disorder)
C0238309|Ischemic peripheral neuropathy (disorder)
C0238309|Ischemic peripheral neuropathy
C0393807|CMT6
C0393807|Hereditary motor and sensory neuropathy with optic atrophy (disorder)
C0393807|HMSN VI
C0393807|Peripheral Neuropathy And Optic Atrophy
C0393807|Charcot-Marie-Tooth Disease, Type 6
C0393807|HMSN6
C0393807|Hereditary Motor And Sensory Neuropathy VI
C0393807|Hereditary motor and sensory neuropathy with optic atrophy
C0393807|hereditary motor and sensory neuropathy with optic atrophy (diagnosis)
C0393807|NEUROPATHY, HEREDITARY MOTOR AND SENSORY, TYPE VI
C0393807|HSMN6
C0393807|Hereditary motor and sensory neuropathy type VI
C0393807|Hereditary motor-sensory neuropathy with optic atrophy
C0393807|Hereditary motor-sensory neuropathy, type VI
C0393807|Hereditary sensory and motor neuropathy, type VI
C0392553|hereditary peripheral neuropathy (diagnosis)
C0392553|hereditary peripheral neuropathy
C0392553|Hered periph neuropathy
C0392553|Hereditary peripheral neuropathy NOS
C0392553|Hereditary peripheral neuropathy NOS (disorder)
C0392553|Peripheral neuropathy hereditary
C0392553|Hereditary peripheral neuropathy (disorder)
C0392553|Hereditary peripheral neuropathy, NOS
C0154690|Idiopathic peripheral autonomic neuropathy
C0154690|idiopathic peripheral autonomic neuropathy (diagnosis)
C0154690|Idiopathic peripheral autonomic neuropathy NOS
C0154690|Idiopathic peripheral autonomic neuropathy (disorder)
C0154690|Idiopathic peripheral autonomic neuropathy NOS (disorder)
C0154690|neuropathy; peripheral, autonomic, idiopathic
C0154754|Hereditary and idiopathic peripheral neuropathy
C0154754|Hereditary and idiopathic neuropathy
C0154754|Hereditary and idiopathic neuropathy, unspecified
C0154754|Hereditary and idiopathic peripheral neuropathy (disorder)
C0154691|Peripheral autonomic neuropathy in disorders classified elsewhere
C0154691|Aut neuropthy in oth dis
C0154757|Other specified idiopathic peripheral neuropathy
C0154757|Idio periph neurpthy NEC
C0041848|Unspecified idiopathic peripheral neuropathy
C0041848|neuropathy; idiopathic
C0041848|Idiopathic Neuropathy
C0235024|Neuritis cranial
C0235024|Cranial neuritis
C0235024|Cranial neuritis (disorder)
C0235024|Cranial neuritis, NOS
C0235880|Mononeuritis of unspecified site
C0235880|Mononeuritis
C0235880|mononeuritis (diagnosis)
C0235880|Mononeuritides
C0235880|Mononeuritis NOS
C0235880|Mononeuritis of unspecified site NOS (disorder)
C0235880|Mononeuritis of unspecified site NOS
C0235880|Mononeuritis (disorder)
C0235880|Mononeuritis, NOS
C0270921|Axonal neuropathy
C0270921|Axonal neuropathy (disorder)
C0270921|Axonal neuropathy, NOS
C0001198|Acrodynia
C0001198|Feers Disease
C0001198|Swifts Disease
C0001198|FEERS DIS
C0001198|SWIFTS DIS
C0001198|PINK DIS
C0001198|SWIFT DIS
C0001198|FEER DIS
C0001198|Erythema, Acrodynic
C0001198|Childhood Mercurialism, Chronic
C0001198|Mercurialism, Chronic Childhood
C0001198|Childhood Mercurialisms, Chronic
C0001198|Chronic Childhood Mercurialisms
C0001198|Acrodynia [Disease/Finding]
C0001198|Swift Disease
C0001198|Chronic Childhood Mercurialism
C0001198|Swift's Disease
C0001198|Acrodynic Erythema
C0001198|Feer's Disease
C0001198|Feer Disease
C0001198|Pink Disease
C0001198|Selter's disease
C0001198|Swift-Feer disease
C0001198|Disease pink
C0001198|Erythredema polyneuropathy
C0001198|Bilderbeck's disease
C0001198|Acrodynia caused by mercury (disorder)
C0001198|Acrodynia caused by mercury poisoning
C0001198|Acrodynia due to mercury (disorder)
C0001198|Acrodynia due to mercury
C0001198|Acrodynia due to mercury poisoning
C0001198|Erythroedema polyneuropathy
C0001198|Acrodynia caused by mercury
C0001198|Swift
C0001198|Feer
C0001198|disease; pink
C0001198|erythredema; polyneuritic
C0001198|erythredema
C0001198|pink; disease
C0002768|Pain Insensitivity, Congenital
C0002768|Congenital Pain Insensitivity
C0002768|ANALGESIA CONGEN
C0002768|PAIN INSENSITIVITY CONGEN
C0002768|CONGEN PAIN INSENSITIVITY
C0002768|CONGEN ANALGESIA
C0002768|INSENSITIVITY CONGEN PAIN
C0002768|PAIN INDIFFERENCE CONGEN
C0002768|Congenital Pain Indifferences
C0002768|Congenital Indifference to Pain
C0002768|Analgesia, Congenital
C0002768|Congenital Analgesia
C0002768|Congenital Pain Indifference
C0002768|Insensitivity, Congenital Pain
C0002768|Pain Indifference, Congenital
C0002768|Pain Insensitivity, Congenital [Disease/Finding]
C0002768|Insensitivity To Pain, Congenital
C0002768|Channelopathy-Associated Insensitivity To Pain
C0002768|Congenital Insensitivity To Pain
C0002768|Congenital indifference to pain (finding)
C0002768|Congenital pain asymbolia
C0002768|Asymbolia
C0027743|Compression Syndrome, Nerve
C0027743|Compression Syndromes, Nerve
C0027743|Nerve Compression Syndrome
C0027743|Nerve Compression Syndromes
C0027743|Syndrome, Nerve Compression
C0027743|Syndromes, Nerve Compression
C0027743|Nerve Compression Syndromes [Disease/Finding]
C0027831|Neurofibromatosis 1
C0027831|von Recklinghausens Disease
C0027831|Recklinghausen's disease
C0027831|neurofibromatosis type 1 (NF1)
C0027831|NF1
C0027831|NEUROFIBROMATOSIS, TYPE I
C0027831|RECKLINGHAUSENS DIS OF NERVE
C0027831|NEUROFIBROMATOSIS A 01
C0027831|RECKLINGHAUSEN DIS OF NERVE
C0027831|VON RECKLINGHAUSENS DIS
C0027831|VON RECKLINGHAUSEN DIS
C0027831|von Recklinghausen's disease
C0027831|Recklinghausen's neurofibromatosis
C0027831|type I neurofibromatosis (diagnosis)
C0027831|neurofibromatosis type I (von Recklinghausen's disease)
C0027831|type I neurofibromatosis
C0027831|Type 1 Neurofibromatosis
C0027831|Type 1, Neurofibromatosis
C0027831|I, Neurofibromatosis Type
C0027831|Neurofibromatoses, Type I
C0027831|Type I Neurofibromatoses
C0027831|Type I, Neurofibromatosis
C0027831|Neurofibromatoses, Peripheral
C0027831|Neurofibromatosis, Peripheral
C0027831|Peripheral Neurofibromatoses
C0027831|Neurofibromatosis type I
C0027831|Recklinghausen Disease of Nerve
C0027831|Neurofibromatosis, Peripheral, NF 1
C0027831|NF1 (Neurofibromatosis 1)
C0027831|Neurofibromatosis, Peripheral, NF1
C0027831|Recklinghausen's Disease of Nerve
C0027831|Recklinghausens Disease of Nerve
C0027831|Neurofibromatosis 1 [Disease/Finding]
C0027831|Peripheral Neurofibromatosis
C0027831|Neurofibromatosis Type 1
C0027831|Neurofibromatosis, Type 1
C0027831|Recklinghausen Disease, Nerve
C0027831|von Recklinghausen Disease
C0027831|Neurofibromatosis I
C0027831|Neurofibromatosis, type 1 [von recklinghausen's disease]
C0027831|Neurofibromatosis, Peripheral Type
C0027831|Molluscum Fibrosum
C0027831|Clinical von Reclinghausen's disease
C0027831|Neurofibromatosis (nonmalignant) type
C0027831|[M]Von Recklinghausen's disease
C0027831|Neurofibromatosis 1 (disorder)
C0027831|Neurofibromatosis, type 1 (von Recklinghausen's disease)
C0027831|Von Recklinghausen's disease (of nerve)
C0027831|Neurofibromatosis, type 1 (disorder)
C0027831|disease; Von Recklinghausen
C0027831|Von Recklinghausen; disease
C0031118|Neoplasm, Peripheral Nerve
C0031118|Neoplasms, Peripheral Nerve
C0031118|Nerve Neoplasm, Peripheral
C0031118|Nerve Neoplasms, Peripheral
C0031118|Peripheral Nerve Neoplasm
C0031118|PERIPHERAL NERVE NEOPL
C0031118|PNS NEOPL
C0031118|neoplasm of peripheral nervous system
C0031118|neoplasm of peripheral nervous system (diagnosis)
C0031118|neoplasm of PNS
C0031118|Peripheral Nervous System Neoplasms
C0031118|Peripheral Nerve Neoplasms
C0031118|Peripheral Nerve Tumors
C0031118|Peripheral Nervous System Neoplasms [Disease/Finding]
C0031118|Nerves, Peripheral--Tumors
C0031118|CNS-excluded nervous sys. cancer
C0031118|CNS-excluded nervous system cancer, NOS
C0031118|Tumor of the peripheral nervous system
C0031118|Neoplasm of the peripheral nervous system
C0031118|Peripheral nervous system neoplasm NOS
C0031118|Peripheral nervous system neoplasm
C0031118|Tumor of peripheral nerve
C0031118|Tumour of peripheral nerve
C0031118|Neoplasm of peripheral nerve (disorder)
C0031118|Neoplasm of peripheral nerve
C0031118|Peripheral Nerve Tumor
C0031118|Neoplasm of the PNS
C0031118|Neoplasm of the Peripheral Nerve
C0031118|Neoplasms, PNS
C0031118|Neoplasms, Peripheral Nervous System
C0031118|PNS Neoplasms
C0031118|PNS Neoplasm
C0031118|PNS Tumor
C0031118|Peripheral Nervous System Tumor
C0031118|Tumor of PNS
C0031118|Tumor of Peripheral Nervous System
C0031118|Tumor of the PNS
C0031118|Tumor of the Peripheral Nerve
C0031118|Nerve Tumor, Peripheral
C0031118|Nerve Tumors, Peripheral
C0031118|Tumor, Peripheral Nerve
C0031118|Tumors, Peripheral Nerve
C0152025|Polyneuropathy
C0152025|Polyneuropathy, unspecified
C0152025|polyneuropathy (diagnosis)
C0152025|Polyneuropathies
C0152025|Polyneuropathies [Disease/Finding]
C0152025|Polyneuropathy (multiple nerve disorder)
C0152025|Polyneuropathy unspecified
C0152025|Polyneuropathy (disorder)
C0152025|[X]Polyneuropathy, unspecified (disorder)
C0152025|Polyneuropathy unspecified (disorder)
C0152025|[X]Polyneuropathy, unspecified
C0152025|Polyneuropathy NOS
C0152025|neuropathy; multiple
C0152025|Polyneuropathy, NOS
C0700594|Radiculopathy
C0700594|radiculopathy (diagnosis)
C0700594|Radiculopathies
C0700594|Radiculopathy, site unspecified
C0700594|Radiculopathy [Disease/Finding]
C0700594|Radicular syndrome
C0700594|Radiculopathy (disorder)
C0700594|Radiculopathy NOS
C0700594|Spinal nerve root disorder NOS
C0700594|neuropathy; radicular
C0700594|radicular; neuropathic
C0700594|radicular; syndrome
C0700594|syndrome; radicular
C0700594|Radiculopathy, NOS
C0206247|Amyloid Neuropathies
C0206247|Amyloid Polyneuropathy
C0206247|Neuropathy, Amyloid
C0206247|Polyneuropathies, Amyloid
C0206247|Amyloid Neuropathy
C0206247|Polyneuropathy, Amyloid
C0206247|amyloid polyneuropathy (diagnosis)
C0206247|Amyloid Polyneuropathies
C0206247|Neuropathies, Amyloid
C0206247|Amyloid Neuropathies [Disease/Finding]
C0206247|Amyloid polyneuropathy (disorder)
C0206247|Polyneuropathy in amyloidosis
C0206247|Polyneuropathy in amyloidosis (disorder)
C3542501|Guillain-Barre Syndrome
C3542501|Syndrome, Guillain-Barre
C3542501|Guillain Barre Syndrome
C3542501|acute idiopathic polyneuritis
C3542501|AIDP
C3542501|ACUTE INFLAMM POLYRADICULONEUROPATHY
C3542501|DEMYELINATING POLYRADICULONEUROPATHY ACUTE INFLAMM
C3542501|INFLAMM POLYNEUROPATHY ACUTE
C3542501|POLYNEUROPATHY ACUTE INFLAMM
C3542501|POLYRADICULONEUROPATHY ACUTE INFLAMM DEMYELINATING
C3542501|INFLAMM DEMYELINATING POLYRADICULONEUROPATHY ACUTE
C3542501|ACUTE INFLAMM POLYNEUROPATHY
C3542501|POLYRADICULONEUROPATHY ACUTE INFLAMM
C3542501|ACUTE INFLAMM DEMYELINATING POLYRADICULONEUROPATHY
C3542501|acute postinfectious polyneuropathy
C3542501|Landry's paralysis
C3542501|postinfectious polyneuritis
C3542501|Infectious neuronitis
C3542501|acute infectious polyneuritis (diagnosis)
C3542501|acute infectious polyneuritis
C3542501|Acute Autoimmune Neuropathies
C3542501|Autoimmune Neuropathies, Acute
C3542501|Autoimmune Neuropathy, Acute
C3542501|Neuropathies, Acute Autoimmune
C3542501|Neuropathy, Acute Autoimmune
C3542501|Acute Inflammatory Polyneuropathies
C3542501|Inflammatory Polyneuropathies, Acute
C3542501|Polyneuropathies, Acute Inflammatory
C3542501|Inflammatory Polyneuropathy, Acute
C3542501|Acute Inflammatory Polyradiculoneuropathies
C3542501|Inflammatory Polyradiculoneuropathies, Acute
C3542501|Polyradiculoneuropathies, Acute Inflammatory
C3542501|Landry Guillain Barre Syndrome
C3542501|Syndrome, Landry-Guillain-Barre
C3542501|Guillaine Barre Syndrome
C3542501|Syndrome, Guillaine-Barre
C3542501|Ac infect polyneuritis
C3542501|Acute, Inflammatory Polyneuropathy
C3542501|Polyneuropathy Acute, Inflammatory
C3542501|Inflammatory Polyneuropathy Acutes
C3542501|Inflammatory Demyelinating Polyradiculoneuropathy, Acute
C3542501|Acute Autoimmune Neuropathy
C3542501|Acute Inflammatory Polyneuropathy
C3542501|Demyelinating Polyradiculoneuropathy, Acute Inflammatory
C3542501|Polyneuropathy, Acute Inflammatory
C3542501|Polyradiculoneuropathy, Acute Inflammatory Demyelinating
C3542501|Inflammatory Polyneuropathy Acute
C3542501|Acute Inflammatory Demyelinating Polyradiculoneuropathy
C3542501|Acute Inflammatory Polyradiculoneuropathy
C3542501|Polyradiculoneuropathy, Acute Inflammatory
C3542501|Acute Inflammatory Demyelinating Polyneuropathy
C3542501|Infectious polyneuritis
C3542501|Acute infective polyneuritis (& [Guillain-Barre syndrome]) (disorder)
C3542501|Acute infective polyneuritis
C3542501|Acute inf. polyneuritis
C3542501|Acute inflammatory demyelinating polyneuropathy (disorder)
C3542501|Acute infective polyneuritis NOS
C3542501|Acute infective polyneuritis NOS (disorder)
C3542501|Acute infective polyneuritis (& [Guillain-Barre syndrome])
C3542501|Acute infective polyneuritis (disorder)
C3542501|Ascending paralysis (finding)
C3542501|Ascending paralysis
C3542501|Polyneuropathy, Inflammatory Demyelinating, Acute
C3542501|Acute Inflammatory Demyelinating Polyradiculopathy
C3542501|Paralysis ascending
C3542501|Guillaine-Barre Syndrome
C3542501|Landry-Guillain-Barre Syndrome
C3542501|Guillain-Barre Syndrome, Familial
C3542501|Acute inflammatory neuropathy
C3542501|Acute post-infective radiculoneuropathy
C3542501|Post-infectious polyneuritis
C3542501|Acute idiopathic polyradiculoneuritis
C3542501|Infectious neuronitis (disorder)
C3542501|Post-infectious polyneuritis (disorder)
C3542501|ascending; paralysis
C3542501|Landry; paralysis
C3542501|infective; polyneuritic
C3542501|multiple; neuritis, infective, acute
C3542501|neuritis; multiple, infective, acute
C3542501|paralysis; Landry
C3542501|paralysis; ascending
C3542501|polyneuritis; acute
C3542501|polyneuritis; infective
C3542501|polyneuritis; postinfective
C3542501|postinfective; polyneuritic
C3542501|PNS neuronitis
C0242287|Isaac Syndrome
C0242287|Isaacs Mertens Syndrome
C0242287|Isaacs Syndrome
C0242287|ISAACS-MERTENS SYNDROME
C0242287|Isaacs syndrome (diagnosis)
C0242287|Continuous Myokymia
C0242287|Continuous Myokymias
C0242287|Myokymias, Continuous
C0242287|Gamstorp Wohlfart Syndrome
C0242287|Isaacs Pseudomyotonia Syndrome
C0242287|Pseudomyotonia
C0242287|Isaacs Syndrome [Disease/Finding]
C0242287|Gamstorp-Wohlfart Syndrome
C0242287|Isaacs' Syndrome
C0242287|Myokymia, Continuous
C0242287|Neuromyotonia
C0242287|Pseudomyotonia Syndrome of Isaacs
C0242287|Continuous Muscle Activity Syndrome
C0242287|Syndrome of Continuous Muscle Activity
C0242287|Quantal Squander
C0242287|Syndromes, Gamstorp-Wohlfart
C0242287|Syndromes, Isaacs-Mertens
C0242287|Gamstorp-Wohlfart Syndromes
C0242287|Myokymia, Myotonia, Muscle Wasting, And Hyperhidrosis
C0242287|NMAN
C0242287|NEUROMYOTONIA AND AXONAL NEUROPATHY, AUTOSOMAL RECESSIVE
C0242287|Neuromyotonia (disorder)
C0242287|Gamstorp disease
C0242287|MYOKYMIA, MYOTONIA, AND MUSCLE WASTING
C0242287|Autosomal recessive neuromyotonia with axonal neuropathy
C0242287|Autosomal recessive axonal neuropathy with neuromyotonia (disorder)
C0242287|Myokymia, myotonia and muscle wasting
C0242287|Autosomal recessive axonal neuropathy with neuromyotonia
C0242287|Isaac's syndrome
C0242287|Continuous muscle fiber activity
C0242287|Continuous muscle fibre activity
C0242287|Isaacs syndrome (disorder)
C0242287|Isaacs
C0242287|Neuromyotonia [Ambiguous]
C0494491|Mononeuropathy, unspecified
C0494491|Mononeuropathy
C0494491|Mononeuropathies
C0494491|Mononeuropathies [Disease/Finding]
C0494491|Mononeuropathy (disorder)
C0494491|Mononeuropathy NOS
C0700251|Brachial Plexus Neuropathies
C0700251|Brachial plexus disorders
C0700251|BRACHIAL PLEXUS DIS
C0700251|Brachial Plexus Disease
C0700251|Plexus Disease, Brachial
C0700251|Plexus Diseases, Brachial
C0700251|Brachial Plexus Disorder
C0700251|Plexus Disorder, Brachial
C0700251|Plexus Disorders, Brachial
C0700251|Brachial Plexus Neuropathy
C0700251|Neuropathies, Brachial Plexus
C0700251|Neuropathy, Brachial Plexus
C0700251|Plexus Neuropathies, Brachial
C0700251|Plexus Neuropathy, Brachial
C0700251|Plexopathies, Brachial
C0700251|Plexopathy, Brachial
C0700251|Brachial Plexopathy
C0700251|Brachial Plexus Diseases
C0700251|Brachial Plexus Neuropathies [Disease/Finding]
C0700251|brachial plexus disorder (diagnosis)
C0700251|Brachial plexus--Diseases
C0700251|BPN - Brachial plexus neuropathy
C0700251|Brachial plexus disorder (disorder)
C0700251|brachial plexus; neuropathy
C0700251|brachial plexus; syndrome
C0700251|disease (or disorder); plexus, brachial
C0700251|neuropathy; brachial plexus
C0700251|plexus brachialis; neuropathic
C0700251|syndrome; brachial plexus
C0700251|Brachial plexus neuropathy, NOS
C0458219|Complex regional pain syndrome NOS
C0458219|Complex Regional Pain Syndromes
C0458219|Complex Regional Pain Syndromes [Disease/Finding]
C0458219|CRPS (Complex Regional Pain Syndromes)
C0458219|Pain Syndromes, Regional Complex
C0458219|CRPS
C0458219|Complex Regional Pain Syndrome
C0458219|Complex regional pain syndrome (CRPS)
C0458219|Complex regional pain syndrome (diagnosis)
C0458219|Complex regional pain syndrome (disorder)
C0458219|Complex regional pain syndromes (disorder)
C1363854|Hand Arm Vibration Syndrome
C1363854|Hand-Arm Vibration Syndromes
C1363854|Hand-Arm Vibration Syndrome
C1363854|Syndrome, Hand-Arm Vibration
C1363854|Syndromes, Hand-Arm Vibration
C1363854|Vibration Syndrome, Hand-Arm
C1363854|Vibration Syndromes, Hand-Arm
C1363854|Hand-Arm Vibration Syndrome [Disease/Finding]
C1363854|Hand and arm vibration syndrome
C0031117|Nerve Disease, Peripheral
C0031117|Nerve Diseases, Peripheral
C0031117|Peripheral Nerve Disease
C0031117|Peripheral Nerve Diseases
C0031117|Disorders of the peripheral nervous system
C0031117|Peripheral Nervous System Diseases
C0031117|PNS Disease
C0031117|peripheral neuropathy
C0031117|PNS DIS
C0031117|PERIPHERAL NERVOUS SYSTEM DIS
C0031117|PERIPHERAL NERVE DIS
C0031117|PNS PERIPHERAL NERVOUS SYSTEM DIS
C0031117|peripheral nervous system disorder
C0031117|peripheral neuropathy (diagnosis)
C0031117|peripheral neuropathy (physical finding)
C0031117|Peripheral neuropathies
C0031117|Neuropathy, Peripheral
C0031117|Disorder of peripheral nervous system NOS
C0031117|PNS Diseases
C0031117|Peripheral Nervous System Disease
C0031117|Peripheral Nervous System Diseases [Disease/Finding]
C0031117|PNS (Peripheral Nervous System) Diseases
C0031117|Peripheral Nervous System Disorders
C0031117|Peripheral nerve disorder
C0031117|PN - Peripheral neuropathy
C0031117|Neuropathy;peripheral
C0031117|Peripheral Nerve Disorders
C0031117|disorders of peripheral nervous system
C0031117|disorders of peripheral nervous system (diagnosis)
C0031117|Peripheral nervous system disorders (disorder)
C0031117|Peripheral nervous system disorder NOS
C0031117|Peripheral nervous system disorder NOS (disorder)
C0031117|Nerves, Peripheral--Diseases
C0031117|Disorder of Peripheral Nervous System
C0031117|Neuropathy peripheral
C0031117|Peripheral neuropathy NOS
C0031117|Peripheral nerve disorder NOS
C0031117|Disorder of the peripheral nervous system (disorder)
C0031117|Disorder of the peripheral nervous system
C0031117|Peripheral nerve disease (disorder)
C0031117|neuropathy; peripheral
C0031117|peripheral; nervous system, disorder
C0031117|peripheral; neuropathic
C0031117|Disorder of the peripheral nervous system, NOS
C0031117|Peripheral nerve disorder, NOS
C0031117|Peripheral neuropathy, NOS
C0520720|Perineurial cyst
C0520720|Cyst, Perineural
C0520720|Cysts, Perineural
C0520720|Perineural Cyst
C0520720|Cysts, Tarlov
C0520720|Tarlov Cysts
C0520720|Cyst, Perineurial
C0520720|Cysts, Perineurial
C0520720|Tarlov Cyst
C0520720|Tarlov Cysts [Disease/Finding]
C0520720|Perineural Cysts
C0520720|Perineurial Cysts
C0520720|Cysts, Sacral Tarlov
C0520720|Cysts, Sacral Perineural
C0520720|Cyst, Sacral Perineural
C0520720|Sacral Perineural Cyst
C0520720|Sacral Perineural Cysts
C0520720|Sacral Tarlov Cysts
C0520720|tarlov cyst (diagnosis)
C0520720|Tarlov's cyst
C0520720|Nerve root cyst
C0520720|Perineurial cyst (disorder)
C0520720|Cyst of Nerve Root
C0520720|Cyst of the Nerve Root
C0852421|Acute polyneuropathy
C0852421|Acute polyneuropathies
C0598589|hereditary neuropathy
C0598589|Inherited neuropathies
C0598589|neuropathy; hereditary
C0598589|Inherited Neuropathy
C0853004|Peripheral neuropathies NEC
C1167650|Polyneuropathy chronic
C1167650|Chronic polyneuropathies
C1167650|Chronic Polyneuropathy
C0750944|PERIPHERAL AUTONOMIC NERVOUS SYSTEM DIS
C0750944|AUTONOMIC PERIPHERAL NERVOUS SYSTEM DIS
C0750944|Autonomic Peripheral Nervous System Diseases
C0750944|Disorder of peripheral autonomic nervous system (disorder)
C0750944|Disorder of peripheral autonomic nervous system
C0750944|disease (or disorder); peripheral, autonomic nervous system
C0750944|Disorder of peripheral autonomic nervous system, NOS
C0750944|Peripheral Autonomic Nervous System Diseases
C0393912|Autonomic Dysfunction, Segmental
C0393912|Autonomic Dysfunctions, Segmental
C0393912|Segmental Autonomic Dysfunctions
C0393912|Segmental Autonomic Dysfunction
C0393912|Segmental autonomic dysfunction (disorder)
C0393918|Drug-induced autonomic dysfunction
C0393918|Drug-induced autonomic dysfunction (disorder)
C0393920|Chronic idiopathic anhidrosis
C0393920|Chronic idiopathic anhidrosis (disorder)
C0393921|Idiopathic diffuse hyperhidrosis
C0393921|Idiopathic diffuse hyperhidrosis (disorder)
C0259749|autonomic neuropathy
C0259749|Autonomic neuropathy NOS
C0259749|Autonomic neuropathy (disorder)
C0560614|Autonomic nerve injury
C0560614|Autonomic nerve injury (disorder)
C1269759|Immature autonomic stability
C1269759|Immature autonomic system (disorder)
C1269759|Immature autonomic system
C0542142|Recurrent Laryngeal Nerve Paralysis
C0542142|Recurrent Laryngeal Nerve Palsy
C0542142|Vagus Nerve Laryngeal Paralysis
C0542142|Paralysis recurrent laryngeal nerve
C0542142|Vagus nerve laryngeal paralysis (disorder)
C0542142|Laryngeal Nerve Palsy, Recurrent
C2317111|Peripheral nerve disorder associated with repair of hernia
C2317111|Peripheral nerve disorder associated with repair of hernia (disorder)
C0393911|Bradbury Eggleston Syndrome
C0393911|Syndrome, Bradbury-Eggleston
C0393911|Pure Autonomic Failure
C0393911|AUTONOMIC FAILURE, PURE
C0393911|Bradbury-Eggleston Syndrome
C0393911|Pure Autonomic Failure [Disease/Finding]
C0393911|Autonomic failure
C0393911|Pure autonomic failure (disorder)
C1850386|GAN1
C1850386|GIANT AXONAL NEUROPATHY 1
C1850386|Axonal Neuropathy, Giant (GAN)
C1850386|Axonal Neuropathy, Giant
C1850386|Neuropathy, Giant Axonal (GAN)
C1850386|Giant Axonal Neuropathy
C1850386|Giant Axonal Neuropathy [Disease/Finding]
C1850386|Giant Axonal Neuropathy 1 (GAN1)
C1850386|Neuropathy, Giant Axonal
C1850386|Giant Axonal Neuropathy (GAN)
C1850386|Neuropathy, Giant Axonal, Autosomal Recessive
C1850386|GIANT AXONAL NEUROPATHY 1, AUTOSOMAL RECESSIVE
C1850386|GAN
C1850386|Giant axonal neuropathy (disorder)
C1263833|Phrenic neuropathy
C1263833|Phrenic nerve disorder (disorder)
C1263833|Phrenic nerve disorder
C1263833|n.phrenicus; disorder
C0338551|Leprosy neuropathy
C0338551|Leprosy neuropathy (disorder)
C0542368|amyloidosis with peripheral autonomic neuropathy
C0542368|amyloidosis with peripheral autonomic neuropathy (diagnosis)
C0542368|Autonomic neuropathy due to amyloid
C0542368|Autonomic neuropathy due to amyloid (disorder)
C0154741|Mononeuritis of upper limb and mononeuritis multiplex
C0154741|Mononeuritis of upper limb and mononeuritis multiplex (disorder)
C0553762|Anterior interosseous nerve syndrome
C0553762|Anterior interosseous nerve lesion
C0553762|Anterior interosseous nerve lesion (disorder)
C0553763|Posterior interosseous nerve lesion
C0553763|Posterior interosseous nerve lesion (disorder)
C0423675|Thoracic and lumbosacral neuritis NOS (disorder)
C0423675|Thoracic and lumbosacral neuritis NOS
C0423675|Thoracic and lumbosacral neuritis
C0423675|Thoracic and lumbosacral neuritis (disorder)
C0273529|Injury to peripheral nerve(s) of shoulder girdle and upper limb
C0273529|Injury to unspecified nerve of shoulder girdle and upper limb
C0273529|Injury of nerves at shoulder and upper arm level
C0273529|Injury of unspecified nerve at shoulder and upper arm level
C0273529|Injury of peripheral nerve of shoulder girdle AND/OR upper limb-RETIRED
C0273529|injury of peripheral nerve of shoulder girdle and upper limb
C0273529|injury of peripheral nerve of shoulder girdle and upper limb (diagnosis)
C0273529|Injury to unspecified peripheral nerve of shoulder girdle and upper limb
C0273529|Inj nerve shldr/arm NOS
C0273529|peripheral nerve injury at shoulder and upper arm level (diagnosis)
C0273529|peripheral nerve injury at shoulder and upper arm level
C0273529|peripheral nerve injury shoulder and upper arm level
C0273529|Shoulder girdle peripheral nerve injury
C0273529|Shoulder girdle or upper limb peripheral nerve injury NOS
C0273529|Injury of peripheral nerve of shoulder girdle AND/OR upper limb (disorder)
C0273529|Injury of peripheral nerve of shoulder girdle AND/OR upper limb
C0273529|Arm peripheral nerve injury
C0273529|[X]Injury of unspecified nerve at shoulder and upper arm level
C0273529|Peripheral nerve injury: [shoulder girdle] &/or [upper limb] or [arm]
C0273529|Shoulder girdle and upper limb peripheral nerve injury
C0273529|[X]Injury of unspecified nerve at shoulder and upper arm level (disorder)
C0273529|Shoulder girdle or upper limb peripheral nerve injury NOS (disorder)
C0273529|Peripheral nerve injury: [shoulder girdle] &/or [upper limb] or [arm] (disorder)
C0273529|Injury of nerves at shoulder and upper arm level (disorder)
C0273529|Injury of peripheral nerve of shoulder girdle and upper limb, NOS
C0273529|Injury to peripheral nerve of shoulder girdle and upper limb
C0273529|Injury to peripheral nerves of shoulder girdle and upper limb
C0393802|Hereditary or idiopathic peripheral neuropathy NOS
C0393802|Peripheral neuropathy - hereditary or idiopathic
C0393802|Hereditary or idiopathic peripheral neuropathy NOS (disorder)
C0393802|Peripheral neuropathy - hereditary or idiopathic (disorder)
C2239188|BURNING, FEET SYNDROME
C2239188|Burning feet syndrome
C2239188|Burning feet syndrome (disorder)
C2239188|Strachan's syndrome
C2239188|burning feet; syndrome
C2239188|burning; feet syndrome
C2239188|foot; burning (syndrome)
C2239188|foot; syndrome, burning
C2239188|syndrome; burning feet
C0338553|Intercostal post-herpetic neuralgia
C0338553|Intercostal post-herpetic neuralgia (disorder)
C0472363|Ischaemic neuropathy due to arterial steal
C0472363|Ischemic neuropathy due to arterial steal
C0472363|Ischemic neuropathy due to arterial steal (disorder)
C0553760|Lumbosacral plexus neuropathy
C0553760|Lumbosacral plexus neuropathy (disorder)
C0393880|Peripheral nerve compression arm
C0393880|Compression neuropathy of upper limb
C0393880|Compression neuropathy of upper limb (disorder)
C0393896|Compression neuropathy of trunk
C0393896|Compression neuropathy of trunk (disorder)
C0393897|Intercostal neuropathy
C0393897|intercostal neuropathy (diagnosis)
C0393897|Intercostal neuropathy (disorder)
C0393897|disease (or disorder); intercostal nerve
C0393919|PARANEOPL AUTONOMIC DYSFUNCTION
C0393919|AUTONOMIC DYSFUNCTION PARANEOPL
C0393919|Autonomic Dysfunctions, Paraneoplastic
C0393919|Paraneoplastic Autonomic Dysfunctions
C0393919|Autonomic Dysfunction, Paraneoplastic
C0393919|Paraneoplastic autonomic dysfunction
C0393919|Paraneoplastic autonomic dysfunction (disorder)
C0270922|Demyelinating peripheral neuropathy
C0270922|Demyelinating neuropathy
C0270922|Peripheral demyelinating neuropathy
C0270922|Demyelinating polyneuropathy
C0270922|Demyelinating polyneuropathy NOS
C0270922|Peripheral demyelinating neuropathy (disorder)
C0270922|Demyelinating neuropathy, NOS
C0270922|Demyelinating polyneuropathy, NOS
C0266517|Congenital peripheral nerve disorders
C0266517|Congenital anomaly of peripheral nerve (disorder)
C0266517|Congenital anomaly of peripheral nerve
C0266517|Congenital anomaly of nerve, NOS
C0413275|Peripheral nerve decompression injury
C0413275|Peripheral nerve decompression injury (disorder)
C0423709|Cruralgia
C0423709|Cruralgia (disorder)
C0344306|Intercostal neuralgia
C0344306|Intercostal neuralgia (disorder)
C0394021|Disorder of peripheral nerve graft
C0394021|Disorder of peripheral nerve graft (disorder)
C0565585|Neuralgia/neuritis - shoulder (disorder)
C0565585|Neuralgia/neuritis - shoulder
C0565586|Neuralgia/neuritis - upper arm (disorder)
C0565586|Neuralgia/neuritis - upper arm
C0565590|Neuralgia/neuritis - lower leg
C0565590|Neuralgia/neuritis - lower leg (disorder)
C0565591|Neuralgia/neuritis -ankle/foot
C0565591|Neuralgia/neuritis - ankle/foot
C0565591|Neuralgia/neuritis - ankle/foot (disorder)
C0574717|Upper limb nerve lesion
C0574717|Upper limb nerve lesion (disorder)
C0574718|Lower limb nerve lesion
C0574718|Lower limb nerve lesion (disorder)
C0574920|Thoracoabdominal neuropathy
C0574920|Thoracoabdominal neuropathy (disorder)
C0153097|polyneuropathy due to mumps
C0153097|polyneuropathy due to mumps (diagnosis)
C0153097|Polyneuropathy mumps
C0153097|Mumps polyneuropathy
C0153097|Polyneuropathy in mumps (disorder)
C0153097|Polyneuropathy in mumps
C0153097|Mumps polyneuropathy (disorder)
C0271686|Diabetic autonomic neuropathy
C0271686|diabetes mellitus with autonomic neuropathy (diagnosis)
C0271686|diabetes mellitus with autonomic neuropathy
C0271686|Autonomic Neuropathies, Diabetic
C0271686|Autonomic Neuropathy, Diabetic
C0271686|Diabetic Autonomic Neuropathies
C0271686|Neuropathies, Diabetic Autonomic
C0271686|Neuropathy, Diabetic Autonomic
C0271686|Autonomic neuropathy due to diabetes
C0271686|Diabetic autonomic neuropathy (disorder)
C0037887|Sphenopalatine neuralgia
C0037887|Neuralgia, Sphenopalatine
C0037887|Neuralgias, Sphenopalatine
C0037887|Sphenopalatine Neuralgias
C0037887|Sluder's neuralgia
C0037887|Sphenopalatine ganglion neuralgia
C0037887|Sluder's syndrome
C0037887|Sphenopalatine neuralgia (disorder)
C0037887|Sluder
C0037887|neuralgia; sphenopalatine
C0037887|sphenopalatine; neuralgia
C1527351|NERVE ROOT DIS
C1527351|Nerve Root Disorders
C1527351|Nerve root disorder
C1527351|Nerve root disorder (disorder)
C1527351|Nerve root disorder, NOS
C0262593|Peripheral nerve injury
C0262593|injury of peripheral nerve (diagnosis)
C0262593|injury of peripheral nerve
C0262593|Injury;nerve;peripheral
C0262593|Nerve Injuries, Peripheral
C0262593|Nerve Injury, Peripheral
C0262593|Injury, Peripheral Nerve
C0262593|Injuries, Peripheral Nerve
C0262593|Peripheral Nerve Injuries
C0262593|Peripheral Nerve Injuries [Disease/Finding]
C0262593|Peripheral nerve injury NOS
C0262593|Peripheral nerve injury NOS (disorder)
C0262593|Peripheral nerve injury (disorder)
C0262593|PNI - Peripheral nerve injury
C0262593|injury; nerve, peripheral
C0262593|nerve; injury, peripheral
C0262593|Peripheral nerve injury, NOS
C0338536|neuralgia superior laryngeal
C0338536|superior laryngeal neuralgia (diagnosis)
C0338536|superior laryngeal neuralgia
C0338536|Superior laryngeal neuralgia (disorder)
C0270910|idiopathic peripheral neuropathy
C0270910|idiopathic peripheral neuropathy (diagnosis)
C0270910|Idiopathic peripheral neuropathy (disorder)
C0270910|neuropathy; peripheral, idiopathic
C0270910|Idiopathic peripheral neuropathy, NOS
C1868426|PERONEAL NERVE, ACCESSORY DEEP
C1868426|Accessory deep peroneal nerve
C0795950|ACCPN
C0795950|AGENESIS OF THE CORPUS CALLOSUM WITH PERIPHERAL NEUROPATHY
C0795950|Corpus callosum agenesis neuronopathy
C0795950|Andermann syndrome
C0795950|Charlevoix disease
C0795950|Polyneuropathy, sensorimotor, with or without agenesis of the corpus callosum
C0795950|Corpus Callosum, Agenesis of, with Neuronopathy
C0795950|Agenesis of Corpus Callosum with Peripheral Neuropathy
C0795950|Agenesis of Corpus Callosum with Polyneuropathy
C0795950|Agenesis of Corpus Callosum with Neuronopathy
C0795950|Hereditary Motor and Sensory Neuropathy with Agenesis of the Corpus Callosum
C0795950|Agenesis of corpus callosum with peripheral neuropathy (disorder)
C0796123|CATARACT-ATAXIA-DEAFNESS-RETARDATION SYNDROME
C0796123|Cataract ataxia deafness
C0796123|Begeer syndrome
C0796123|Cataract ataxia deafness syndrome
C0796123|Polyneuropathy, cataract, deafness syndrome
C0796123|Polyneuropathy-Cataract-Deafness Syndrome
C1850406|NN
C1850406|NAVAJO NEUROHEPATOPATHY
C1850406|Navajo neuropathy
C1850406|NNH
C1850406|MITOCHONDRIAL DNA DEPLETION SYNDROME 6 (HEPATOCEREBRAL TYPE)
C1850406|MTDPS6
C1850406|MPV17-Associated Hepatocerebral MDS
C1850406|MPV17-Related Hepatocerebral Mitochondrial DNA Depletion Syndrome
C1850406|Mitochondrial Dna Depletion Syndrome 6
C2932678|Inherited Peripheral Neuropathy
C0006091|Brachial plexus lesions
C0006091|Lesion;brachial plexus
C0006091|Brachial plexus lesions NOS
C0006091|Brachial plexus lesions NOS (disorder)
C0006091|Brachial plexus lesion
C0006091|brachial plexus; lesion
C0006091|lesion; brachial plexus
C0006091|plexus brachialis; lesion
C0006091|Brachial plexus lesion, NOS
C0006091|lesion of brachial plexus
C2959948|Ependymal cyst of spinal nerve (disorder)
C2959948|Ependymal cyst of spinal nerve
C0271676|Abdominal Polyradiculopathies
C0271676|Abdominal Polyradiculopathy
C0271676|Polyradiculopathies, Abdominal
C0271676|Abdominal polyradiculopathy (disorder)
C0271676|Polyradiculopathy, Abdominal
C2119284|uncontrolled type I diabetes mellitus with peripheral neuropathy (diagnosis)
C2119284|type 1 diabetic peripheral neuropathy, uncontrolled
C2119284|uncontrolled type 1 diabetes mellitus with peripheral neuropathy (diagnosis)
C2119284|uncontrolled type 1 diabetes mellitus with peripheral neuropathy
C1827029|Entrapment neuropathy of upper limb (disorder)
C1827029|Entrapment neuropathy of upper limb
C0154758|Inflammatory and toxic neuropathy
C0154758|Unspecified inflammatory and toxic neuropathies
C0154758|Inflam/tox neuropthy NOS
C0154758|Unspecified inflammatory and toxic neuropathy
C0154758|Inflammatory &/or toxic neuropathy (disorder)
C0154758|Toxic or inflammatory neuropathy NOS
C0154758|Toxic or inflammatory neuropathy NOS (disorder)
C0154758|Inflammatory &/or toxic neuropathy
C0154758|Inflammatory and toxic neuropathy (disorder)
C0270109|Phrenic nerve paralysis due to birth injury
C0270109|Phrenic nerve paralysis as birth trauma
C0270109|Phrenic nerve paralysis as birth trauma (disorder)
C0270109|Phrenic nerve paralysis due to birth trauma
C0393852|Neuropathy due to infection
C0393852|Neuropathy due to infection (disorder)
C0273522|Cauda equina injury without bony injury (disorder)
C0273522|Cauda equina injury without bony injury
C0273522|Cauda equina injury without bone injury
C0273522|Cauda equina injury without bone injury (disorder)
C0393841|Neuropathy in liver disease
C0393841|Neuropathy in liver disease (disorder)
C0393841|Hepatic neuropathy (disorder)
C0393841|Hepatic neuropathy
C0160799|Late effect of injury to peripheral nerve of shoulder girdle and upper limb
C0160799|Sequelae of injury of nerve of upper limb
C0160799|late effects of injury of peripheral nerve of shoulder girdle and upper limb (diagnosis)
C0160799|late effects of injury of peripheral nerve of shoulder girdle and upper limb
C0160799|Late effect of injury of peripheral nerve of shoulder girdle and upper limb
C0160799|Lt eff nerv inj shld/arm
C0160799|Late effect of injury to peripheral nerve of shoulder girdle AND/OR upper limb (disorder)
C0160799|Late effect of injury to peripheral nerve of shoulder girdle AND/OR upper limb
C0270102|Birth injury to peripheral nervous system
C0270102|Birth injury to peripheral nervous system, unspecified
C0270102|peripheral nerve injury due to birth trauma (diagnosis)
C0270102|peripheral nerve injuries due to birth trauma
C0270102|peripheral nerve injury due to birth trauma
C0270102|Peripheral nerve injury as birth trauma
C0270102|Peripheral nerve injury as birth trauma (disorder)
C0270102|Peripheral nerve injury due to birth trauma (disorder)
C0270102|birth; injury, laceration, peripheral nerve
C0270102|birth; injury, nerve, peripheral
C0270102|injury; birth, laceration, peripheral nerve
C0270102|injury; birth, nerve, peripheral
C0347066|malignant infiltration of peripheral nerve
C0347066|neoplasm - pns malignant infiltration
C0347066|malignant infiltration of peripheral nerve (diagnosis)
C0347066|Malignant infiltration of peripheral nerve (disorder)
C0270933|Inflammatory neuropathy
C0270933|Inflammatory neuropathy (disorder)
C0270933|Inflammatory neuropathy, NOS
C0393410|Other specified disorders of peripheral nervous system (disorder)
C0393410|Other specified disorders of peripheral nervous system
C0560607|Intercostal post-herpetic neuritis
C0560607|Intercostal post-herpetic neuritis (disorder)
C0582681|Lesions of nerves plexuses and roots
C0582681|Lesions of nerves plexuses and roots (disorder)
C1510429|Neuropathies, Entrapment
C1510429|Neuropathy, Entrapment
C1510429|Nerve entrapment syndromes
C1510429|Compression neuropathy (disorder)
C1510429|Compression neuropathy
C1510429|Entrapment neuropathies
C1510429|Entrapment neuropathy
C1510429|Nerve entrapment syndrome
C1510429|Trapped nerve
C1510429|Peripheral nerve entrapment syndrome (disorder)
C1510429|Peripheral nerve entrapment syndrome
C1510429|neuropathy; entrapment
C1510429|Entrapment syndrome, NOS
C1510429|Entrapment neuropathy, NOS
C0271684|Diabetic pseudotabes
C0271684|Diabetic pseudotabes (disorder)
C0564741|Other peripheral nerve disease
C0564741|Other peripheral nerve disease (disorder)
C3647370|neuropathy peripheral in association with hereditary ataxia (diagnosis)
C3647370|neuropathy peripheral in association with hereditary ataxia
C3662005|Neuropathy of lower limb
C3662005|Neuropathy of lower limb (disorder)
C1282521|Pudendal nerve neuropathy (disorder)
C1282521|Pudendal nerve neuropathy
C3662002|Neuropathy of upper limb (disorder)
C3662002|Neuropathy of upper limb
C3661994|Disorder of nerve root and/or plexus (disorder)
C3661994|Disorder of nerve root and/or plexus
C0574905|Long thoracic nerve lesion
C0574905|Long thoracic nerve lesion (disorder)
C3670522|Dysmyelinogenesis (disorder)
C3670522|Dysmyelinogenesis
C2931445|Sacral plexopathy
C1845095|DFNX5
C1845095|AUNX1
C1845095|DEAFNESS, X-LINKED 5
C1845095|DEAFNESS, X-LINKED 5 (disorder)
C1845095|Auditory Neuropathy, X-Linked, 1, with Peripheral Sensory Neuropathy
C1833831|OPTIC ATROPHY, HEARING LOSS, AND PERIPHERAL NEUROPATHY, AUTOSOMAL DOMINANT
C1855885|HYPERTROPHIC NEUROPATHY AND CATARACT
C1850383|NEUROPATHY, PAINFUL
C1834180|NEUROPATHY, WITH PARAPROTEIN IN SERUM, CEREBROSPINAL FLUID AND URINE
C1850022|PERIPHERAL NEUROPATHY, ATAXIA, FOCAL NECROTIZING ENCEPHALOPATHY, AND SPONGY DEGENERATION OF BRAIN
C1866770|SPINOCEREBELLAR ATAXIA WITH RIGIDITY AND PERIPHERAL NEUROPATHY
C0031315|Limb, Phantom
C0031315|Limbs, Phantom
C0031315|Phantom Limb
C0031315|Phantom Limbs
C0031315|Phantom limb (syndrome)
C0031315|Phantom limb syndrome with pain
C0031315|phantom limb syndrome
C0031315|phantom limb syndrome (diagnosis)
C0031315|Pseudomelias
C0031315|Phantom limb syndrome NOS
C0031315|Phantom Limb [Disease/Finding]
C0031315|Pseudomelia
C0031315|phantom limb syndrome with pain (diagnosis)
C0031315|Phantom limb syndrome with pain (finding)
C0031315|Phantom limb (disorder)
C0031315|Phantom limb pain
C0031315|PLS - Phantom limb pain syndrome
C0031315|Stump hallucination
C0031315|Phantom pain
C0031315|PLS - Phantom limb syndrome
C0031315|Phantom limb syndrome (disorder)
C0031315|FLS - Phantom limb syndrome
C0031315|pain; phantom limb syndrome
C0031315|phantom limb syndrome; pain
C0031315|phantom limb; syndrome, with pain
C0031315|phantom limb; syndrome
C0031315|syndrome; phantom limb, with pain
C0031315|syndrome; phantom limb
C3873567|Peripheral neuropathy due to chemotherapy
C3873567|Chemotherapy-induced peripheral neuropathy
C3873567|Peripheral neuropathy due to chemotherapy (disorder)
C3873567|CIPN - Chemotherapy-induced peripheral neuropathy
C4024907|Mixed demyelinating and axonal polyneuropathy
C0271683|Motor polyneuropathy
C0271683|Motor Polyneuropathies
C0271683|Polyneuropathies, Motor
C0271683|Polyneuropathy, Motor
C0271683|Motor polyneuropathy (disorder)
C0020580|Hypesthesia
C0020580|Hypesthesias
C0020580|Hypoesthesias
C0020580|HYPOESTHESIA
C0020580|Hypoaesthesia
C0020580|Decreased Sensitivity
C0020580|[D]Hypoesthesia (context-dependent category)
C0020580|Sensory impairment
C0020580|Hypesthesias, Tactile
C0020580|Tactile Hypesthesia
C0020580|Tactile Hypesthesias
C0020580|Impaired Sensations
C0020580|Sensation, Impaired
C0020580|Sensations, Impaired
C0020580|Reduced Sensations
C0020580|Sensation, Reduced
C0020580|Sensations, Reduced
C0020580|Hypesthesia, Tactile
C0020580|Impaired Sensation
C0020580|Numbness
C0020580|Hypesthesia [Disease/Finding]
C0020580|Reduced Sensation
C0020580|Decreased;sensation
C0020580|Reduced sensation of skin (finding)
C0020580|Reduced sensation of skin
C0020580|[D]Hypesthesia
C0020580|Hypoaesthesia (reduced sensation)
C0020580|Hypoesthesia (reduced sensation)
C0020580|[D]Hypoesthesia
C0020580|Limited sensation
C0020580|[D]Hypoaesthesia
C0020580|[D]Hypoaesthesia (situation)
C0020580|[D]Hypoesthesia (situation)
C0020580|Cutaneous hypoesthesia
C0020580|Hypaesthesia
C0020580|Hypesthesia (finding)
C0020580|Tactile hypaesthesia
C0020580|Tactile hypesthesia (finding)
C0020580|decreased sensation
C1867971|Acute episodes of neuropathic symptoms
C1848695|Episodic peripheral neuropathy
C4024974|Sensorimotor polyneuropathy affecting arms more than legs
C1112256|Sensorimotor peripheral neuropathy
C1112256|Peripheral sensorimotor neuropathy
C1112256|Sensorimotor neuropathy
C1112256|Mixed polyneuropathy
C4024967|Congenital peripheral neuropathy
C4025794|Chronic sensorineural polyneuropathy
C1263857|Peripheral axonal neuropathy
C1263857|Axonal peripheral neuropathy
C1263857|Peripheral axonal neuropathy (disorder)
C1859178|Progressive polyneuropathy
C1859178|Progressive peripheral neuropathy
C1859178|Peripheral neuropathy, progressive
C4039742|Peripheral neuropathy caused by toxin (disorder)
C4039742|Peripheral neuropathy caused by toxin
C3495442|Phantom pain
C3495442|Phantom pain (finding)
C3495442|Phantom limb syndrome
C3495442|Phantom pain (disorder)
C4039352|Peripheral neuropathy due to inflammation
C4039352|Peripheral neuropathy due to inflammation (disorder)
C3276706|SFNP
C3276706|NEUROPATHY, SMALL FIBER
C3276706|Small fibre neuropathy
C3276706|Small fiber neuropathy
C3276706|Small fiber neuropathy (disorder)
C3276706|Small Nerve Fiber Neuropathy
C4040658|Peripheral neuropathy due to metabolic disorder
C4040658|Peripheral neuropathy due to metabolic disorder (disorder)
C0271375|Fourth or trochlear nerve palsy
C0271375|Fourth [trochlear] nerve palsy
C0271375|fourth nerve palsy
C0271375|fourth cranial nerve palsy
C0271375|fourth nerve palsy (diagnosis)
C0271375|IVth nerve paralysis
C0271375|Fourth Nerve Palsies
C0271375|Palsies, Fourth Nerve
C0271375|Palsy, Fourth Nerve
C0271375|Palsies, Trochlear Nerve
C0271375|Palsy, Trochlear Nerve
C0271375|Trochlear Nerve Palsies
C0271375|Trochlear Nerve Disorder
C0271375|IVth Cranial Nerve Disorder
C0271375|Trochlear Nerve Diseases
C0271375|Fourth Cranial Nerve Diseases
C0271375|Trochlear Nerve Disorders
C0271375|Trochlear Nerve Diseases [Disease/Finding]
C0271375|Trochlear Neuropathy
C0271375|Cranial Nerve IV Diseases
C0271375|Palsy;IV nerve
C0271375|Fourth cranial nerve paresis (disorder)
C0271375|Disorder of trochlear nerve
C0271375|Fourth cranial nerve disease (disorder)
C0271375|Fourth cranial nerve disease
C0271375|Superior oblique muscle innervation disorder (disorder)
C0271375|IVth nerve paresis
C0271375|Superior oblique muscle innervation disorder
C0271375|Disorder of trochlear nerve (disorder)
C0271375|Fourth cranial nerve paresis
C0271375|Disorder of cranial nerve 4
C0271375|IVth nerve disorder
C0271375|Trochlear nerve palsy
C0271375|Superior oblique palsy
C0271375|Trochlear nerve paralysis
C0271375|Paresis of fourth cranial nerve
C0271375|IVth nerve palsy
C0271375|Fourth nerve paresis
C0271375|Fourth nerve paralysis
C0271375|Fourth cranial nerve paralysis
C0271375|Fourth cranial nerve disorder
C0271375|Trochlear nerve weakness
C0271375|4th nerve palsy
C0271375|IV nerve palsy
C0271375|Fourth nerve palsy (disorder)
C0271375|Trochlear nerve disease
C0271375|disease (or disorder); cranial nerve, fourth
C0271375|disease (or disorder); trochlear nerve
C0271375|n.trochlearis; paralysis
C0271375|paralysis; cranial nerve, fourth
C0271375|paralysis; trochlear nerve
C0271375|Fourth cranial nerve disease, NOS
C0271375|Fourth cranial nerve disorder, NOS
C0271375|Trochlear nerve disease, NOS
C0271375|Trochlear nerve disorder, NOS
C0271375|IV thnerve palsy
C0270937|Celiac plexus syndrome
C0270937|Solar plexus syndrome
C0270937|Coeliac plexus syndrome
C0270937|Celiac plexus syndrome (disorder)
C0271353|Third cranial nerve disorder
C0271353|Disorder of oculomotor nerve
C0271353|Disorder of oculomotor nerve (disorder)
C0271353|IIIrd nerve disorder
C0271353|Disorder of cranial nerve 3
C0271353|Oculomotor nerve disorder
C0271353|Oculomotor nerve disease
C0271353|Third cranial nerve disease (disorder)
C0271353|Third cranial nerve disease
C0271353|cranial nerve; disorder, third (oculomotor)
C0271353|disease (or disorder); cranial nerve, third (oculomotor)
C0271353|disease (or disorder); nerve, oculomotor
C0271353|n.oculomotorius; disorder
C0271353|Oculomotor nerve disease, NOS
C0271353|Oculomotor nerve disorder, NOS
C0271353|Third cranial nerve disease, NOS
C0271353|Third cranial nerve disorder, NOS
C0152179|Disorders of pneumogastric (10th) nerve
C0152179|Disorders of vagus nerve
C0152179|TENTH CRANIAL NERVE DIS
C0152179|PNEUMOGASTRIC NERVE DIS
C0152179|CRANIAL NERVE X DIS
C0152179|VAGUS NERVE DIS
C0152179|Vagus nerve disorders
C0152179|Vagus Nerve Disease
C0152179|Vagus Nerve Diseases
C0152179|Disorder, Pneumogastric Nerve
C0152179|Disorders, Pneumogastric Nerve
C0152179|Pneumogastric Nerve Disorder
C0152179|Vagus Nerve Disorder
C0152179|Neuropathies, Vagus
C0152179|Neuropathy, Vagus
C0152179|Vagus Neuropathies
C0152179|Disorders of pneumogastric [10th] nerve
C0152179|Tenth Cranial Nerve Diseases
C0152179|Vagus Neuropathy
C0152179|Vagus Nerve Diseases [Disease/Finding]
C0152179|Cranial Nerve X Diseases
C0152179|Pneumogastric Nerve Disorders
C0152179|disorder of vagus nerve (diagnosis)
C0152179|disorder vagus nerve
C0152179|disorder of vagus nerve
C0152179|Disorder of cranial nerve 10
C0152179|Vagus nerve disorder NOS
C0152179|Disorders of the Xth cranial nerve
C0152179|Disorders of the tenth nerve
C0152179|Vagus nerve lesion
C0152179|Disorder of pneumogastric nerve
C0152179|Disorder of the tenth cranial nerve
C0152179|Disorder of vagus nerve (disorder)
C0152179|cranial nerve; disorder, tenth (vagus)
C0152179|disease (or disorder); cranial nerve, tenth (vagus)
C0152179|disease (or disorder); nerve, pneumogastric
C0152179|disease (or disorder); nerve, vagus
C0152179|n.vagus; disorder
C0152179|Disorder of pneumogastric nerve, NOS
C0152179|Disorder of the tenth cranial nerve, NOS
C0152179|Disorder of vagus nerve, NOS
C0152179|Disorder of pneumogastric nerve (disorder)
C0152179|n.pneumogastric; disorder
C0152179|Disorders of 10th nerve
C0152179|Disorders of pneumogastric nerve
C0152179|Disorders of vagal nerve
C0270923|Secondary peripheral neuropathy (disorder)
C0270923|Secondary peripheral neuropathy
C0270923|Secondary peripheral neuropathy, NOS
C0152177|Trigeminal nerve disorders
C0152177|Disorder of trigeminal nerve, unspecified
C0152177|Disorders of trigeminal nerve
C0152177|CRANIAL NERVE V DIS
C0152177|TRIGEMINAL NERVE DIS
C0152177|FIFTH CRANIAL NERVE DIS
C0152177|Trigeminal disorders
C0152177|Trigeminal Nerve Disease
C0152177|Trigeminal Nerve Diseases
C0152177|Trigeminal Nerve Disorder
C0152177|Neuropathies, Trigeminal
C0152177|Neuropathy, Trigeminal
C0152177|Trigeminal Neuropathies
C0152177|Trigeminal nerve dis NOS
C0152177|disorders of 5th cranial nerve
C0152177|Trigeminal Nerve Diseases [Disease/Finding]
C0152177|Cranial Nerve V Diseases
C0152177|Trigeminal Neuropathy
C0152177|Fifth Cranial Nerve Diseases
C0152177|disorder trigeminal nerve
C0152177|disorder of trigeminal nerve
C0152177|disorder of trigeminal nerve (diagnosis)
C0152177|Trigeminal nerve disorder NOS (disorder)
C0152177|Trigeminal nerve disorder NOS
C0152177|Disorder of trigeminal nerve (disorder)
C0152177|Disorder of cranial nerve 5
C0152177|Trigeminal nerve--Diseases
C0152177|Trigeminal nerve disorder, unspecified
C0152177|Disorders of the Vth cranial nerve
C0152177|Disorders of the fifth nerve
C0152177|Disorder of the fifth cranial nerve
C0152177|Trigeminal nerve disorder (disorder)
C0152177|disease (or disorder); cranial nerve, fifth
C0152177|disease (or disorder); trigeminal nerve
C0152177|Disorder of the fifth cranial nerve, NOS
C0152177|Trigeminal nerve disorder, NOS
C0031121|Peripheral neuralgia
C0031121|Peripheral neuralgia (disorder)
C4076016|Disorder of peripheral nervous system co-occurrent with human immunodeficiency virus infection (disorder)
C4076016|Disorder of peripheral nervous system co-occurrent with human immunodeficiency virus infection
C0271355|Sixth or abducens nerve palsy
C0271355|Sixth [abducent] nerve palsy
C0271355|Lateral rectus palsy
C0271355|ABDUCENS NERVE DIS
C0271355|SIXTH CRANIAL NERVE DIS
C0271355|VITH CRANIAL NERVE DIS
C0271355|CRANIAL NERVE VI DIS
C0271355|sixth nerve palsy (diagnosis)
C0271355|sixth nerve palsy
C0271355|sixth cranial nerve palsy
C0271355|Abducens paralysis
C0271355|VIth nerve paralysis
C0271355|Abducens Nerve Disease
C0271355|Abducens Nerve Diseases
C0271355|Abducens Nerve Palsies
C0271355|Palsies, Abducens Nerve
C0271355|Palsy, Abducens Nerve
C0271355|Lateral Rectus Palsies
C0271355|Palsies, Lateral Rectus
C0271355|Palsy, Lateral Rectus
C0271355|Palsies, Sixth Nerve
C0271355|Palsy, Sixth Nerve
C0271355|Sixth Nerve Palsies
C0271355|Palsy, VI Nerve
C0271355|Nerve Palsies, VI
C0271355|Nerve Palsy, VI
C0271355|Palsies, VI Nerve
C0271355|Nerve Palsy, 6th
C0271355|Palsies, 6th Nerve
C0271355|Palsy, 6th Nerve
C0271355|6th Nerve Palsies
C0271355|Nerve Palsies, 6th
C0271355|Abducens Nerve Palsy
C0271355|VIth Cranial Nerve Diseases
C0271355|Cranial Nerve VI Diseases
C0271355|Sixth Cranial Nerve Disorders
C0271355|Sixth Cranial Nerve Diseases
C0271355|Abducens Nerve Diseases [Disease/Finding]
C0271355|Cranial Nerve VI Palsy
C0271355|6th Nerve Palsy
C0271355|VI Nerve Palsy
C0271355|Abducens nerve weakness
C0271355|Sixth cranial nerve weakness
C0271355|Sixth cranial nerve disorder
C0271355|Disorder of abducent nerve
C0271355|Abducens (sixth) nerve palsy
C0271355|Sixth cranial nerve disease
C0271355|Disorder of abducent nerve (disorder)
C0271355|Lateral rectus muscle denervation paresis
C0271355|Abducens nerve paralysis
C0271355|Abducens nerve disorder
C0271355|Sixth cranial nerve paralysis
C0271355|Lateral rectus muscle innervation disorder
C0271355|VIth nerve disorder
C0271355|Lateral rectus muscle denervation paresis (disorder)
C0271355|Lateral rectus muscle innervation disorder (disorder)
C0271355|Abducens nerve paresis
C0271355|Sixth cranial nerve disease (disorder)
C0271355|Sixth nerve palsy (disorder)
C0271355|Disorder of abducens nerve
C0271355|Disorder of cranial nerve 6
C0271355|Sixth nerve paralysis
C0271355|VIth nerve palsy
C0271355|Abducent nerve paralysis
C0271355|Abducens nerve disorder (disorder)
C0271355|Abducens nerve palsy (disorder)
C0271355|Abducens nerve weakness (disorder)
C0271355|disease (or disorder); abducent nerve
C0271355|disease (or disorder); cranial nerve, sixth
C0271355|paralysis; abducent nerve
C0271355|paralysis; cranial nerve, sixth
C0271355|Abducens nerve disease, NOS
C0271355|Abducens nerve disorder, NOS
C0271355|Sixth cranial nerve disease, NOS
C0271355|Sixth cranial nerve disorder, NOS
C0751941|Disorders of glossopharyngeal nerve
C0751941|CRANIAL NERVE IX DIS
C0751941|GLOSSOPHARYNGEAL NERVE DIS
C0751941|NINTH CRANIAL NERVE DIS
C0751941|CRANIAL NERVE VIIII DISEASES
C0751941|Glossopharyngeal nerve disorders
C0751941|Glossopharyngeal Nerve Disease
C0751941|Glossopharyngeal Nerve Diseases
C0751941|Cranial Nerve IX Diseases
C0751941|Cranial Nerve IX Disorders
C0751941|Ninth Cranial Nerve Diseases
C0751941|Glossopharyngeal Nerve Diseases [Disease/Finding]
C0751941|disorder of glossopharyngeal nerve
C0751941|disorder of glossopharyngeal nerve (diagnosis)
C0751941|disorder glossopharyngeal nerve
C0751941|Glossopharyngeal nerve disorder
C0751941|Disorder of cranial nerve 9
C0751941|Glossopharyngeal nerve disorder NOS
C0751941|Disorder of the ninth cranial nerve
C0751941|Disorder of IXth cranial nerve
C0751941|Disorder of ninth nerve
C0751941|Glossopharyngeal nerve lesion
C0751941|Disorder of glossopharyngeal nerve (disorder)
C0751941|cranial nerve; disorder, ninth (glossopharyngeal)
C0751941|disease (or disorder); cranial nerve, ninth (glossopharyngeal)
C0751941|disease (or disorder); nerve, glossopharyngeal
C0751941|n.glossopharyngeus; disorder
C0751941|IX Nerve Disorder
C0751941|Ninth Nerve Disorder
C0015464|Diseases, Facial Nerve
C0015464|Facial Nerve Disease
C0015464|Facial Nerve Diseases
C0015464|Facial nerve disorders
C0015464|Disease, Facial Nerve
C0015464|Disorder of facial nerve, unspecified
C0015464|Disorder of seventh cranial nerve
C0015464|Facial nerve disorder
C0015464|Facial nerve disorder (disorder)
C0015464|Facial neuropathy
C0015464|Disorders of the VIIth cranial nerve
C0015464|Disorders of the seventh nerve
C0015464|Disorder of facial nerve
C0015464|SEVENTH CRANIAL NERVE DIS
C0015464|CRANIAL NERVE VII DIS
C0015464|FACIAL NERVE DIS
C0015464|Disorder, Facial Nerve
C0015464|Disorders, Facial Nerve
C0015464|Facial Neuropathies
C0015464|Neuropathies, Facial
C0015464|Neuropathy, Facial
C0015464|Facial nerve dis NOS
C0015464|disorders of 7th cranial nerve
C0015464|Seventh Cranial Nerve Diseases
C0015464|Cranial Nerve VII Disorders
C0015464|Facial Nerve Diseases [Disease/Finding]
C0015464|Cranial Nerve VII Diseases
C0015464|LMNL of VIIth nerve
C0015464|Facial cranial nerve disorders
C0015464|disorder of facial nerve (diagnosis)
C0015464|disorder facial nerve
C0015464|Facial nerve disorders NOS
C0015464|Facial nerve disorder NOS (disorder)
C0015464|Disorder of facial nerve (disorder)
C0015464|Facial nerve disorder NOS
C0015464|Facial neuropathy (disorder)
C0015464|Disorder of cranial nerve 7
C0015464|Facial nerve--Diseases
C0015464|Facial nerve disorder, unspecified
C0015464|disease (or disorder); cranial nerve, seventh
C0015464|disease (or disorder); facial nerve
C0015464|Disorder of seventh cranial nerve, NOS
C0015464|Facial nerve disorder, NOS
C0015464|Disorder of of seventh cranial nerve, NOS
C0152181|Disorders of hypoglossal (12th) nerve
C0152181|Disorders of hypoglossal nerve
C0152181|HYPOGLOSSAL NERVE DIS
C0152181|CRANIAL NERVE XII DIS
C0152181|TWELFTH CRANIAL NERVE DIS
C0152181|Hypoglossal nerve disorders
C0152181|Hypoglossal Nerve Disease
C0152181|Hypoglossal Nerve Diseases
C0152181|Disorders of 12th cranial nerve
C0152181|Twelfth Cranial Nerve Disorder
C0152181|Cranial Nerve XII Diseases
C0152181|Cranial Nerve XII Disorders
C0152181|Hypoglossal Nerve Diseases [Disease/Finding]
C0152181|Twelfth Cranial Nerve Diseases
C0152181|disorder of hypoglossal nerve (diagnosis)
C0152181|disorder of hypoglossal nerve
C0152181|disorder hypoglossal nerve
C0152181|Hypoglossal nerve disorder
C0152181|Disorder of cranial nerve 12
C0152181|Hypoglossal nerve disorder NOS
C0152181|Disorders of the XIIth cranial nerve
C0152181|Disorders of the twelfth cranial nerve
C0152181|Hypoglossal nerve lesion
C0152181|Disorder of hypoglossal nerve (disorder)
C0152181|Disorder of the twelfth cranial nerve
C0152181|cranial nerve; disorder, twelfth (hypoglossal)
C0152181|disease (or disorder); cranial nerve, twelfth (hypoglossal)
C0152181|disease (or disorder); nerve, hypoglossal
C0152181|n.hypoglossus; disorder
C0152181|Disorder of hypoglossal nerve, NOS
C0152181|Disorder of the twelfth cranial nerve, NOS
C0152181|Disorder of XII Nerve
C0152181|Twelfth Nerve Disorder
C0152181|Disorder of the XII Nerve
C0152181|Disorders of hypoglossal [12th] nerve
C0152181|Disorders of 12th nerve
C0266834|Familial visceral neuropathy
C0266834|Familial visceral neuropathy (disorder)
C0001163|Disorders of acoustic nerve
C0001163|VESTIBULOCOCHLEAR NERVE DIS
C0001163|CRANIAL NERVE VIII DIS
C0001163|EIGHTH CRANIAL NERVE DIS
C0001163|Auditory nerve disorders
C0001163|VIIIth cranial nerve disorders
C0001163|Vestibulocochlear Nerve Disease
C0001163|Vestibulocochlear Nerve Diseases
C0001163|Acoustic nerve disorders
C0001163|Eighth Cranial Nerve Diseases
C0001163|Cranial Nerve VIII Diseases
C0001163|Cranial Nerve VIII Disorders
C0001163|Vestibulocochlear Nerve Diseases [Disease/Finding]
C0001163|disorder of acoustic nerve (diagnosis)
C0001163|Disorder of acoustic nerve
C0001163|Acoustic nerve disorder NOS
C0001163|Acoustic nerve disorder NOS (disorder)
C0001163|Disorder of auditory nerve
C0001163|Disorder of vestibulocochlear nerve
C0001163|Disorder of eighth cranial nerve
C0001163|Disorder of cranial nerve 8
C0001163|Disorder of eighth nerve
C0001163|Disorder of acoustovestibular nerve
C0001163|Disorder of acoustic nerve (disorder)
C0001163|Disorder of the vestibulocochlear nerve
C0001163|auditory nerve; disorder
C0001163|auditory; nerve
C0001163|cranial nerve; disorder, eighth (auditory)
C0001163|disease (or disorder); cranial nerve, eighth (auditory)
C0001163|disease (or disorder); nerve, acoustic
C0001163|disease (or disorder); nerve, auditory
C0001163|disorder; vestibulocochlear nerve
C0001163|disturbance; vestibulocochlear nerve
C0001163|n.vestibulocochlearis; disorder
C0001163|Disorder of acoustic nerve, NOS
C0001163|Disorder of eighth nerve, NOS
C0001163|Disorder of the vestibulocochlear nerve, NOS
C0001163|Acoustic Nerve Disorder
C0001163|Vestibulocochlear Nerve Disorder
C0001163|Disorder of acoustic or eighth nerve
C0495832|Injury of peripheral nerves of thorax
C0495832|peripheral nerve injury of thorax (diagnosis)
C0495832|peripheral nerve injury of thorax
C0495832|peripheral nerve injury thorax
C0495832|injury; nerve, thorax, peripheral
C0677499|radial tunnel syndrome (diagnosis)
C0677499|radial tunnel syndrome
C0677499|Supinator syndrome
C0677499|Radial tunnel syndrome (disorder)
C0677499|Radial tunnel syndrome (supinator syndrome)
C0149940|SCIATIC NERVE DIS
C0149940|Nerve Disease, Sciatic
C0149940|Nerve Diseases, Sciatic
C0149940|Sciatic Nerve Disease
C0149940|Neuropathies, Sciatic
C0149940|Neuropathy, Sciatic
C0149940|Sciatic Neuropathies
C0149940|Sciatic Neuropathy
C0149940|Sciatic Neuropathy [Disease/Finding]
C0149940|Sciatic Nerve Diseases
C0149940|Sciatic nerve neuropathy
C0149940|Sciatic nerve--Diseases
C0149940|Sciatic neuropathy (disorder)
C0149940|disease (or disorder); nerve, sciatic
C0149940|n.ischiadicus; neuropathic
C0149940|neuropathy; sciatic nerve
C0027881|neuronitis
C0393804|Polyneuropathy in disease NOS (disorder)
C0393804|Polyneuropathy in disease NOS
C0477401|Other disorders of peripheral nervous system
C0477401|[X]Other disorders of the peripheral nervous system
C0477401|[X]Other disorders of the peripheral nervous system (disorder)
C0392555|Hypertrophic interstitial neuropathy
C0392555|Onion bulb hypertrophy
C0392555|Hypertrophic interstitial neuropathy (disorder)
C0263899|Radicular syndrome of lower limbs
C0263899|Radicular syndrome of lower limbs (disorder)
C0271348|Strachan's syndrome
C0271348|Strachan's syndrome (diagnosis)
C0271348|Strachan syndrome
C0271348|Amblyopia, neuropathy, orogenital dermatitis syndrome
C0271348|Howes-Pallister-Landor syndrome
C0271348|Strachan's syndrome (disorder)
C0266513|Defective development of cauda equina
C0266513|Defective development of cauda equina (disorder)
C0266513|Defective development of the cauda equina
C0266513|Defective development of the cauda equina (disorder)
C0266513|development; defective, congenital, cauda equina
C0394022|Disorder of nerve repair
C0394022|Disorder of nerve repair (disorder)
C0393866|Injection neuropathy
C0393866|Injection neuropathy (disorder)
C0555208|Fibrolipoma of filum terminale
C0555208|Fibrolipoma of filum terminale (disorder)
C0266516|congenital malformations anomaly of peripheral nervous system
C0266516|congenital anomaly of peripheral nervous system
C0266516|congenital anomaly of peripheral nervous system (diagnosis)
C0266516|Congenital peripheral nervous system anomaly NOS
C0266516|Congenital anomaly of the peripheral nervous system (disorder)
C0266516|Congenital anomaly of the peripheral nervous system
C0266516|Congenital anomaly of the peripheral nervous system, NOS
C1145628|ANS Disease
C1145628|Autonomic Nervous System Diseases
C1145628|Disorders of the autonomic nervous system
C1145628|Autonomic Disease
C1145628|Disorder of autonomic nervous system, unspecified
C1145628|Disorders of autonomic nervous system
C1145628|autonomic disorder
C1145628|Autonomic dysfunction
C1145628|DIS AUTONOMIC NERVOUS SYSTEM
C1145628|AUTONOMIC NERVOUS SYSTEM DIS
C1145628|ANS DIS
C1145628|NERVOUS SYSTEM DIS AUTONOMIC
C1145628|CENTRAL AUTONOMIC NERVOUS SYSTEM DIS
C1145628|AUTONOMIC DIS
C1145628|autonomic nervous system disorder (diagnosis)
C1145628|autonomic nervous system disorder
C1145628|ANS disorder
C1145628|Autonomic nervous system disorders
C1145628|Autonomic nerve dis NEC
C1145628|Disorder of the autonomic nervous system, unspecified
C1145628|Autonomic Central Nervous System Diseases
C1145628|Autonomic Nervous System Diseases [Disease/Finding]
C1145628|ANS Diseases
C1145628|Autonomic Diseases
C1145628|Nervous System Diseases, Autonomic
C1145628|Central Autonomic Nervous System Diseases
C1145628|ANS (Autonomic Nervous System) Diseases
C1145628|AUTONOMIC CNS DIS
C1145628|Autonomic nervous system disorder NOS (disorder)
C1145628|Autonomic nervous system disorder NOS
C1145628|Autonomic nervous system--Diseases
C1145628|Unspecified disorder of autonomic nervous system
C1145628|Disorder of autonomic nervous system (disorder)
C1145628|Disorder of autonomic nervous system
C1145628|Disorder of vegetative system
C1145628|autonomic; nervous system, disorder
C1145628|disease (or disorder); autonomic nervous system
C1145628|disease (or disorder); nervous system, autonomic
C1145628|disease (or disorder); nervous system, vegetative
C1145628|nervous system; disorder, autonomic
C1145628|Disorder of autonomic nervous system, NOS
C1145628|Disorder of vegetative system, NOS
C1278821|Infectious disorder of the peripheral nervous system
C1278821|Infectious disorder of the peripheral nervous system (disorder)
C1278821|Peripheral nerve infection
C1278821|Infectious peripheral neuropathy
C1278821|Infectious disorder of the peripheral nervous system [Ambiguous]
C1278821|Peripheral Nervous System Infectious Disorder
C0270891|ElectroPhys: Nerve plexus disorder
C0270891|Nerve plexus disorder (disorder)
C0270891|Nerve plexus disorder
C0270891|Nerve plexus disorder, NOS
C0751950|NEUROMUSCULAR TRANSM DIS
C0751950|NEUROMUSCULAR JUNCTION DIS
C0751950|Neuromuscular Junction Disease
C0751950|Neuromuscular Junction Diseases
C0751950|Neuromuscular Junction Disorder
C0751950|Neuromuscular Transmission Disorder
C0751950|Neuromuscular Transmission Disorders
C0751950|Neuromuscular Junction Diseases [Disease/Finding]
C0751950|Neuromuscular Junction Disorders
C0751950|Neuromuscular junction disorder (disorder)
C0034931|Dystrophies, Reflex Sympathetic
C0034931|Dystrophy, Reflex Sympathetic
C0034931|Reflex Sympathetic Dystrophies
C0034931|Reflex Sympathetic Dystrophy
C0034931|Shoulder Hand Syndrome
C0034931|Sudeck's Atrophy
C0034931|Sympathetic Dystrophies, Reflex
C0034931|Sympathetic Dystrophy, Reflex
C0034931|Syndrome, Shoulder-Hand
C0034931|Shoulder-Hand Syndromes
C0034931|Syndromes, Shoulder-Hand
C0034931|CRPS TYPE I
C0034931|Reflex sympathetic dystrophy of upper extremity
C0034931|Sudeck's atrophy (diagnosis)
C0034931|shoulder-hand syndrome (diagnosis)
C0034931|shoulder-hand syndrome
C0034931|Complex regional pain syndrome type I of the upper limb
C0034931|Atrophy, Sudek
C0034931|Atrophy, Sudek's
C0034931|Sudeks Atrophy
C0034931|I, CPRS Type
C0034931|Type I, CPRS
C0034931|Reflex Dystrophia, Sympathetic
C0034931|Sympathetic Reflex Dystrophias
C0034931|Unsp rflx sympth dystrph
C0034931|Rflx sym dystrph up limb
C0034931|Sudek's Atrophy
C0034931|CPRS Type I
C0034931|Pain Syndrome Type I, Regional, Complex
C0034931|Complex Regional Pain Syndrome, Type I
C0034931|RSD (Reflex Sympathetic Dystrophy)
C0034931|Syndrome, Reflex Sympathetic Dystrophy
C0034931|Sympathetic Reflex Dystrophia
C0034931|Type I Complex Regional Pain Syndrome
C0034931|Reflex Sympathetic Dystrophy [Disease/Finding]
C0034931|Pain Syndrome Type I, Complex Regional
C0034931|Reflex Sympathetic Dystrophy Syndrome
C0034931|Sudek Atrophy
C0034931|Dystrophy;reflex sympathetic
C0034931|Atrophies, Sudek's
C0034931|CPRS Type Is
C0034931|Is, CPRS Type
C0034931|RSDs (Reflex Sympathetic Dystrophy)
C0034931|Sudek's Atrophies
C0034931|Type Is, CPRS
C0034931|Algodystrophy
C0034931|Sudeck's atrophy (disorder)
C0034931|Reflex sympathetic dystrophy (disorder)
C0034931|Reflex sympathetic dystrophy (& Sudek's atrophy) (disorder)
C0034931|CRPS - Complex regional pain syndrome type I
C0034931|Reflex sympathetic dystrophy (& Sudek's atrophy)
C0034931|Sudek's atrophy (disorder)
C0034931|Shoulder-hand syndrome (disorder)
C0034931|RSD - Reflex sympathetic dystrophy
C0034931|Complex regional pain syndrome type I
C0034931|Algoneurodystrophy
C0034931|complex regional pain syndrome type I of upper limb (diagnosis)
C0034931|Complex regional pain syndrome type I (diagnosis)
C0034931|complex regional pain syndrome type I of upper limb
C0034931|Reflex sympathetic dystrophy of the upper limb
C0034931|Reflex sympathetic dystrophy, unspecified
C0034931|Reflex Neurovascular Dystrophy
C0034931|CRPS I
C0034931|RND
C0034931|RSDS
C0034931|Complex Regional Pain Syndrome I
C0034931|Steinbrocker's syndrome
C0034931|Algodystrophy (disorder)
C0034931|Reflex sympathetic dystrophy of upper extremity (disorder)
C0034931|atrophy; Sudeck
C0034931|Sudeck; atrophy
C0034931|Sudeck
C0034931|hand-shoulder; syndrome
C0034931|shoulder-hand; syndrome
C0034931|syndrome; hand-shoulder
C0034931|syndrome; shoulder-hand
C0034931|Reflex sympathetic dystrophy [Ambiguous]
C0494493|Idiopathic progressive neuropathy
C0494493|idiopathic peripheral neuropathy progressive
C0494493|idiopathic progressive neuropathy (diagnosis)
C0494493|idiopathic; neuropathic, progressive
C0494493|neuropathy; idiopathic, progressive
C0436023|compartment syndrome of buttock
C0436023|compartment syndrome buttock
C0436023|compartment syndrome of buttock (diagnosis)
C0436023|Compartment syndrome, buttock
C0436023|Compartment syndrome, buttock (disorder)
C0436024|compartment syndrome of thigh (diagnosis)
C0436024|Compartment syndrome of thigh
C0436024|Compartment syndrome of thigh (disorder)
C0086957|Scalenus Anticus Syndrome
C0086957|Syndrome, Scalenus Anticus
C0086957|scalenus anticus syndrome (diagnosis)
C0086957|Cervical rib syndrome
C0086957|Cervical rib syndrome (disorder)
C0086957|Scalenus anticus syndrome (disorder)
C0086957|scalenus anticus; syndrome
C0086957|syndrome; scalenus anticus
C0086957|Naffziger's syndrome
C0751932|POSTERIOR TIBIAL NERVE DIS
C0751932|TIBIAL NERVE DIS
C0751932|Nerve Disease, Tibial
C0751932|Nerve Diseases, Tibial
C0751932|Tibial Nerve Disease
C0751932|Internal Popliteal Neuropathies
C0751932|Neuropathies, Internal Popliteal
C0751932|Neuropathy, Internal Popliteal
C0751932|Popliteal Neuropathies, Internal
C0751932|Popliteal Neuropathy, Internal
C0751932|Medial Popliteal Neuropathies
C0751932|Neuropathies, Medial Popliteal
C0751932|Neuropathy, Medial Popliteal
C0751932|Popliteal Neuropathies, Medial
C0751932|Popliteal Neuropathy, Medial
C0751932|Neuropathies, Posterior Tibial
C0751932|Neuropathy, Posterior Tibial
C0751932|Posterior Tibial Neuropathies
C0751932|Tibial Neuropathies, Posterior
C0751932|Tibial Neuropathy, Posterior
C0751932|Neuropathies, Tibial
C0751932|Neuropathy, Tibial
C0751932|Tibial Neuropathies
C0751932|Tibial Neuropathy
C0751932|Tibial Nerve Diseases
C0751932|Tibial Neuropathy [Disease/Finding]
C0751932|Internal Popliteal Neuropathy
C0751932|Posterior Tibial Nerve Diseases
C0751932|Posterior Tibial Neuropathy
C0751932|Medial Popliteal Neuropathy
C0751932|Tibial neuropathy (disorder)
C0751932|Posterior tibial neuropathy (disorder)
C0751932|Tibial neuropathy (disorder) [Ambiguous]
C1275816|Common peroneal nerve paralysis
C1275816|Common peroneal nerve paralysis (disorder)
C0205930|Algoneurodystrophy
C0205930|Algoneurodystrophy, unspecified site
C0205930|Algoneurodystrophy NOS
C0205930|Algoneurodystrophy NOS (disorder)
C0205930|Algoneurodystrophy (disorder)
C0434564|closed dislocation of lumbar vertebra with cauda equina lesion (diagnosis)
C0434564|closed dislocation of lumbar vertebra with cauda equina lesion
C0434564|dislocation vertebra lumbar closed with cauda equina lesion
C0434564|Closed spinal dislocation with cauda equina lesion
C0434564|Closed spinal dislocation with cauda equina lesion (disorder)
C0434571|open dislocation of lumbar vertebra with cauda equina lesion
C0434571|dislocation vertebra open with cauda equina lesion
C0434571|open dislocation of lumbar vertebra with cauda equina lesion (diagnosis)
C0434571|dislocation vertebra lumbar open with cauda equina lesion
C0434571|open dislocation of vertebra with cauda equina lesion
C0434571|Open spinal dislocation with cauda equina lesion
C0434571|Open spinal dislocation with cauda equina lesion (disorder)
C0270907|Acute radial nerve palsy
C0270907|Acute radial nerve palsy (disorder)
C0751922|Median neuropathy (finding)
C0751922|MEDIAN NERVE DIS
C0751922|nerve palsy median
C0751922|median nerve palsy
C0751922|median nerve palsy (diagnosis)
C0751922|Median Nerve Disease
C0751922|Nerve Disease, Median
C0751922|Nerve Diseases, Median
C0751922|Median Neuropathies
C0751922|Median Neuropathy
C0751922|Neuropathies, Median
C0751922|Neuropathy, Median
C0751922|Median Nerve Diseases
C0751922|Median Neuropathy [Disease/Finding]
C0751922|Median neuropathy (disorder)
C0751922|disease (or disorder); median nerve
C0740447|Diabetic peripheral neuropathy (disorder)
C0740447|Diabetic peripheral neuropathy
C0740447|diabetic peripheral neuropathy (diagnosis)
C0553761|Median nerve compression in forearm
C0553761|Median nerve compression in forearm (disorder)
C1384669|lateral popliteal nerve palsy (diagnosis)
C1384669|nerve palsy lateral popliteal
C1384669|nerve palsy common peroneal
C1384669|common peroneal nerve palsy
C1384669|lateral popliteal nerve palsy
C1384669|common peroneal nerve palsy (diagnosis)
C1335029|Non-Neoplastic Peripheral Nervous System Disease
C1335029|Non-Neoplastic Peripheral Nervous System Disorder
C0026849|Muscular dystrophies and other myopathies
C0026849|Other muscular dystrophies and myopathies
C0026849|Muscular dystrophies and other myopathies, unspecified
C0026849|Muscular dystrophy/myopathies
C0026849|Other myopathies and muscular dystrophies
C0026849|Other myopathies and muscular dystrophies (disorder)
C0026849|Muscular dystrophies and other myopathies (disorder)
C0154730|Disorders of other cranial nerves
C0154730|Other cranial nerve disorders
C0154730|Other cranial nerve disorders (disorder)
C0154747|mononeuritis of lower limb (diagnosis)
C0154747|mononeuritis lower limb
C0154747|mononeuritis of lower limb
C0154747|mononeuritis of a lower limb
C0154747|Unspecified mononeuritis of lower limb
C0154747|Mononeuritis leg NOS
C0154747|Mononeuritis;legs
C0154747|Unspecified mononeuritis lower limb (disorder)
C0154747|Mononeuritis lower limb (disorder)
C0154747|Unspecified mononeuritis lower limb
C0154747|Mononeuritis of lower limb (disorder)
C0154747|Mononeuritis of lower limb, unspecified
C0154747|lower limb; mononeuritis
C0154747|mononeuritis; lower limb
C0154747|Mononeuritis of lower limb, NOS
C0154747|mononeuritis of the legs
C0270890|Nerve root and plexus disorders
C0270890|Nerve root and plexus disorder, unspecified
C0270890|nerve root and plexus disorder (diagnosis)
C0270890|nerve root and plexus disorder
C0270890|Nerv root/plexus dis NOS
C0270890|Nerve root or plexus disorder NOS
C0270890|Nerve root or plexus disorder NOS (disorder)
C0270890|Unspecified nerve root and plexus disorder
C0270890|disease (or disorder); plexus
C0435513|Closed fracture of coccyx with complete cauda equina lesion
C0435513|Closed fracture of coccyx with complete cauda equina lesion (disorder)
C0435518|Open fracture of coccyx with complete cauda equina lesion
C0435518|Open fracture of coccyx with complete cauda equina lesion (disorder)
C1960872|Sural neuropathy
C1960872|Sural neuropathy (disorder)
C0435504|Open fracture of sacrum with complete cauda equina lesion
C0435504|Open fracture of sacrum with complete cauda equina lesion (disorder)
C1268588|porphyric polyneuropathy
C1268588|porphyric polyneuropathy (diagnosis)
C1268588|Polyneuropathy in porphyria (disorder)
C1268588|Polyneuropathy in porphyria
C1268588|Porphyric polyneuropathy (disorder)
C0032587|Polyradiculoneuropathies
C0032587|Polyradiculoneuropathy
C0032587|Polyradiculoneuropathy [Disease/Finding]
C0032587|Polyradiculoneuropathy (disorder)
C0394023|Disruption of nerve repair
C0394023|Disruption of nerve repair (disorder)
C0394025|Neuroma of nerve repair
C0394025|Neuroma of nerve repair (disorder)
C0751929|Neuropathies, Superficial Peroneal
C0751929|Peroneal Neuropathies, Superficial
C0751929|Peroneal Neuropathy, Superficial
C0751929|Superficial Peroneal Neuropathies
C0751929|Superficial Peroneal Neuropathy
C0751929|Superficial peroneal nerve neuropathy (disorder)
C0751929|Superficial peroneal nerve lesion
C0751929|Superficial peroneal nerve neuropathy
C0751929|Superficial peroneal nerve disorder
C0751929|Superficial peroneal nerve disorder (disorder)
C0751929|Neuropathy, Superficial Peroneal
C2102996|disorders of peripheral nerve, neuromuscular junction and muscle (diagnosis)
C2102996|disorders of peripheral nerve, neuromuscular junction and muscle
C0442874|Neuropathy
C0442874|nerve disorders
C0442874|nerve disorders (diagnosis)
C0442874|Neuropathy - (NOS)
C0442874|Neuropathy NOS
C0442874|neuropathy (diagnosis)
C0442874|Neuropathy (nerve damage)
C0442874|Neuropathy (disorder)
C0442874|nerve; disorder
C0442874|Neuropathy, NOS
