C0364639|Iron[Mass/volume] in Serum or Plasma
C0428578|Iron level result
C0853169|Blood iron measurement
C1318312|Serum iron measurement
C0373658|Iron binding capacity measurement
C0428579|Iron measurement, urine
C1272108|Plasma iron level 
C0364639|Iron [Mass/volume] in Serum or Plasma
C0364639|Iron SerPl-mCnc
C0364639|Iron:MCnc:Pt:Ser/Plas:Qn
C0364639|Iron:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0853169|Blood iron measurement
C0853169|Blood iron
C1283048|Total iron binding capacity
C1283048|Iron binding capacity total
C1283048|Iron binding capacity.total
C1283048|IBCT
C1283048|Total iron binding capacity measurement
C1283048|Total iron binding capacity measurement (procedure)
C1283048|Iron binding capacity total measurement
C1283048|TIBC - Total iron binding capacity
C1283048|Total iron binding capacity each test
C1283048|tot iron bndng cpct ea.tst
C1318312|serum iron
C1318312|serum iron measurement (lab test)
C1318312|serum iron measurement
C1318312|Serum iron level
C1318312|(Serum iron tests) or (serum iron level) (procedure)
C1318312|(Serum iron tests) or (serum iron level)
C1318312|Serum iron: [tests] or [level] (procedure)
C1318312|Serum iron level (procedure)
C1318312|Serum iron: [tests] or [level]
C1318312|Serum iron measurement (procedure)
C1277709|iron saturation
C1277709|iron saturation (lab test)
C1277709|Transferrin saturation
C1277709|Transferrin Saturation Measurement
C1277709|Transferrin saturation index (procedure)
C1277709|Transferrin saturation index
C1277709|Saturation of iron binding capacity (procedure)
C1277709|Saturation of iron binding capacity
C1277709|Iron Saturation Percent
C1277709|TFRRNSAT
C1277709|Serum Iron to TIBC Ratio
C1277709|Transferrin Iron Saturation
C1277709|Iron Binding Capacity Saturation
C1277709|Percentage iron saturation
C1277709|Serum transferrin saturation
C0202106|Unsaturated Iron Binding Capacity Measurement
C0202106|Unsaturated iron binding capacity
C0202106|Unsaturated iron binding capacity (procedure)
C0202106|Transferrin saturation measurement
C0202106|Iron/total iron binding capacity ratio measurement
C0202106|Unsaturated iron binding capacity measurement (procedure)
C0202106|Iron, percent saturation, calculated
C0202106|IBCU
C0202106|Iron, percent saturation measurement
C0202106|UIBC - Unsaturated iron binding capacity
C1990893|Iron binding capacity.unsaturated &#x7C; bld-ser-plas
C1990892|Iron binding capacity &#x7C; bld-ser-plas
C0373658|Iron binding capacity
C0373658|IBC
C0373658|Measurement of iron binding capacity
C0373658|IRON BINDING TEST
C0373658|IBC - Iron binding capacity
C0373658|Iron binding capacity measurement
C0428579|Urine iron
C0428579|Urine iron (& level)
C0428579|Iron - urine
C0428579|Urine iron (& level) (procedure)
C0428579|Iron measurement, urine
C0428579|Urine iron level
C0428579|Iron measurement, urine (procedure)
C1278240|24 hour urine iron output (procedure)
C1278240|24 hour urine iron output
C1278240|24 hour urine iron output measurement (procedure)
C1278240|24 hour urine iron output measurement
C1272108|Plasma iron level
C1272108|Plasma iron level (procedure)
