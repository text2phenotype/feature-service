Position|above|epi||epigastric|above, on top of
Position|above|supra||suprapubic|above, upward
Position|around|peri||periodontis|around, surrounding
Position|around|circum||circumoral|around
Position|away|ana|||away, up, apart
Position|away|ab|||away from
Position|away|apo||apocrine|away from, separate
Position|back|retro||retroflexion|backward
Position|between|inter||intercostal|between
Position|down|infra||infraspinous|down
Position|front|pre|||before, in front of
Position|front|ante||anteversion|forward, in front of
Position|front|front||frontonasal|forehead, front
Position|in|in|||in, not
Position|in|en|||in
Position|in|eso||esotropia|inward 
Position|lateral|laterali||laterality|of, at, toward, or from side(s)
Position|lateral||lateral|laterality|of, at, toward, or from side(s)
Position|left|levo||levocardia|left
Position|near|par|||near, beside
Position|out|ex||| 
Position|out|exo||exostosis|out
Position|out|ec|||out, outward
Position|out|ecto||ectomorph|out, outward
Position|out|extra||extracorporeal|outside
Position|right|dextro|||
Position|same|ipsi||ipsilateral|same
Position|through|dia||dialysis|complete, through
Position|through|trans||transcutaneous|accross, through
Position|through|per|||through
Position|toward|ad||adduction|toward
Position|under|sub||subcutaneous|under, below
Position|within|end||endarterectomy|within
Position|within|endo||endometriosis|within
Position|within|intra||intracerebral|within
