C0009555|Complete Blood Count
C0545131|complete blood count with differential (lab test)
C0545131|CBC with differential
C0545131|complete blood count with differential
C0545131|Blood Cell Count with Differential
C0545131|CBC with Diff
C0009555|complete blood count
C0009555|CBC
C0009555|Blood Counts, Complete
C0009555|Complete Blood Counts
C0009555|Count, Complete Blood
C0009555|Counts, Complete Blood
C0009555|Full blood count
C0009555|CBC (complete blood count)
C0009555|complete blood count (CBC)
C0009555|complete blood count (CBC) (lab test)
C0009555|FBC
C0009555|Test;full blood count
C0009555|Full blood count NOS (procedure)
C0009555|Full blood count NOS
C0009555|Full blood count (procedure)
C0009555|blood cell count
C0009555|FBC - Full blood count
C0009555|Complete blood count (procedure)
C0009555|Complete blood count, NOS
C0009555|CBC, NOS
C0009555|Blood Count, Complete
C0523113|blood blast count
C0523113|blood blast count (lab test)
C0523113|Blast Count
C0523113|BLAST
C0523113|Blasts
C0523113|Blast cells
C0523113|Blast cells NOS
C0523113|Blast count, blood
C0523113|Blast count, blood (procedure)
C0523113|Blast count procedure
C2698870|Precursor Plasma Cell Count
C2698870|Precursor Plasma Cells
C2698870|PLSPCE
C2698870|Plasmablast
C2698029|Mature Plasma Cell Count
C2698029|Mature Plasma Cells
C2698029|Plasmacytes
C2698029|PLSMCE
C2827509|Eosinophilic Metamyelocyte Count
C2827509|Eosinophilic Metamyelocytes
C2827509|EOSMM
C2827509|Metamyelocytes.eosinophilic
C2827510|Eosinophilic Myelocyte Count
C2827510|Eosinophilic Myelocytes
C2827510|EOSMYL
C2827511|Neutrophilic Metamyelocyte Count
C2827511|Neutrophilic Metamyelocytes
C2827511|NEUTMM
C2827512|Neutrophilic Myelocyte Count
C2827512|Neutrophilic Myelocytes
C2827512|NEUTMY
C0014772|Count, Erythrocyte
C0014772|Counts, Erythrocyte
C0014772|Erythrocyte Count
C0014772|Erythrocyte Counts
C0014772|Erythrocyte Numbers
C0014772|Red blood cell count
C0014772|RBC count NOS (procedure)
C0014772|erythrocyte count (lab test)
C0014772|RBC count
C0014772|Red Cell Count
C0014772|Red blood cell count (procedure)
C0014772|RBC count NOS
C0014772|Red blood cell count NOS (procedure)
C0014772|Red blood cell count NOS
C0014772|Erythrocytes
C0014772|RBC
C0014772|Red Blood Cells
C0014772|Erythrocyte Number
C0014772|Blood Cell Count, Red
C0014772|Whole Blood Erythrocytic Cell Counts
C0014772|RBC - Red blood cell count
C0014772|Red Blood Cell Count measurement
C0518015|Haemoglobin
C0518015|Haem
C0518015|Hemoglobin Measurement
C0518015|hemoglobin
C0518015|hemoglobin measurement (lab test)
C0518015|Test;haemoglobin
C0518015|BLOOD COUNT HEMOGLOBIN
C0518015|Hemoglobin level
C0518015|Measurement of hemoglobin (Hgb)
C0518015|Hemoglobin determination (procedure)
C0518015|Hemoglobin determination
C0518015|Haemoglobin determination
C0518015|HGB
C0518015|Blood count; hemoglobin (Hgb)
C0518015|FHGB
C0518015|Free Hemoglobin
C0518015|Hemoglobin determination, NOS
C0518015|Haemoglobin determination, NOS
C0518015|Test;hemoglobin
C0518015|haemoglobin test
C0518015|hemoglobin test
C0018935|Hct
C0018935|Erythrocyte Volumes, Packed
C0018935|Hematocrit
C0018935|Hematocrits
C0018935|Packed Erythrocyte Volume
C0018935|Packed Erythrocyte Volumes
C0018935|Packed Red Cell Volume
C0018935|Packed Red-Cell Volumes
C0018935|Red-Cell Volume, Packed
C0018935|Red-Cell Volumes, Packed
C0018935|Volume, Packed Erythrocyte
C0018935|Volume, Packed Red-Cell
C0018935|Volumes, Packed Erythrocyte
C0018935|Volumes, Packed Red-Cell
C0018935|Haematocrit
C0018935|Hematocrit procedure
C0018935|hematocrit (lab test)
C0018935|Hematocrit Measurement
C0018935|BLOOD COUNT HEMATOCRIT
C0018935|Measurement of hematocrit (Hct)
C0018935|Packed cell volume (observable entity)
C0018935|Haematocrit - PCV - NOS
C0018935|Packed cell volume
C0018935|Haematocrit (observable entity)
C0018935|Haematocrit (procedure)
C0018935|Hematocrit - PCV - NOS
C0018935|Haematocrit - PCV - NOS (procedure)
C0018935|Hematocrit - PCV - NOS (procedure)
C0018935|hematocrit packed cell volume (lab test)
C0018935|hematocrit packed cell volume
C0018935|EVF
C0018935|PCV
C0018935|Erythrocyte Volume Fraction
C0018935|Blood count; hematocrit (Hct)
C0018935|Packed Red-Cell Volume
C0018935|Erythrocyte Volume, Packed
C0018935|Whole Blood Hematocrit Test
C0018935|Hematocrit determination
C0018935|Haematocrit - PCV
C0018935|Hct - Haematocrit
C0018935|Hct - Hematocrit
C0018935|Hematocrit - PCV
C0018935|Haematocrit determination
C0018935|Hematocrit determination (procedure)
C0018935|Packed cell volume measurement (procedure)
C0018935|Packed cell volume measurement
C0023508|White Blood Cell Count
C0023508|Count, Leukocyte
C0023508|Counts, Leukocyte
C0023508|Leukocyte Count
C0023508|Leukocyte Counts
C0023508|Leukocyte Numbers
C0023508|Number, Leukocyte
C0023508|Numbers, Leukocyte
C0023508|White Blood Cell Count procedure
C0023508|leukocyte count (lab test)
C0023508|WBC count
C0023508|White blood cell count (procedure)
C0023508|Leukocytes
C0023508|White Blood Cells
C0023508|WBC
C0023508|White cells
C0023508|Leukocyte count NOS
C0023508|White blood cell count NOS
C0023508|White blood cell analysis
C0023508|Leucocyte count
C0023508|Leukocyte Number
C0023508|Blood Cell Count, White
C0023508|Whole Blood Leukocyte Counts
C0023508|WBC - White blood cell count
C0023508|WCC - White blood cell count
C0023508|White blood cell count - observation
C2097083|complete blood count with manual differential and indices (lab test)
C2097083|CBC with manual differential and indices
C2097083|manual CBC with differential and indices
C2097083|complete blood count with manual differential and indices
C2030595|hemogram indices (lab test)
C2030595|hemogram indices
C2984931|Myeloid to Erythroid Ratio Measurement
C2984931|MYPCERPC
C2984931|Myeloid/Erythroid Ratio
C3272957|Immature Plasma Cell Count
C3272957|Immature Plasma Cells
C3272957|PLSIMCE
C0200694|Measurement of total hemoglobin concentration and hematocrit (procedure)
C0200694|Hemoglobin and hematocrit determination
C0200694|Measurement of total hemoglobin concentration and hematocrit
C0200694|Measurement of total haemoglobin concentration and haematocrit
C0200694|Hemoglobin and hematocrit determination (procedure)
C0200694|Haemoglobin and haematocrit determination
C0200694|H & H determination
C0200694|total hemoglobin concentration and hematocrit
C0200694|total hemoglobin concentration and hematocrit (lab test)
C0200694|Haemoglobin and hematocrit determination
C2228885|mean corpuscular diameter (MCD)
C2228885|mean corpuscular diameter (MCD) (lab test)
C2228885|mean corpuscular diameter
C2228299|erythrocyte volume distribution width (RDW)
C2228299|RBC volume distribution width (RDW)
C2228299|erythrocyte volume distribution width (RDW) (lab test)
C2228299|RBC volume distribution width
C0883120|Hemoglobin & Hematocrit panel
C0883120|hemoglobin and hematocrit panel (lab test)
C0883120|hemoglobin and hematocrit panel
C0369183|Mean cell haemoglobin
C0369183|MCH - NOS (procedure)
C0369183|Erythrocyte Mean Corpuscular Hemoglobin
C0369183|Erythrocyte Mean Corpuscular Hemoglobin Test
C0369183|mean corpuscular hemoglobin (MCH)
C0369183|mean corpuscular hemoglobin (MCH) (lab test)
C0369183|Mean corpuscular haemoglobin (MCH) - NOS (procedure)
C0369183|MCH
C0369183|MCH - NOS
C0369183|Mean corpuscular hemoglobin (MCH) - NOS
C0369183|Mean cell haemoglobin (& level)
C0369183|Mean corpuscular haemoglobin (MCH) - NOS
C0369183|Mean cell haemoglobin (& level) (procedure)
C0369183|Mean cell hemoglobin (& level)
C0369183|Mean corpuscular hemoglobin NOS
C0369183|Mean cell hemoglobin
C0369183|Mean corpuscular haemoglobin NOS
C0369183|Mean corpuscular hemoglobin NOS (procedure)
C0369183|Ery. Mean Corpuscular Hemoglobin
C0369183|Mean corpuscular hemoglobin
C0369183|Mean corpuscular haemoglobin
C0369183|Mean corpuscular hemoglobin determination
C0369183|MCH determination
C0369183|MCH - Mean cell haemoglobin
C0369183|MCH - Mean cell hemoglobin
C0369183|Mean corpuscular haemoglobin determination
C0369183|MCH - Mean corpuscular haemoglobin
C0369183|MCH - Mean corpuscular hemoglobin
C0369183|Mean corpuscular hemoglobin determination (procedure)
C1948043|Erythrocyte Mean Corpuscular Volume
C1948043|Erythrocyte Mean Corpuscular Volume Measurement
C1948043|mean corpuscular volume (MCV) (lab test)
C1948043|mean corpuscular volume (MCV)
C1948043|mean corpuscular volume
C1948043|Ery. Mean Corpuscular Volume
C1948043|RBC Mean Corpuscular Volume
C1948043|MCV
C1948043|Erythrocytes Mean Corpuscular Volume
C2030597|CBC with platelet count
C2030597|CBC with platelet count (lab test)
C4031906|cbc automated
C4031906|automated CBC (lab test)
C4031906|automated CBC
C0200665|Mean platelet volume
C0200665|mean platelet volume (MPV) (lab test)
C0200665|mean platelet volume (MPV)
C0200665|MPV
C0200665|Mean Platelet Volume Measurement
C0200665|Volumes, Mean Platelet
C0200665|Platelet Volumes, Mean
C0200665|Platelet Volume, Mean
C0200665|Volume, Mean Platelet
C0200665|Mean Platelet Volumes
C0200665|MPV - Mean platelet volume
C0200665|Platelet mean volume (observable entity)
C0200665|Platelet mean volume
C0200665|Platelet mean volume determination
C0200665|Platelet mean volume determination (procedure)
C4054355|Neutrophils Band Form/ Neutrophils
C4054355|NEUTBNE
C4054355|Neutrophils Band Form to Neutrophils Ratio Measurement
C4054477|Monocytoid Cells/Leukocytes
C4054477|Monocytoid Cells to Leukocytes Ratio Measurement
C4054477|MOCYCELE
C4054040|NEUTSGNE
C4054040|Neutrophils, Segmented/Neutrophils
C4054040|Segmented Neutrophils to Neutrophils Ratio Measurement
C0200629|complete blood count with manual differential
C0200629|complete blood count with manual differential (lab test)
C0200629|CBC with manual differential
C0200629|Complete blood count with white cell differential, manual
C0200629|Complete blood count with white cell differential, manual (procedure)
C0200630|CBC with automated differential
C0200630|CBC with automated differential (lab test)
C0200630|Complete blood count with white cell differential, automated
C0200630|Complete blood count with white cell differential, automated (procedure)
C0200631|Hemogram
C0200631|Complete blood count without differential
C0200631|CBC without differential
C0200631|Haemogram
C0200631|Complete blood count without differential (procedure)
C0032181|Blood Platelet Counts
C0032181|Blood Platelet Numbers
C0032181|Count, Blood Platelet
C0032181|Count, Platelet
C0032181|Counts, Blood Platelet
C0032181|Counts, Platelet
C0032181|Number, Blood Platelet
C0032181|Number, Platelet
C0032181|Numbers, Blood Platelet
C0032181|Numbers, Platelet
C0032181|Platelet Count
C0032181|Platelet Count, Blood
C0032181|Platelet Counts
C0032181|Platelet Counts, Blood
C0032181|Platelet Number, Blood
C0032181|Platelet Numbers
C0032181|Platelet Numbers, Blood
C0032181|platelets
C0032181|platelet count (lab test)
C0032181|Platelet count NOS (procedure)
C0032181|Platelet count NOS
C0032181|Platelet count (procedure)
C0032181|PLAT
C0032181|Anucleated Thrombocytes
C0032181|Thrombocyte count
C0032181|Platelet Number
C0032181|Blood Platelet Count
C0032181|Blood Platelet Number
C0032181|Whole Blood Platelet Counts
C0032181|Plt - Platelet count
C0032181|Platelet count - observation
C0032181|Platelet Count measurement
C1879889|Blood Cell Count Ratio Measurement
