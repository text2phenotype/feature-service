C1305855|Body mass index
C0005893|Body mass index procedure
C4229017|Normal BMI
C0424671|Body mass index 30+ obesity
C1561729|Body mass index (BMI) 40 or greater, adult
C2724372|Body Mass Index (BMI), documented (PV)
C2240399|Encounter for body mass index [BMI]
C0578022|Finding of body mass index
C1305855|Quetelet index
C1305855|Body mass index
C1305855|BMI
C1305855|body mass index (physical finding)
C1305855|Quetelet index (observable entity)
C1305855|Body mass index - observation
C1305855|Body mass index (observable entity)
C1305855|BMI - Body mass index
C1305855|Body mass index, NOS
C1305855|Body mass index [dup] (observable entity)
C2227318|BMI ___ percentile
C2227318|body mass index percentile (physical finding)
C2227318|body mass index percentile
C0578022|Observation of body mass index
C0578022|Finding of body mass index (finding)
C0578022|Finding of body mass index
C0424670|Weight for height
C0424670|Weight for height (observable entity)
C0424670|Ponderal index
C3695134|body mass index screening score (physical finding)
C3695134|body mass index screening score
C0231255|Body mass index decreased
C0231255|body mass index decreased (physical finding)
C0231255|body mass index low (physical finding)
C0231255|body mass index low
C0231255|Decreased body mass index
C0231255|Low body mass index
C0231255|Decreased body mass index (finding)
C0231253|Body mass index normal
C0231253|Normal body mass index (physical finding)
C0231253|Normal body mass index
C0231253|Normal body mass index (finding)
C0231254|Body mass index increased
C0231254|Increased body mass index
C0231254|body mass index increased (physical finding)
C0231254|body mass index high
C0231254|body mass index high (physical finding)
C0231254|Increase in body mass index
C0231254|Increased body mass index (finding)
C2911062|Body Mass Index, pediatric
C2911062|Body mass index (BMI) pediatric
C2911062|body mass index pediatric
C2911062|body mass index, pediatric (physical finding)
C0005893|Body Mass Index
C0005893|Index, Body Mass
C0005893|Quetelets Index
C0005893|Quetelet's Index
C0005893|Quetelet Index
C0005893|Body mass index procedure
C0005893|Index, Quetelet
C0424671|Body mass index 30+ - obesity
C0424671|Obesity (BMI>30)
C0424671|Body mass index 30+ - obesity (finding)
C0424671|BMI 30+ - obesity
C2362324|Childhood obesity
C2362324|Childhood obesity (disorder)
C2362324|Obesity in Children
C2362324|Pediatric Obesity
C2362324|Obesity, Pediatric
C2362324|Childhood obesity BMI 95-100 percentile
C2362324|childhood obesity (diagnosis)
C2362324|Pediatric Obesity [Disease/Finding]
C2362324|Obesity in adolescence
C2362324|Obesity, Adolescent
C2362324|Onset Obesity, Childhood
C2362324|Obesity, Infantile
C2362324|Obesity, Child
C2362324|Obesity, Infant
C2362324|Obesity, Childhood
C2362324|Obesity, Childhood Onset
C2362324|Infantile Obesity
C2362324|Child Obesity
C2362324|Infant Obesity
C2362324|Childhood Onset Obesity
C2362324|Adolescent Obesity
C2362324|Obesity in Childhood
C2921312|BMI 40.0-44.9, adult
C2921312|Body Mass Index 40.0-44.9, adult
C2921313|Body Mass Index 45.0-49.9, adult
C2921313|BMI 45.0-49.9, adult
C2921314|BMI 50.0-59.9, adult
C2921314|Body Mass Index 50.0-59.9, adult
C2921315|Body Mass Index 60.0-69.9, adult
C2921315|BMI 60.0-69.9, adult
C2921316|BMI 70 and over, adult
C2921316|Body Mass Index 70 and over, adult
C2977643|Body mass index (BMI) 40.0-44.9, adult
C2977644|Body mass index (BMI) 45.0-49.9, adult
C2977645|Body mass index (BMI) 50-59.9 , adult
C2977646|Body mass index (BMI) 60.0-69.9, adult
C2977647|Body mass index (BMI) 70 or greater, adult
C2724372|BODY MASS INDEX DOCD
C2724372|Body Mass Index (BMI), documented (PV)
C2724372|BODY MASS INDEX DOCUMENTED
C2911038|Body mass index (BMI) 19 or less, adult
C2911039|Body mass index (BMI) 20-29, adult
C2911050|Body mass index (BMI) 30-39, adult
C1561729|Body Mass Index 40 and over, adult
C1561729|Body mass index (BMI) 40 or greater, adult
C2240399|BODY MASS INDEX
C2240399|Body mass index [BMI]
C2240399|Encounter for body mass index [BMI]
C2240399|Body mass index [BMI] (Z68)
C1561711|BMI between 19-24,adult
C1561711|Body Mass Index between 19-24, adult
C1561717|Body Mass Index between 25-29, adult
C1561728|Body Mass Index between 30-39, adult
C1561710|BMI less than 19,adult
C1561710|Body Mass Index less than 19, adult
C1319441|Body mass index 40+ - morbidly obese
C1319441|Obese class III
C1319441|Body mass index 40+ - severely obese (finding)
C1319441|Body mass index 40+ - severely obese
C0587773|Body mass index less than 20 (finding)
C0587773|Body mass index less than 20
C0587773|BMI less than 20
C0424672|Body mass index 25-29 - overweight (finding)
C0424672|Body mass index index 25-29 - overweight
C0424672|Body mass index 25-29 - overweight
C0424672|Body mass index index 25-29 - overweight (finding)
C0424672|BMI 25-29 - overweight
C1445936|Body mass index 20-24 - normal (finding)
C1445936|Body mass index 20-24 - normal
C0424674|Body mass index high K/M2
C0424674|Body mass index high K/M2 (finding)
C0424673|Body mass index low K/M2
C0424673|Body mass index low K/M2 (finding)
C0424675|Body mass index normal K/M2 (finding)
C0424675|Body mass index normal K/M2
