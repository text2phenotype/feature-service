C0237154|Sharing contaminated personal items
C0237154|Homelessness
C0237154|Homeless
C0032854|Poverty
C2911663|Encounter due to homelessness
C0237154|homeless
C0237154|Homelessness
C0237154|homeless (history)
C0237154|Lack (of);housing
C0237154|Housing lack NOS (finding)
C0237154|Living on the street
C0237154|Housing lack NOS
C0237154|Housing lack
C0237154|Homeless (finding)
C0237154|(Housing lack) or (homeless) (finding)
C0237154|(Housing lack) or (homeless)
C0237154|Living on the street (finding)
C0237154|lack of housing (history)
C0237154|lack of housing
C0237154|Housing lack (finding)
C0237154|housing; lack of
C0237154|lack of; housing
C0237154|lack of; shelter
C0237154|shelter; lack of
C1550450|Transient
C1550450|Living Arrangement - Transient
C1550451|Nomadic
C0425241|Homeless family
C0425241|Homeless family (finding)
C0425241|homeless family (history)
C0425242|Homeless single person
C0425242|Homeless single person (finding)
C0425242|homeless individual
C0425242|homeless individual (history)
C0425242|Single homeless person
C0557220|Living rough
C0557220|living rough (history)
C0557220|Living rough (finding)
C0038077|Squatter
C0038077|Illegal tennant
C0038077|Lives in squat (finding)
C0038077|[Squatter] or [illegal tennant]
C0038077|Lives in squat
C0038077|[Squatter] or [illegal tennant] (environment)
C0038077|Squatter (history)
C0038077|homeless - lives in squat
C0038077|Squatters
C1956419|Illegal migrant
C1956419|Illegal migrant (finding)
C0217846|Vagabond
C0217846|Tramps
C0217846|Social migrant (finding)
C0217846|Tramp
C0217846|Tramp (life style)
C0217846|Social migrant
C0217846|Tramp (life style) [Ambiguous]
C1287167|Finding of temporary shelter arrangements
C1287167|Finding of temporary shelter arrangements (finding)
C1287167|Temporary shelter arrangements - finding
C0870659|Homeless Mentally Ill
C0870659|Mentally Ill Homeless
C0032855|Area, Poverty
C0032855|Areas, Poverty
C0032855|Poverty Area
C0032855|Poverty Areas
C0032854|Poverty
C0032854|Poverty status
C0032854|Low Income
C0032854|Poor
C0032854|Financially poor
C0032854|Financially poor (finding)
C0032854|Social problem - poverty
C0032854|Economic deprivation
C0032854|Pauper
C0032854|Severe lack of money
C0032854|Living in poverty
C3539555|extreme poverty (history)
C3539555|Extreme poverty
C0557161|destitution
C0557161|destitution (history)
C0557161|Destitute
C0557161|Destitute (finding)
C2184145|living in poverty conditions (history)
C2184145|living in poverty conditions
C2184145|lives in poverty conditions
C2911663|Homelessness
C2911663|Encounter due to homelessness
C1394678|homelessness; problem
C1394678|problem; homelessness
C1399807|care providing; lack of housing
C0687129|[V]Lack of housing (context-dependent category)
C0687129|Lack of housing
C0687129|Encounter due to vagabond status
C0687129|[V]Tramp
C0687129|[V]Social transient
C0687129|[V]Lack of housing
C0687129|[V]Hobo
C0687129|[V]Lack of housing (situation)
C0687129|[V]Vagabond
C0687129|[V]Social migrant
C0687129|hobo
C0687129|transient
C0687129|Transients
C0687129|Tramps
C0687129|Hobos
C0687129|Social migrants
C0687129|Vagabonds
C1410737|vagebond
C0026093|Migrant
C0026093|Nomad
C0026093|Nomads
C0026093|Migrant (person)
C0026093|Migrants
