C0010294|Creatinine
C0201975|Creatinine
C1561535|Creatinine
C0201975|Creatinine measurement
C0239150|Creatinine low
C0428279|Finding of creatinine level
C0428279|Creatinine level
C0428279|Creatinine level in blood
C0555149|Creatinine in sample (finding)
C0742904|creatinine rising
C0201975|Creatinine measurement
C0201976|Creatinine measurement, serum (procedure)
C0236408|CHEM-7 Creatinine Measurement
C0010294|Creatinine
C0010294|4H-Imidazol-4-one, 2-amino-1,5-dihydro-1-methyl-
C0010294|Creatinine [Chemical/Ingredient]
C0010294|Creatinine (substance)
C0062932|1-carboxyethyl-2-iminoimidazolidine
C0062932|1H-Imidazole-1-propanoic acid, 2-amino-4,5-dihydro-
C0062932|homocyclocreatine
C0062932|1-carboxyethyl-2-imino-imidazolidine
C0666701|NA 22598A
C0666701|NA-22598A
C0666701|NA22598A
C0482524|Creatinine [Mass/volume] in 24 hour Urine --pre 2 mg dexamethasone PO 2.5 day high dose q6h
C0482524|Creatinine^pre 2 mg dexamethasone PO 2.5 day high dose q6h:MCnc:24H:Urine:Qn
C0482524|Creatinine^pre 2 mg dexamethasone Oral 2.5 day high dose q6h:Mass Concentration:24 hours:Urine:Quantitative
C0482524|Creat pre 2 mg Dex high 24h Ur-mCnc
C1543983|Creatinine [Mass/volume] in Serum or Plasma --10 hours post XXX challenge
C1543983|Creatinine^10H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543983|Creatinine^10H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543983|Creat 10h p chal SerPl-mCnc
C1543998|Creatinine [Mass/volume] in Urine --1.5 hours post XXX challenge
C1543998|Creatinine^1.5H post XXX challenge:MCnc:Pt:Urine:Qn
C1543998|Creatinine^1 1/2 hour post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1543998|Creat 1.5h p chal Ur-mCnc
C1542940|Creatinine^1H pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542940|Creatinine [Moles/volume] in Serum or Plasma --1 hour pre XXX challenge
C1542940|Creat 1h pre chal SerPl-sCnc
C1542940|Creatinine^1 hour pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544117|Creatinine^10H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544117|Creatinine [Moles/volume] in Serum or Plasma --10 hours post XXX challenge
C1544117|Creatinine^10H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544117|Creat 10h p chal SerPl-sCnc
C1544120|Creatinine^18H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544120|Creatinine [Moles/volume] in Serum or Plasma --18 hours post XXX challenge
C1544120|Creat 18h p chal SerPl-sCnc
C1544120|Creatinine^18H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544231|Creatinine^3H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544231|Creatinine [Mass/volume] in Serum or Plasma --3 hours post XXX challenge
C1544231|Creatinine^3 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544231|Creat 3h p chal SerPl-mCnc
C1544242|Creatinine [Moles/volume] in Serum or Plasma --1 hour post XXX challenge
C1544242|Creatinine^1H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544242|Creatinine^1 hour post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544242|Creat 1h p chal SerPl-sCnc
C1986128|Creatinine &#x7C; XXX
C1986123|Creatinine &#x7C; Stool
C1543979|Creatinine^5.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543979|Creatinine [Mass/volume] in Serum or Plasma --5.5 hours post XXX challenge
C1543979|Creatinine^5.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543979|Creat 5.5h p chal SerPl-mCnc
C1543987|Creatinine [Mass/volume] in Serum or Plasma --2 days post XXX challenge
C1543987|Creatinine^2D post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543987|Creat 2D p chal SerPl-mCnc
C1543987|Creatinine^2 days post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544004|Creatinine^4.5H post XXX challenge:MCnc:Pt:Urine:Qn
C1544004|Creatinine [Mass/volume] in Urine --4.5 hours post XXX challenge
C1544004|Creatinine^4.5 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544004|Creat 4.5h p chal Ur-mCnc
C1544137|Creatinine^4.5H post XXX challenge:SCnc:Pt:Urine:Qn
C1544137|Creatinine [Moles/volume] in Urine --4.5 hours post XXX challenge
C1544137|Creatinine^4.5 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544137|Creat 4.5h p chal Ur-sCnc
C1544229|Creatinine [Mass/volume] in Serum or Plasma --2 hours post XXX challenge
C1544229|Creatinine^2H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544229|Creatinine^2 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544229|Creat 2h p chal SerPl-mCnc
C1544230|Creatinine [Mass/volume] in Serum or Plasma --2.5 hours post XXX challenge
C1544230|Creatinine^2.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544230|Creatinine^2 1/2 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544230|Creat 2.5h p chal SerPl-mCnc
C0363589|Creatinine^48H post 2 mg dexamethasone PO 2.5 day high dose q6h:MCnc:24H:Urine:Qn
C0363589|Creatinine [Mass/volume] in 24 hour Urine --48 hours post 2 mg dexamethasone PO 2.5 day high dose q6h
C0363589|Creatinine^48H post 2 mg dexamethasone Oral 2.5 day high dose q6h:Mass Concentration:24 hours:Urine:Quantitative
C0363589|Creat 48h p 2 mg Dex 24h Ur-mCnc
C1543973|Creatinine^45M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543973|Creatinine [Mass/volume] in Serum or Plasma --45 minutes post XXX challenge
C1543973|Creat 45M p chal SerPl-mCnc
C1543973|Creatinine^45M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543995|Creatinine [Mass/volume] in Urine --baseline
C1543995|Creat BS Ur-mCnc
C1543995|Creatinine^baseline:MCnc:Pt:Urine:Qn
C1543995|Creatinine^baseline:Mass Concentration:Point in time:Urine:Quantitative
C1986126|Creatinine &#x7C; Urine and Serum or Plasma
C1543990|Creatinine [Mass/volume] in Urine --pre XXX challenge
C1543990|Creatinine^pre XXX challenge:MCnc:Pt:Urine:Qn
C1543990|Creat pre chal Ur-mCnc
C1543990|Creatinine^pre XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1542942|Creatinine [Moles/volume] in Serum or Plasma --30 minutes pre XXX challenge
C1542942|Creat 30M pre chal SerPl-sCnc
C1542942|Creatinine^30M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542942|Creatinine^30 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544141|Creatinine^8H post XXX challenge:SCnc:Pt:Urine:Qn
C1544141|Creatinine [Moles/volume] in Urine --8 hours post XXX challenge
C1544141|Creatinine^8 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544141|Creat 8h p chal Ur-sCnc
C0482518|Creatinine^24H post 40 ug corticotropin IM BID 3 day:MCnc:24H:Urine:Qn
C0482518|Creatinine [Mass/volume] in 24 hour Urine --24 hours post 40 ug corticotropin IM BID 3 day
C0482518|Creatinine^24 hours post 40 ug corticotropin Intramuscular BID 3 day:Mass Concentration:24 hours:Urine:Quantitative
C0482518|Creat 1D p 40 ug ACTH IM 24h Ur-mCnc
C1543981|Creatinine^8H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543981|Creatinine [Mass/volume] in Serum or Plasma --8 hours post XXX challenge
C1543981|Creatinine^8 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543981|Creat 8h p chal SerPl-mCnc
C1546313|Creatinine [Mass/volume] in Serum or Plasma --2.25 hours post XXX challenge
C1546313|Creatinine^2.25H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1546313|Creatinine^2.25H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1546313|Creat 2.25h p chal SerPl-mCnc
C1543982|Creatinine^9H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543982|Creatinine [Mass/volume] in Serum or Plasma --9 hours post XXX challenge
C1543982|Creatinine^9H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543982|Creat 9h p chal SerPl-mCnc
C1543986|Creat 18h p chal SerPl-mCnc
C1543986|Creatinine^18H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543986|Creatinine [Mass/volume] in Serum or Plasma --18 hours post XXX challenge
C1543986|Creatinine^18H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544119|Creatinine^16H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544119|Creat 16h p chal SerPl-sCnc
C1544119|Creatinine [Moles/volume] in Serum or Plasma --16 hours post XXX challenge
C1544119|Creatinine^16H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544121|Creatinine^2D post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544121|Creatinine [Moles/volume] in Serum or Plasma --2 days post XXX challenge
C1544121|Creat 2D p chal SerPl-sCnc
C1544121|Creatinine^2 days post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544240|Creat BS SerPl-sCnc
C1544240|Creatinine^baseline:SCnc:Pt:Ser/Plas:Qn
C1544240|Creatinine [Moles/volume] in Serum or Plasma --baseline
C1544240|Creatinine^baseline:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544245|Creatinine [Moles/volume] in Serum or Plasma --2.5 hours post XXX challenge
C1544245|Creatinine^2.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544245|Creatinine^2 1/2 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544245|Creat 2.5h p chal SerPl-sCnc
C3534241|Creatinine in peritoneal fluid &#x7C; Peritoneal fluid and serum or plasma
C1986115|Creatinine &#x7C; cerebral spinal fluid
C1986127|Creatinine &#x7C; vitreous fluid
C1986111|Creatinine &#x7C; amniotic fluid
C1544135|Creatinine^3.5H post XXX challenge:SCnc:Pt:Urine:Qn
C1544135|Creatinine [Moles/volume] in Urine --3.5 hours post XXX challenge
C1544135|Creatinine^3.5 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544135|Creat 3.5h p chal Ur-sCnc
C1986122|Creatinine &#x7C; pleural fluid
C1544000|Creatinine^2.5H post XXX challenge:MCnc:Pt:Urine:Qn
C1544000|Creatinine [Mass/volume] in Urine --2.5 hours post XXX challenge
C1544000|Creatinine^2 1/2 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544000|Creat 2.5h p chal Ur-mCnc
C1544007|Creatinine^6H post XXX challenge:MCnc:Pt:Urine:Qn
C1544007|Creatinine [Mass/volume] in Urine --6 hours post XXX challenge
C1544007|Creatinine^6 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544007|Creat 6h p chal Ur-mCnc
C1544123|Creatinine^7D post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544123|Creat 7D p chal SerPl-sCnc
C1544123|Creatinine [Moles/volume] in Serum or Plasma --7 days post XXX challenge
C1544123|Creatinine^7 days post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544134|Creatinine [Moles/volume] in Urine --3 hours post XXX challenge
C1544134|Creatinine^3H post XXX challenge:SCnc:Pt:Urine:Qn
C1544134|Creatinine^3 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544134|Creat 3h p chal Ur-sCnc
C1986112|Creatinine &#x7C; bld-ser-plas
C0482520|Creatinine [Mass/volume] in 24 hour Urine --48 hours post 500 ug dexamethasone PO 2.5 day low dose q6h
C0482520|Creatinine^48H post 500 ug dexamethasone PO 2.5 day low dose q6h:MCnc:24H:Urine:Qn
C0482520|Creatinine^48H post 500 ug dexamethasone Oral 2.5 day low dose q6h:Mass Concentration:24 hours:Urine:Quantitative
C0482520|Creat 48h p 500 ug Dex 24h Ur-mCnc
C1543975|Creatinine^3.75H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543975|Creatinine [Mass/volume] in Serum or Plasma --3.75 hours post XXX challenge
C1543975|Creatinine^3.75H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543975|Creat 3.75h p chal SerPl-mCnc
C1544005|Creatinine^5H post XXX challenge:MCnc:Pt:Urine:Qn
C1544005|Creatinine [Mass/volume] in Urine --5 hours post XXX challenge
C1544005|Creatinine^5 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544005|Creat 5h p chal Ur-mCnc
C1544008|Creatinine^8H post XXX challenge:MCnc:Pt:Urine:Qn
C1544008|Creatinine [Mass/volume] in Urine --8 hours post XXX challenge
C1544008|Creatinine^8 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544008|Creat 8h p chal Ur-mCnc
C1542943|Creatinine [Moles/volume] in Serum or Plasma --45 minutes post XXX challenge
C1542943|Creat 45M p chal SerPl-sCnc
C1542943|Creatinine^45M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542943|Creatinine^45M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0550308|Creat BS DiafP-mCnc
C0550308|Creatinine^baseline:MCnc:Pt:Dial fld prt:Qn
C0550308|Creatinine [Mass/volume] in Peritoneal dialysis fluid --baseline
C0550308|Creatinine^baseline:Mass Concentration:Point in time:Peritoneal dialysis fluid:Quantitative
C1543970|Creatinine [Mass/volume] in Serum or Plasma --1 hour pre XXX challenge
C1543970|Creat 1h pre chal SerPl-mCnc
C1543970|Creatinine^1H pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543970|Creatinine^1 hour pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543989|Creat 7D p chal SerPl-mCnc
C1543989|Creatinine^7D post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543989|Creatinine [Mass/volume] in Serum or Plasma --7 days post XXX challenge
C1543989|Creatinine^7 days post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543992|Creatinine [Mass/volume] in Urine --1.5 hours pre XXX challenge
C1543992|Creatinine^1.5H pre XXX challenge:MCnc:Pt:Urine:Qn
C1543992|Creat 1.5h pre chal Ur-mCnc
C1543992|Creatinine^1 1/2 hour pre XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1542945|Creatinine^4H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542945|Creatinine [Moles/volume] in Serum or Plasma --4 hours post XXX challenge
C1542945|Creatinine^4 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542945|Creat 4h p chal SerPl-sCnc
C1831325|Creat sp1 p chal Ur-mCnc
C1831325|Creatinine [Mass/volume] in Urine --1st specimen post XXX challenge
C1831325|Creatinine^1st specimen post XXX challenge:MCnc:Pt:Urine:Qn
C1831325|Creatinine^1st specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1831326|Creatinine^3rd specimen post XXX challenge:MCnc:Pt:Urine:Qn
C1831326|Creat sp3 p chal Ur-mCnc
C1831326|Creatinine [Mass/volume] in Urine --3rd specimen post XXX challenge
C1831326|Creatinine^3rd specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C0482522|Creatinine^pre 40 ug corticotropin IM 3 day:MCnc:24H:Urine:Qn
C0482522|Creatinine [Mass/volume] in 24 hour Urine --pre 40 ug corticotropin IM 3 day
C0482522|Creatinine^pre 40 ug corticotropin Intramuscular 3 day:Mass Concentration:24 hours:Urine:Quantitative
C0482522|Creat pre 40 ug ACTH IM 24h Ur-mCnc
C1543996|Creatinine^30M post XXX challenge:MCnc:Pt:Urine:Qn
C1543996|Creat 30M p chal Ur-mCnc
C1543996|Creatinine [Mass/volume] in Urine --30 minutes post XXX challenge
C1543996|Creatinine^30 minutes post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544002|Creatinine [Mass/volume] in Urine --3.5 hours post XXX challenge
C1544002|Creatinine^3.5H post XXX challenge:MCnc:Pt:Urine:Qn
C1544002|Creatinine^3.5 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544002|Creat 3.5h p chal Ur-mCnc
C1542944|Creatinine [Moles/volume] in Serum or Plasma --3.5 hours post XXX challenge
C1542944|Creatinine^3.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542944|Creatinine^3.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542944|Creat 3.5h p chal SerPl-sCnc
C1544125|Creatinine [Moles/volume] in Urine --1.5 hours pre XXX challenge
C1544125|Creat 1.5h pre chal Ur-sCnc
C1544125|Creatinine^1.5H pre XXX challenge:SCnc:Pt:Urine:Qn
C1544125|Creatinine^1 1/2 hour pre XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544131|Creatinine^1.5H post XXX challenge:SCnc:Pt:Urine:Qn
C1544131|Creatinine [Moles/volume] in Urine --1.5 hours post XXX challenge
C1544131|Creatinine^1 1/2 hour post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544131|Creat 1.5h p chal Ur-sCnc
C1544248|Creatinine^6H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544248|Creatinine [Moles/volume] in Serum or Plasma --6 hours post XXX challenge
C1544248|Creatinine^6 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544248|Creat 6h p chal SerPl-sCnc
C3534240|Creatinine in pleural fluid &#x7C; Bld-Ser-Plas
C1986117|Creatinine &#x7C; dialysis fluid
C1986114|Creatinine &#x7C; body fluid
C1986121|Creatinine &#124; peritoneal fluid
C1986121|Creatinine &#x7C; peritoneal fluid
C0482519|Creatinine^48H post 40 ug corticotropin IM BID 3 day:MCnc:24H:Urine:Qn
C0482519|Creatinine [Mass/volume] in 24 hour Urine --48 hours post 40 ug corticotropin IM BID 3 day
C0482519|Creatinine^48H post 40 ug corticotropin Intramuscular BID 3 day:Mass Concentration:24 hours:Urine:Quantitative
C0482519|Creat 2D p 40 ug ACTH IM 24h Ur-mCnc
C1543994|Creatinine [Mass/volume] in Urine --30 minutes pre XXX challenge
C1543994|Creat 30M pre chal Ur-mCnc
C1543994|Creatinine^30M pre XXX challenge:MCnc:Pt:Urine:Qn
C1543994|Creatinine^30 minutes pre XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1543999|Creatinine^2H post XXX challenge:MCnc:Pt:Urine:Qn
C1543999|Creatinine [Mass/volume] in Urine --2 hours post XXX challenge
C1543999|Creatinine^2 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1543999|Creat 2h p chal Ur-mCnc
C1544133|Creatinine [Moles/volume] in Urine --2.5 hours post XXX challenge
C1544133|Creatinine^2.5H post XXX challenge:SCnc:Pt:Urine:Qn
C1544133|Creatinine^2 1/2 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544133|Creat 2.5h p chal Ur-sCnc
C1544249|Creat 1D p chal SerPl-sCnc
C1544249|Creatinine^1D post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544249|Creatinine [Moles/volume] in Serum or Plasma --1 day post XXX challenge
C1544249|Creatinine^1 day post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0482523|Creatinine [Mass/volume] in 24 hour Urine --pre 500 ug dexamethasone PO 2.5 day low dose q6h
C0482523|Creatinine^pre 500 ug dexamethasone PO 2.5 day low dose q6h:MCnc:24H:Urine:Qn
C0482523|Creatinine^pre 500 ug dexamethasone Oral 2.5 day low dose q6h:Mass Concentration:24 hours:Urine:Quantitative
C0482523|Creat pre 500 ug Dex 24h Ur-mCnc
C1543972|Creatinine [Mass/volume] in Serum or Plasma --30 minutes pre XXX challenge
C1543972|Creatinine^30M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543972|Creat 30M pre chal SerPl-mCnc
C1543972|Creatinine^30 minutes pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544226|Creat 30M p chal SerPl-mCnc
C1544226|Creatinine [Mass/volume] in Serum or Plasma --30 minutes post XXX challenge
C1544226|Creatinine^30M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544226|Creatinine^30 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544233|Creatinine [Mass/volume] in Serum or Plasma --6 hours post XXX challenge
C1544233|Creatinine^6H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544233|Creatinine^6 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544233|Creat 6h p chal SerPl-mCnc
C1986120|Creatinine &#x7C; gastric fluid
C1986125|Creatinine &#x7C; urine
C1544115|Creatinine^8H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544115|Creatinine [Moles/volume] in Serum or Plasma --8 hours post XXX challenge
C1544115|Creatinine^8 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544115|Creat 8h p chal SerPl-sCnc
C1544118|Creatinine [Moles/volume] in Serum or Plasma --12 hours post XXX challenge
C1544118|Creatinine^12H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544118|Creatinine^12 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544118|Creat 12h p chal SerPl-sCnc
C1544124|Creatinine^pre XXX challenge:SCnc:Pt:Urine:Qn
C1544124|Creat pre chal Ur-sCnc
C1544124|Creatinine [Moles/volume] in Urine --pre XXX challenge
C1544124|Creatinine^pre XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544243|Creatinine [Moles/volume] in Serum or Plasma --1.5 hours post XXX challenge
C1544243|Creatinine^1.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544243|Creatinine^1 1/2 hour post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544243|Creat 1.5h p chal SerPl-sCnc
C2924902|Creatinine reduction ratio &#x7C; Bld-Ser-Plas
C1543976|Creatinine [Mass/volume] in Serum or Plasma --4 hours post XXX challenge
C1543976|Creatinine^4H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543976|Creatinine^4 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543976|Creat 4h p chal SerPl-mCnc
C1542939|Creat 1.5h pre chal SerPl-sCnc
C1542939|Creatinine [Moles/volume] in Serum or Plasma --1.5 hours pre XXX challenge
C1542939|Creatinine^1.5H pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542939|Creatinine^1 1/2 hour pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544126|Creatinine^1H pre XXX challenge:SCnc:Pt:Urine:Qn
C1544126|Creatinine [Moles/volume] in Urine --1 hour pre XXX challenge
C1544126|Creat 1h pre chal Ur-sCnc
C1544126|Creatinine^1 hour pre XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544116|Creatinine [Moles/volume] in Serum or Plasma --9 hours post XXX challenge
C1544116|Creatinine^9H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544116|Creatinine^9H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544116|Creat 9h p chal SerPl-sCnc
C1544246|Creatinine [Moles/volume] in Serum or Plasma --3 hours post XXX challenge
C1544246|Creatinine^3H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544246|Creatinine^3 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544246|Creat 3h p chal SerPl-sCnc
C1831329|Creat sp6 p chal Ur-mCnc
C1831329|Creatinine [Mass/volume] in Urine --6th specimen post XXX challenge
C1831329|Creatinine^6th specimen post XXX challenge:MCnc:Pt:Urine:Qn
C1831329|Creatinine^6th specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C2357242|Creatinine &#x7C; Dialysis fluid + Serum or Plasma
C2357241|Creatinine &#x7C; Dialysis fluid peritoneal + Serum or Plasma
C1831341|Creatinine [Mass/volume] in Urine --5th specimen post XXX challenge
C1831341|Creat sp5 p chal Ur-mCnc
C1831341|Creatinine^5th specimen post XXX challenge:MCnc:Pt:Urine:Qn
C1831341|Creatinine^5th specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544003|Creatinine^4H post XXX challenge:MCnc:Pt:Urine:Qn
C1544003|Creatinine [Mass/volume] in Urine --4 hours post XXX challenge
C1544003|Creatinine^4 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544003|Creat 4h p chal Ur-mCnc
C1544234|Creat 1D p chal SerPl-mCnc
C1544234|Creatinine [Mass/volume] in Serum or Plasma --1 day post XXX challenge
C1544234|Creatinine^1D post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544234|Creatinine^1 day post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C3169509|Creatinine^post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C3169509|Creat p chal SerPl-sCnc
C3169509|Creatinine^post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3169509|Creatinine [Moles/volume] in Serum or Plasma --post XXX challenge
C0482521|Creatinine^72H post 40 ug corticotropin IM BID 3 day:MCnc:24H:Urine:Qn
C0482521|Creatinine [Mass/volume] in 24 hour Urine --72 hours post 40 ug corticotropin IM BID 3 day
C0482521|Creatinine^72H post 40 ug corticotropin Intramuscular BID 3 day:Mass Concentration:24 hours:Urine:Quantitative
C0482521|Creat 72h p 40 ug ACTH IM 24h Ur-mCnc
C1543991|Creatinine [Mass/volume] in Urine --2.25 hours pre XXX challenge
C1543991|Creatinine^2.25H pre XXX challenge:MCnc:Pt:Urine:Qn
C1543991|Creatinine^2.25H pre XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1543991|Creat 2.25h pre chal Ur-mCnc
C1544009|Creatinine^1D post XXX challenge:MCnc:Pt:Urine:Qn
C1544009|Creatinine [Mass/volume] in Urine --1 day post XXX challenge
C1544009|Creat 1D p chal Ur-mCnc
C1544009|Creatinine^1 day post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544227|Creatinine^1H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544227|Creatinine [Mass/volume] in Serum or Plasma --1 hour post XXX challenge
C1544227|Creatinine^1 hour post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544227|Creat 1h p chal SerPl-mCnc
C1543985|Creatinine [Mass/volume] in Serum or Plasma --16 hours post XXX challenge
C1543985|Creat 16h p chal SerPl-mCnc
C1543985|Creatinine^16H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543985|Creatinine^16H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544130|Creatinine [Moles/volume] in Urine --1 hour post XXX challenge
C1544130|Creatinine^1H post XXX challenge:SCnc:Pt:Urine:Qn
C1544130|Creatinine^1 hour post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544130|Creat 1h p chal Ur-sCnc
C1544132|Creatinine^2H post XXX challenge:SCnc:Pt:Urine:Qn
C1544132|Creatinine [Moles/volume] in Urine --2 hours post XXX challenge
C1544132|Creatinine^2 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544132|Creat 2h p chal Ur-sCnc
C1544136|Creatinine^4H post XXX challenge:SCnc:Pt:Urine:Qn
C1544136|Creatinine [Moles/volume] in Urine --4 hours post XXX challenge
C1544136|Creatinine^4 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544136|Creat 4h p chal Ur-sCnc
C1544232|Creatinine [Mass/volume] in Serum or Plasma --5 hours post XXX challenge
C1544232|Creatinine^5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544232|Creatinine^5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544232|Creat 5h p chal SerPl-mCnc
C1986113|Creatinine &#x7C; blood arterial
C1543988|Creatinine^4D post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543988|Creatinine [Mass/volume] in Serum or Plasma --4 days post XXX challenge
C1543988|Creat 4D p chal SerPl-mCnc
C1543988|Creatinine^4 days post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543993|Creatinine [Mass/volume] in Urine --1 hour pre XXX challenge
C1543993|Creatinine^1H pre XXX challenge:MCnc:Pt:Urine:Qn
C1543993|Creat 1h pre chal Ur-mCnc
C1543993|Creatinine^1 hour pre XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544001|Creatinine [Mass/volume] in Urine --3 hours post XXX challenge
C1544001|Creatinine^3H post XXX challenge:MCnc:Pt:Urine:Qn
C1544001|Creatinine^3 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544001|Creat 3h p chal Ur-mCnc
C1544247|Creatinine^5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544247|Creatinine [Moles/volume] in Serum or Plasma --5 hours post XXX challenge
C1544247|Creatinine^5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544247|Creat 5h p chal SerPl-sCnc
C2925718|Creat sp2 Ur-mCnc
C2925718|Creatinine^2nd specimen:MCnc:Pt:Urine:Qn
C2925718|Creatinine [Mass/volume] in Urine --2nd specimen
C2925718|Creatinine^2nd specimen:Mass Concentration:Point in time:Urine:Quantitative
C1986118|Creatinine &#124; dialysis fluid peritoneal
C1986118|Creatinine &#x7C; dialysis fluid peritoneal
C1543968|Creat pre chal SerPl-mCnc
C1543968|Creatinine^pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543968|Creatinine [Mass/volume] in Serum or Plasma --pre XXX challenge
C1543968|Creatinine^pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543977|Creatinine^4.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543977|Creatinine [Mass/volume] in Serum or Plasma --4.5 hours post XXX challenge
C1543977|Creatinine^4.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543977|Creat 4.5h p chal SerPl-mCnc
C1542941|Creatinine^45M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542941|Creatinine [Moles/volume] in Serum or Plasma --45 minutes pre XXX challenge
C1542941|Creat 45M pre chal SerPl-sCnc
C1542941|Creatinine^45M pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544138|Creatinine^5H post XXX challenge:SCnc:Pt:Urine:Qn
C1544138|Creatinine [Moles/volume] in Urine --5 hours post XXX challenge
C1544138|Creatinine^5 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544138|Creat 5h p chal Ur-sCnc
C1544140|Creatinine^6H post XXX challenge:SCnc:Pt:Urine:Qn
C1544140|Creatinine [Moles/volume] in Urine --6 hours post XXX challenge
C1544140|Creatinine^6 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544140|Creat 6h p chal Ur-sCnc
C1544225|Creat BS SerPl-mCnc
C1544225|Creatinine [Mass/volume] in Serum or Plasma --baseline
C1544225|Creatinine^baseline:MCnc:Pt:Ser/Plas:Qn
C1544225|Creatinine^baseline:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544228|Creatinine [Mass/volume] in Serum or Plasma --1.5 hours post XXX challenge
C1544228|Creatinine^1.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544228|Creatinine^1 1/2 hour post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544228|Creat 1.5h p chal SerPl-mCnc
C1544006|Creatinine^5.5H post XXX challenge:MCnc:Pt:Urine:Qn
C1544006|Creatinine [Mass/volume] in Urine --5.5 hours post XXX challenge
C1544006|Creatinine^5.5 hours post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1544006|Creat 5.5h p chal Ur-mCnc
C1544127|Creatinine [Moles/volume] in Urine --30 minutes pre XXX challenge
C1544127|Creatinine^30M pre XXX challenge:SCnc:Pt:Urine:Qn
C1544127|Creat 30M pre chal Ur-sCnc
C1544127|Creatinine^30 minutes pre XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544142|Creatinine [Moles/volume] in Urine --1 day post XXX challenge
C1544142|Creat 1D p chal Ur-sCnc
C1544142|Creatinine^1D post XXX challenge:SCnc:Pt:Urine:Qn
C1544142|Creatinine^1 day post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1831324|Creatinine^2nd specimen post XXX challenge:MCnc:Pt:Urine:Qn
C1831324|Creatinine [Mass/volume] in Urine --2nd specimen post XXX challenge
C1831324|Creat sp2 p chal Ur-mCnc
C1831324|Creatinine^2nd specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1543971|Creatinine [Mass/volume] in Serum or Plasma --45 minutes pre XXX challenge
C1543971|Creat 45M pre chal SerPl-mCnc
C1543971|Creatinine^45M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543971|Creatinine^45M pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543974|Creatinine [Mass/volume] in Serum or Plasma --3.5 hours post XXX challenge
C1543974|Creatinine^3.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543974|Creatinine^3.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543974|Creat 3.5h p chal SerPl-mCnc
C1543997|Creatinine^1H post XXX challenge:MCnc:Pt:Urine:Qn
C1543997|Creatinine [Mass/volume] in Urine --1 hour post XXX challenge
C1543997|Creatinine^1 hour post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C1543997|Creat 1h p chal Ur-mCnc
C1543978|Creatinine [Mass/volume] in Serum or Plasma --5.25 hours post XXX challenge
C1543978|Creatinine^5.25H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543978|Creatinine^5.25H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543978|Creat 5.25h p chal SerPl-mCnc
C1542938|Creatinine^pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542938|Creatinine [Moles/volume] in Serum or Plasma --pre XXX challenge
C1542938|Creat pre chal SerPl-sCnc
C1542938|Creatinine^pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544139|Creatinine^5.5H post XXX challenge:SCnc:Pt:Urine:Qn
C1544139|Creatinine [Moles/volume] in Urine --5.5 hours post XXX challenge
C1544139|Creatinine^5.5 hours post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544139|Creat 5.5h p chal Ur-sCnc
C1544244|Creatinine^2H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544244|Creatinine [Moles/volume] in Serum or Plasma --2 hours post XXX challenge
C1544244|Creatinine^2 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544244|Creat 2h p chal SerPl-sCnc
C1986124|Creatinine &#x7C; synovial fluid
C1543969|Creatinine^1.5H pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543969|Creat 1.5h pre chal SerPl-mCnc
C1543969|Creatinine [Mass/volume] in Serum or Plasma --1.5 hours pre XXX challenge
C1543969|Creatinine^1 1/2 hour pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544129|Creatinine [Moles/volume] in Urine --30 minutes post XXX challenge
C1544129|Creatinine^30M post XXX challenge:SCnc:Pt:Urine:Qn
C1544129|Creat 30M p chal Ur-sCnc
C1544129|Creatinine^30 minutes post XXX challenge:Substance Concentration:Point in time:Urine:Quantitative
C1544241|Creatinine^30M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544241|Creat 30M p chal SerPl-sCnc
C1544241|Creatinine [Moles/volume] in Serum or Plasma --30 minutes post XXX challenge
C1544241|Creatinine^30 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1543980|Creatinine^6.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543980|Creatinine [Mass/volume] in Serum or Plasma --6.5 hours post XXX challenge
C1543980|Creatinine^6.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543980|Creat 6.5h p chal SerPl-mCnc
C1543984|Creatinine [Mass/volume] in Serum or Plasma --12 hours post XXX challenge
C1543984|Creatinine^12H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1543984|Creatinine^12 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543984|Creat 12h p chal SerPl-mCnc
C1544122|Creatinine^4D post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544122|Creatinine [Moles/volume] in Serum or Plasma --4 days post XXX challenge
C1544122|Creat 4D p chal SerPl-sCnc
C1544122|Creatinine^4 days post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544128|Creat BS Ur-sCnc
C1544128|Creatinine^baseline:SCnc:Pt:Urine:Qn
C1544128|Creatinine [Moles/volume] in Urine --baseline
C1544128|Creatinine^baseline:Substance Concentration:Point in time:Urine:Quantitative
C1831327|Creatinine^4th specimen post XXX challenge:MCnc:Pt:Urine:Qn
C1831327|Creatinine [Mass/volume] in Urine --4th specimen post XXX challenge
C1831327|Creat sp4 p chal Ur-mCnc
C1831327|Creatinine^4th specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative
C0299232|2-amino-2-imidazolin-4-one
C0299232|2-iminoimidazolidin-4-one
C0082119|2-amino-5-hydroxy-1-methylimidazol-4(5H)-one
C0082119|creatol
C0082119|5-hydroxycreatinine
C0056742|1-carboxymethyl-2-iminoimidazolidine
C0056742|cyclocreatine
C0655900|5,7-DHT-CR
C0655900|5,7-dihydroxytryptamine creatinine
C4044173|1-(4-aminobutyl)-2-iminoimidazolidin-4-one
C0201976|serum creatinine
C0201976|Serum Creatinine Measurement
C0201976|Creatinine measurement, serum (procedure)
C0201976|serum creatinine level
C0201976|serum creatinine measurement (lab test)
C0201976|Creatinine.serum
C0201976|Serum creatinine (& level) (procedure)
C0201976|Creatinine - serum
C0201976|Serum creatinine NOS (procedure)
C0201976|Serum creatinine NOS
C0201976|Serum creatinine (& level)
C0201976|Serum Creatinine Test
C0201976|Creatinine measurement, serum
C1318439|Urine Creatinine Measurement
C1318439|urine creatinine measurement (lab test)
C1318439|urine creatinine
C1318439|creatinine level
C1318439|Creatinine urine
C1318439|Urine creatinine (& level) (procedure)
C1318439|Urine creatinine (& level)
C1318439|Creatinine - urine
C1318439|Creatinine measurement, urine
C1318439|Urine creatinine measurement (procedure)
C1318439|Urine creatinine level
C4050528|Creatinine^overnight dwell:SCnc:Pt:Dial fld prt:Qn
C4050528|Creat DiafP-sCnc
C4050528|Creatinine^overnight dwell:Substance Concentration:Point in time:Peritoneal dialysis fluid:Quantitative
C4050528|Creatinine [Moles/volume] in Peritoneal dialysis fluid --overnight dwell
C0010295|Salt, Creatinine Sulfate
C0010295|Sulfate Salt, Creatinine
C0010295|Creatinine Sulfate Salt
C0765512|2-amino-1,5-dihydro-1-methyl-4H-imidazol-4-one cpd with 3-(2-aminoethyl)-1H-indol-5-ol sulfate
C0765512|serotonin-creatinine sulfate
C0765512|5-hydroxytryptamine creatinine sulphate
C0765512|5-HTQ
C0765512|creatinine sulfate - serotonin
C0765512|creatinine sulfate, serotonin drug combination
C0765512|5-hydroxytryptamine creatinine sulfate
C0201975|Creatinine measurement
C0201975|Creatinine; blood
C0201975|Blood creatinine
C0201975|Creatinine
C0201975|Test;creatinine
C0201975|CREATININE BLOOD
C0201975|Blood creatinine level
C0201975|Measurement of creatinine
C0201975|Cr
C0201975|lab-based chem measurements creatinine
C0201975|measurement of creatinine (lab test)
C0201975|CREAT
C0201975|blood creatinine level (lab test)
C0201975|Creatinine measurement (procedure)
C0201975|Creatinine measurement, NOS
C0201975|ASSAY OF CREATININE
C0201975|creatinine test
C2732591|Urea, electrolytes and creatinine measurement
C2732591|Measurement of urea, sodium, potassium, chloride, bicarbonate and creatinine
C2732591|Measurement of urea, sodium, potassium, chloride, bicarbonate and creatinine (procedure)
C2732591|lab-based chem measure urea, na, potassium chloride, bicarbonate, creatinine
C2732591|measurement of urea, sodium, potassium chloride, bicarbonate, and creatinine
C2732591|measurement of urea, sodium, potassium chloride, bicarbonate, and creatinine (lab test)
C2981749|Urinary Creatinine Assay
C2981751|Serum Creatinine Assay
C1278055|plasma creatinine measurement
C1278055|Plasma creatinine level
C1278055|Plasma creatinine level (procedure)
C1278055|plasma creatinine
C1278055|Plasma creatinine measurement (lab test)
C1278055|Plasma creatinine measurement (procedure)
C0201977|urine creatinine 12-hour
C0201977|12-hour urine creatinine measurement
C0201977|12-hour urine creatinine measurement (lab test)
C0201977|12-hour creatinine level
C0201977|Creatinine measurement, 12 hour urine
C0201977|Creatinine measurement, 12 hour urine (procedure)
C3694999|creatinine concentration (serum or plasma)
C3694999|serum or plasma creatinine concentration (lab test)
C3694999|serum or plasma creatinine concentration
C3694393|lab-based chem measurements creatinine clearance - glomerular filtration (lab test)
C3694393|lab-based chem measurements creatinine clearance - glomerular filtration
C0373594|Creatinine; other source
C0373594|CREATININE OTHER SOURCE
C0373594|ASSAY OF URINE CREATININE
C0373595|Creatinine; clearance
C0373595|Creatinine renal clearance
C0373595|Measurement of renal clearance of creatinine
C0373595|Creatinine clearance test
C0373595|Creatinine clearance test (procedure)
C0373595|Measurement of renal clearance of creatinine (procedure)
C0373595|Creatinine clearance measurement
C0373595|Creatinine renal clearance measurement (procedure)
C0373595|Creatinine clearance-glom filt
C0373595|Creatinine clearance study (procedure)
C0373595|Creatinine renal clearance measurement
C0373595|Creatinine clearance
C0373595|Creatinine clearance study
C0373595|CREATCLR
C0373595|renal function creatinine clearance
C0373595|creatinine renal clearance (procedure)
C0428279|Finding of creatinine level
C0428279|lab-based chem measurements creatinine level finding
C0428279|creatinine level finding (lab test)
C0428279|creatinine level finding
C0428279|Creatinine level
C0428279|Creatinine level - finding
C0428279|Finding of creatinine level (finding)
C0523586|Creatinine challenge tests
C0523586|Creatinine challenge tests (procedure)
C1278053|Corrected plasma creatinine level
C1278053|Corrected plasma creatinine level (procedure)
C1278053|Corrected plasma creatinine measurement (procedure)
C1278053|Corrected plasma creatinine measurement
C1261396|Fluid sample creatinine measurement
C1261396|Body Fluid Creatinine Test
C1261396|Creatinine measurement, body fluid
C1261396|Fluid sample creatinine measurement (procedure)
C1261396|Fluid sample creatinine level
C1293927|Measurement of ratio of analyte to creatinine (procedure)
C1293927|Measurement of ratio of analyte to creatinine
C0428613|Calcium to Creatinine Ratio Measurement
C0428613|Calcium/creatinine ratio
C0428613|Calcium/creatinine ratio (procedure)
C0428613|CACREAT
C0428613|Calcium/Creatinine
C0428613|Calcium/creatinine ratio measurement (procedure)
C0428613|Calcium/creatinine ratio measurement
C1446045|5-Hydroxyindoleacetic acid/creatinine ratio measurement (procedure)
C1446045|5-Hydroxyindoleacetic acid/creatinine ratio measurement
C1446045|5HIAA/creatinine ratio
C1446063|Aminolaevulinic acid / creatinine ratio measurement
C1446063|Aminolaevulinic acid/creatinine ratio measurement
C1446063|Aminolevulinic acid / creatinine ratio measurement
C1446063|Aminolevulinic acid/creatinine ratio measurement (procedure)
C1446063|Aminolevulinic acid/creatinine ratio measurement
C1446063|ALA/creatinine ratio
C1446080|Magnesium to Creatinine Ratio Measurement
C1446080|Magnesium/Creatinine
C1446080|MGCREAT
C1446080|Magnesium / creatinine ratio measurement (procedure)
C1446080|Magnesium / creatinine ratio measurement
C1446080|Magnesium/creatinine ratio
C1446178|Retinol binding protein / creatinine ratio measurement (procedure)
C1446178|Retinol binding protein / creatinine ratio measurement
C1531635|Citrate:creatinine ratio (procedure)
C1531635|Citrate:creatinine ratio
C1531635|Measurement of ratio of citrate to creatinine (procedure)
C1531635|Measurement of ratio of citrate to creatinine
C1531635|Meausrement of ratio of citrate to creatinine
C1531635|Meausrement of ratio of citrate to creatinine (procedure)
C1531635|Citrate/Creatinine
C1531635|Citrate to Creatinine Ratio Measurement
C1531635|Citric Acid/Creatinine
C1531635|CITCREAT
C1559901|CTCAE Grade 1 Creatinine
C1559901|Grade 1 Creatinine
C1559903|CTCAE Grade 3 Creatinine
C1559903|Grade 3 Creatinine
C1559905|CTCAE Grade 5 Creatinine
C1559905|Grade 5 Creatinine
C1559902|CTCAE Grade 2 Creatinine
C1559902|Grade 2 Creatinine
C1559904|CTCAE Grade 4 Creatinine
C1559904|Grade 4 Creatinine
C0852810|Blood creatinine decreased
C0852810|Creatinine blood decreased
C0239150|Creatinine low
C0239150|Creatinine decreased
C3671034|Ascitic fluid creatinine concentration above normal (finding)
C3671034|Ascitic fluid creatitine increased above normal
C3671034|Ascitic fluid creatinine concentration above normal
C0555149|Creatinine in sample (finding)
C0555149|Creatinine in sample
C0600061|Serum creatinine
C0600061|Serum creatinine level
C0600061|Finding of serum creatinine level
C0600061|serum creatinine level finding
C0600061|serum creatinine level finding (lab test)
C0600061|Finding of serum creatinine level (finding)
C0600061|Serum creatinine level - finding
C2114518|previously (less than 3 months) normal creatinine now rising daily
C2114518|previously (less than 3 months) normal creatinine now rising daily (lab test)
C2114518|previously (< 3 months) normal creatinine now rising daily
C2114518|previously (< 3mo.) normal creatinine now rising daily
C2114518|a previously (< 3mo.) normal creatinine is now rising daily
C2097688|serum creatinine was obtained pre-procedure (lab test)
C2097688|serum creatinine was obtained pre-procedure
C2097688|a serum creatinine was obtained pre-procedure
C1278054|Corrected serum creatinine level (procedure)
C1278054|Corrected serum creatinine level
C1278054|Corrected serum creatinine measurement (procedure)
C1278054|Corrected serum creatinine measurement
