C0546647|Iron, total, measurement
C0546647|Iron total
C1446028|serum iron / total iron binding capacity (TIBC) ratio (lab test)
C2229883|serum total iron binding capacity (TIBC)
C0036835|Serum Total Iron-Binding Capacity result
C1277709|iron saturation
C1277709|iron saturation (lab test)
C1277709|Transferrin saturation
C1277709|Transferrin Saturation Measurement
C1277709|Transferrin saturation index (procedure)
C1277709|Transferrin saturation index
C1277709|Saturation of iron binding capacity (procedure)
C1277709|Saturation of iron binding capacity
C1277709|Iron Saturation Percent
C1277709|TFRRNSAT
C1277709|Serum Iron to TIBC Ratio
C1277709|Transferrin Iron Saturation
C1277709|Iron Binding Capacity Saturation
C1277709|Percentage iron saturation
C1277709|Serum transferrin saturation
C0036835|TIBC
C0036835|Serum Total Iron-Binding Capacity result
