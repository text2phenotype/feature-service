C0033707|Protime
C0033707|Prothrombin time
C0033707|Prothrombin time assay
C0151872|Prothrombin time increased
C2346191|CUVETTES,PROTIME DISPOSABLE 3-CHANNEL
C0482694|Coagulation tissue factor induced:Time:Pt:PPP:Qn:Coag
C0482694|Coagulation tissue factor induced
C0482694|Coagulation time
C0482694|LOINC 5902-2
C0482694|LNC 5902-2
C0482694|5902-2
C0482694|Prothrombin time
C0236454|Plasma Control Prothrombin Test
C0236453|Plasma Patient Prothrombin Test
C0033707|Prothrombin Time
C0033707|Prothrombin Times
C0033707|Time, Prothrombin
C0033707|Times, Prothrombin
C0033707|Prothrombin time (PT)
C0033707|PT
C0033707|Prothrombin Time Test
C0033707|prothrombin time (PT) (lab test)
C0033707|Test;prothrombin time
C0033707|Prothrombin time assay
C0033707|PT assay
C0033707|Protime
C0033707|PTT - Prothrombin time
C0033707|Quick one stage prothrombin time
C0033707|PT - Prothrombin time
C0033707|Prothrombin time (procedure)
C0033707|One stage prothrombin time
C0033707|One stage prothrombin time (procedure)
C0033707|Pro-thrombin time
C0033707|Prothrombin test
C0033707|Plasma Prothrombin Test
C1271785|Prothrombin time - reference
C1271785|Prothrombin time - reference (procedure)
C0373814|Prothrombin time; substitution, plasma fractions, each
C0373814|Prothrombin time assay; substitution, plasma fractions, each
C0373814|PROTHROMBIN TIME SUBSTITUTION PLASMA FRCTJ EACH
C0373814|PROTHROMBIN TEST
C4027891|prothrombin time in platelet-poor plasma by coagulation assay
C4027891|prothrombin time (pt) in platelet-poor plasma by coagulation assay
C4027891|prothrombin time in platelet-poor plasma by coagulation assay (lab test)
C4027892|prothrombin time (pt) in capillary blood (lab test)
C4027892|prothrombin time (pt) in capillary blood
C1319577|PT 50:50 mix (procedure)
C1319577|Prothrombin time 50:50 mix (procedure)
C1319577|Prothrombin time 50:50 mix
C1319577|PT 50:50 mix
C1319577|Prothrombin time with 50:50 mix
C1319578|PT 80:20 mix
C1319578|Prothrombin time with 80:20 mix (procedure)
C1319578|Prothrombin time with 80:20 mix
C3853850|International Normalized Ratio of Prothrombin Time
C3853850|Prothrombin Intl. Normalized Ratio
C0151872|Prolonged prothrombin time
C0151872|Prothrombin time inc
C0151872|PT inc
C0151872|Prothrombin level increased
C0151872|Prothrombin time prolonged
C0151872|PT prolonged
C0151872|Prothrombin time increased
C0151872|Coagulation factor II level increased
C0151872|Prothrombin increased
C0151872|PT increased
C0151872|prolonged; prothrombin time
C0151872|prothrombin time; prolonged
C0151872|Prothrombin time increased (finding)
C0151872|Abnormal or prolonged prothrombin time
C0151872|Abnormal or prolonged PT
C3670570|OSPT increased
C3670570|One stage prothrombin time increased
C3670570|One stage prothrombin time increased (finding)
C3670543|Thrombotest prolonged
C3670543|PIVKA test prolonged
C3670543|Thrombotest prolonged (finding)
C2346191|CUVETTES,PROTIME DISPOSABLE 3-CHANNEL
C2346191|CUVETTES,PROTIME DISPOSABLE 3-CHANNEL [VA Product]
C0482694|Coagulation tissue factor induced:Time:Pt:PPP:Qn:Coag
C0482694|Coagulation tissue factor induced:Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay
C0482694|Prothrombin time
C0482694|Prothrombin time (PT)
