C0427512|Finding of white blood cell number
C0023516|Leukocytes
C3842546|Low blood counts, anemia, low white blood cell count, or low platelet count
C0023508|White Blood Cell Count procedure
C0023518|Leukocytosis
C0151370|CSF white count
C0427512|White blood cell count laboratory result
C0438221|White blood cell count normal
C0438223|Differential white count abnormal
C0517645|White blood count depression
C0580531|White blood cell count abnormal
C0750394|White blood cell count decreased
C0750426|White blood cell count increased (lab result)
C1271681|Total white blood count
C1820731|Differential white blood count
C1820736|Absolute white blood count
C1821144|White blood count
C1882326|Percent in White Blood Count Differential
C4055603|APACHE II - White Blood Count
C0162401|Differential white blood cell count procedure
C0427547|Total white cell count measurement
C0438222|Differential white cell count normal
C0855357|Cerebrospinal fluid white blood cell count (lab test)
C0948695|White blood cell count low
C1318024|Total white cell count result
C1820727|Alterations in differential white blood count
C1861189|Increased total white blood count
C2135995|reported abnormal white blood cell count
C2135996|reported high white blood cell count
C2186576|reported white blood cell count
C2186577|reported low white blood cell count
C3495375|Blood count; leukocyte (WBC), automated
C0200629|Complete blood count with white cell differential, manual
C0200630|Complete blood count with white cell differential, automated
C0523122|White blood cell count, automated, cerebrospinal fluid
C0523124|White blood cell count, automated, peritoneal fluid
C0523128|White blood cell count, automated, pleural fluid
C0523133|White blood cell count, automated, semen
C0523135|White blood cell count, automated, synovial fluid
C0855358|CSF white blood cell count negative
C0855359|CSF white blood cell count positive
C0857573|White blood cell count NOS CSF normal
C0857792|White blood cell count NOS CSF abnormal
C0860796|Differential white blood cell count abnormal
C0860797|Differential white blood cell count normal
C0860829|CSF white blood cell count increased
C0860856|White blood cell count semen normal
C0860859|White blood cell count semen high
C1096498|CSF white blood cell count decreased
C1144711|Blood count; automated differential WBC count
C1719330|Other decreased white blood cell count
C1719336|Elevated white blood cell count, unspecified
C1719341|Other elevated white blood cell count
C1719725|Decreased white blood cell count, unspecified
C1822245|Urinary tract infection(<100,000 white blood count)
C2097084|Manual differential white blood cell count
C3516389|Manual white blood cell count and evaluation
C3525567|Buffy coat differential white blood cell count
C3525569|Manual differentiated white blood cell count
C3525788|Manual white blood cell (WBC) count
C3807998|Elevated white cell count in cerebrospinal fluid
C0373807|Leukocyte Alkaline Phosphatase with Count
C0523137|WBC differential count, peripheral blood buffy coat smear
C1303089|Total B lymphocyte count
C1504163|Natural killer (NK) cells, total count
C2676078|WHITE BLOOD CELL COUNT QUANTITATIVE TRAIT LOCUS 1
C3516387|Microscopic examination for white blood cells with manual cell count
C3842546|Low blood counts, anemia, low white blood cell count, or low platelet count
C0523102|Hemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and manual WBC differential
C0523103|Hemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and automated partial WBC differential
C0523104|Hemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and automated complete WBC differential
C1843217|Total white blood cell count less than 25,000/cubic mm with 30-70% eosinophils
C3516392|Automated complete blood cell count
C0151683|Neutrophil count increased
C0151683|Neutrophilia
C0151683|Neutrophils increased
C0151683|Neutrophilia (finding)
C0151683|Granulocytosis
C0151683|Neutrophil count above reference range
C0151683|Neutrophil count high
C0151683|Neutrophilic leukocytosis
C0151683|Neutrophilic leucocytosis
C0001824|Agranulocytoses
C0001824|Agranulocytosis
C0001824|Granulocytopenia
C0001824|Granulocytopenias
C0001824|agranulocytosis (diagnosis)
C0001824|granulocytopenia (diagnosis)
C0001824|Agranulocytosis [Disease/Finding]
C0001824|Agranulocytosis NOS (disorder)
C0001824|Agranulocytosis (finding)
C0001824|Agranulocytosis (disorder)
C0001824|Granulocytopenia (disorder)
C0001824|Granulopenia
C0001824|Agranulocytosis NOS
C0001824|Schultz
C0001824|Granulocytopenic disorder (disorder)
C0001824|Granulocytopenic disorder
C0853697|Peripheral neutropenia
C0853697|Neutropenia
C0853697|Neutrophil count decreased
C0853697|Neutrophils decreased
C0853697|Granulocytopenia
C0853697|Neutrophil count low
C0853697|Neutrophils reduced
C0853697|Neutropenia (finding)
C0853697|Neutrophil count below reference range
C0853986|Decreased lymphocytes
C0853986|Lymphocyte count decreased
C0853986|Lymphocytopenia
C0853986|Lymphocytes decreased below normal range
C0853986|Decreased blood lymphocyte count
C0853986|Lymphopenia
C0853986|Decreased blood lymphocyte count (finding)
C0853986|lymphocytic leukopenia
C0853986|Lymphocyte count low
C0750426|Elevated white blood cell count
C0750426|White blood count elevation
C0750426|White blood cell count increased
C0750426|WBC inc
C0750426|Increased white blood cell count
C0750426|Leukocytosis
C0750426|White blood cell count increased (lab result)
C0750426|White blood cell numbers increased
C0750426|WBC numbers increased
C0750426|Leucocytosis
C0750426|Increased blood leukocyte number
C0750426|Increased blood leucocyte number
C0750426|White blood cell count high
C0750426|White blood cell increased
C0750426|WBC increased
C0750426|Leukocyte count increased
C0750426|Increased white cell count
C0750426|Raised WBC
C0750426|increased; leukocyte count
C0750426|leukocyte count; increased
C0750426|Increased blood leukocyte number (finding)
C0702266|Basophilia
C0702266|basophilia (diagnosis)
C0702266|Basophilia (finding)
C0702266|Circulating basophils increased above normal range
C0702266|Basophilic leukocytosis
C0702266|Basophilic leucocytosis
C0427538|Immature white blood cells NOS (finding)
C0427538|Immature white blood cells (finding)
C0427538|Immature white blood cells NOS
C0427538|Immature white blood cells
C0427548|Relative lymphocytosis
C0427548|Relative lymphocytosis (finding)
C0427549|Reversed differential
C0427549|Reversed differential (finding)
C0750880|Finding of monocyte count
C0750880|Monocyte count result
C0750880|Finding of monocyte count (finding)
C0750880|Monocyte count - finding
C0750880|Monocyte count - observation
C0853698|Lymphocyte count increased
C0853698|Lymphocytes increased above normal range
C0853698|Increased blood lymphocyte number
C0853698|Lymphocytosis
C0853698|Lymphocyte count high
C0853698|Lymphocytes raised
C0853698|Increased blood lymphocyte number (finding)
C0750394|Decreased white blood cell count
C0750394|White blood cell count decreased
C0750394|WBC dec
C0750394|White blood cell numbers decreased
C0750394|WBC numbers decreased
C0750394|leukopenia
C0750394|White blood cell decreased
C0750394|Leucopenia
C0750394|Decreased blood leucocyte number
C0750394|Decreased blood leukocyte number
C0750394|Leukocytopenia
C0750394|Decreased white cell count
C0750394|WBC decreased
C0750394|Leukocyte count decreased
C0750394|Decreased blood leukocyte number (finding)
C2240374|Eosinophil count raised (finding)
C2240374|Eosinophil count increased
C2240374|Eosinophil count raised
C2240374|Eosinophilia
C2240374|Increased blood eosinophil number
C2240374|Increased blood eosinophil number (finding)
C2240374|Increased eosinophils
C2240374|Eosinophilic leukocytosis
C2240374|Eosinophilic leucocytosis
C2240374|Eosinophil count high
C0018183|Granulocyte
C0018183|Granulocytes
C0018183|Granulocytic
C0018183|Granulocytic cells
C0018183|granular leukocyte
C0018183|Granulocytic Cell
C0018183|Granulocyte (cell)
C0018183|Granulocytic cell (cell)
C0018183|Granulocytic cell, NOS
C0018183|Granulocyte (body structure)
C0018183|Granulocytic cell (body structure)
C0018183|Granular Leukocytes
C0022686|K cell
C0022686|killer cell
C0022686|Cytotoxic cell
C0022686|K-cell (cell)
C0022686|K-cell
C0022686|K lymphocyte
C0022686|K lymphocyte (cell)
C0022686|Killer cells
C0022686|K-cell (body structure)
C0024264|Lymphocyte
C0024264|Lymphocytes
C0024264|Lymph Cell
C0024264|Lymphocyte (cell)
C0024264|Lymphocytic cell
C0024264|Lymphocyte, NOS
C0024264|Lymphocytic cell, NOS
C0026473|Monocytes
C0026473|monocyte
C0026473|Blood monocytes
C0026473|Monocyte (cell)
C0026473|Monocyte, NOS
C0031307|Phagocytes
C0031307|phagocyte
C0031307|amebocyte
C0031307|Cell, Phagocytic
C0031307|Cells, Phagocytic
C0031307|Phagocytic Cells
C0031307|Phagocytic Cell
C0031307|Phagocytic cell (cell)
C0031307|Phagocyte, NOS
C0031307|Phagocytic cell, NOS
C0031307|Phagocytic cell (body structure)
C0032112|Plasmacyte
C0032112|Cell, Plasma
C0032112|Cells, Plasma
C0032112|Plasma Cells
C0032112|Plasma Cell
C0032112|plasmocyte
C0032112|plasmacytic
C0032112|Plasma cells.centrocytes
C0032112|Plasma cells.centroblasts
C0032112|Plasmacytes
C0032112|Plasma cell (cell)
C0032112|Plasma cell, NOS
C0032112|Plasma cell (body structure)
C0027950|Leukocyte, Polymorphonuclear
C0027950|Neutrophil
C0027950|Neutrophils
C0027950|Polymorphonuclear Leukocyte
C0027950|Polymorphonuclear cells
C0027950|Neutrophil (cell)
C0027950|Polymorph
C0027950|Polymorphonuclear cells/leukocytes
C0027950|PMN
C0027950|Blood neutrophils
C0027950|Polymorphonuclear Leukocytes
C0027950|Leukocytes, Polymorphonuclear
C0027950|PMN cell
C0027950|Polymorphonuclear leucocyte
C0027950|Polymorphonuclear leukocyte (cell)
C0027950|Neutrophil (body structure)
C0027950|Blood Segmented Neutrophil
C0027950|Neutrophilic Granulocyte
C0027950|Polymorphonuclear Cell
C0027950|Polymorphonuclear Neutrophils
C0027950|Neutrophilic Leukocyte
C0027950|PMN - polymorphonuclear leucocyte
C0027950|PMN - polymorphonuclear leukocyte
C0027950|Polys
C0033416|Promyelocytes
C0033416|Premyelocytes
C0033416|Progranulocytes
C0033416|Promyelocyte
C0033416|Premyelocyte
C0033416|Progranulocyte
C0033416|Promyelocyte (cell)
C0033416|Progranulocyte, NOS
C0033416|Promyelocyte, NOS
C0229635|Metamyelocytes
C0229635|Metamyelocyte
C0229635|Metamyelocyte (cell)
C0369715|Myelocytes
C0369715|myelocyte
C0369715|Myelocyte (cell)
C0023517|Leukocyte, Mononuclear
C0023517|Leukocytes, Mononuclear
C0023517|Mononuclear Leukocyte
C0023517|Nongranular leukocyte
C0023517|agranulocyte
C0023517|Mononuclear Leukocytes
C0023517|Mononucleated Cell
C0023517|Non-Granular Leukocytes
C0023517|Non-Granular Leukocyte
C0368761|Blasts
C0368761|Hematohistioblast
C0368761|Blast cell
C0368761|Ferrata cell
C0368761|Hemocytoblast
C0368761|Haematohistioblast
C0368761|Hemohistioblast
C0368761|Haemocytoblast
C0368761|Polyblast
C0368761|Haemohistioblast
C0368761|blast
C0368761|Blast Cells
C0368761|Blast cell (cell)
C0368761|Blast cell (body structure)
C0023516|Leukocyte
C0023516|WBC
C0023516|Leukocytes
C0023516|Blood Cell, White
C0023516|White Blood Cell
C0023516|Corpuscle, White Blood
C0023516|Blood Corpuscle, White
C0023516|Corpuscles, White Blood
C0023516|White Blood Corpuscle
C0023516|WBC (white blood cell)
C0023516|White blood cell (cell)
C0023516|Leucocytes
C0023516|White blood cells
C0023516|White Blood Corpuscles
C0023516|Blood Corpuscles, White
C0023516|Blood Cells, White
C0023516|Leucocyte
C0023516|WBC - White blood cell
C0023516|Leukocyte (cell)
C0023516|Leukocyte, NOS
C0023516|White blood cell, NOS
C0023516|Reticuloendothelial System, Leukocytes
C0023516|White Cell
C2939172|Lymphocytic (qualifier value)
C2939172|lymphocytic
C0427532|Hypergranular white blood cell
C0427532|Hypergranular white blood cell (cell)
C0427532|Hypergranular white blood cell (body structure)
C0229659|Myelomonocyte
C0229659|Myelomonocyte (cell)
C0229659|Myelomonocyte, NOS
C0229659|Neoplastic Monocyte
C0427534|Agranular white blood cell
C0427534|Agranular white blood cell (cell)
C0427534|Agranular white blood cell (body structure)
C0427533|Hypogranular white blood cell
C0427533|Hypogranular white blood cell (cell)
C0427533|Hypogranular white blood cell (body structure)
C0443777|Neutrophil inclusion
C0443777|Neutrophil inclusion (body structure)
C0443777|Neutrophil inclusion (cell structure)
C0443777|Neutrophil inclusion (cell)
C0427536|White blood cell type (cell)
C0427536|White blood cell type
C0427536|White blood cell type (body structure)
C1268009|Basophilic granulocytic cell (cell)
C1268009|Basophilic granulocytic cell
C1268009|Basophilic granulocytic cell (body structure)
C0229636|Neutrophilic promyelocyte
C0229636|Neutrophilic progranulocyte
C0229636|Neutrophilic promyelocyte (cell)
C1268008|Eosinophilic granulocytic cell (cell)
C1268008|Eosinophilic granulocytic cell
C1268008|Eosinophilic granulocytic cell (body structure)
C1991568|Leukocytes &#x7C; Semen
C1991557|Leukocytes &#124; dialysis fluid peritoneal
C1991557|Leukocytes &#x7C; dialysis fluid peritoneal
C1991567|Leukocytes &#124; peritoneal fluid
C1991567|Leukocytes &#x7C; peritoneal fluid
C1991588|Leukocytes+Platelets &#x7C; Bld-Ser-Plas
C0362942|Leukocytes:NCnc:Pt:Semen:Qn:Manual count
C0362942|Leukocytes [#/volume] in Semen by Manual count
C0362942|WBC # Smn Manual
C0362942|Leukocytes:Number Concentration (count/vol):Point in time:Seminal fluid:Quantitative:Manual count
C1716495|WBC #/area UrnS LPF
C1716495|Leukocytes:Naric:Pt:Urine sed:Qn:Microscopy.light.LPF
C1716495|Leukocytes [#/area] in Urine sediment by Microscopy low power field
C1716495|Leukocytes:Number Aeric (number per area):Point in time:Urine sediment:Quantitative:Microscopy.light.LPF
C1991562|Leukocytes &#x7C; Bone marrow
C2361322|WBC Ur Ql Auto
C2361322|Leukocytes [Presence] in Urine by Automated
C2361322|Leukocytes:ACnc:Pt:Urine:Ord:Automated
C2361322|Leukocytes:Arbitrary Concentration:Point in time:Urine:Ordinal:Automated
C1991558|Leukocytes &#x7C; body fluid
C0362941|WBC # Smn Auto
C0362941|Leukocytes [#/volume] in Semen by Automated count
C0362941|Leukocytes:NCnc:Pt:Semen:Qn:Automated count
C0362941|Leukocytes:Number Concentration (count/vol):Point in time:Seminal fluid:Quantitative:Automated count
C0806987|Mononuclear cells
C1148382|Monocytes+Macrophages
C2361490|Leukocytes.disintegrated
C1114261|Leukocytes [#/volume] in Urine
C1114261|WBC # Ur
C1114261|Leukocytes:NCnc:Pt:Urine:Qn
C1114261|Leukocytes:Number Concentration (count/vol):Point in time:Urine:Quantitative
C2358187|Leukocytes &#x7C; Blood product unit &#x7C; Bld-Ser-Plas
C2358189|Leukocytes &#x7C; Cervix
C1830776|Leukocytes:Number Aeric (number per area):Point in time:Urine sediment:Quantitative:Automated count
C1830776|Leukocytes:Naric:Pt:Urine sed:Qn:Automated count
C1830776|Leukocytes [#/area] in Urine sediment by Automated count
C1830776|WBC #/area UrnS Auto
C1991569|Leukocytes &#124; sputum
C1991569|Leukocytes &#x7C; sputum
C1991574|Leukocytes &#x7C; Vaginal
C1317495|Leukocyte clumps
C1744633|Leukocytes:NCnc:Pt:Urine:Qn:Manual count
C1744633|WBC # Ur Manual
C1744633|Leukocytes [#/volume] in Urine by Manual count
C1744633|Leukocytes:Number Concentration (count/vol):Point in time:Urine:Quantitative:Manual count
C0584614|Finding of large unstained cells
C0584614|Large unstained cells
C0584614|Large unstained cells (qualifier value)
C0584614|Large unstained cells (finding)
C0584614|Finding of large unstained cells (finding)
C3534195|Leukocytes &#x7C; Prostatic fluid
C1991570|Leukocytes &#x7C; stool
C1315523|WBC Ur Ql
C1315523|Leukocytes:ACnc:Pt:Urine:Ord
C1315523|Leukocytes [Presence] in Urine
C1315523|Leukocytes:Arbitrary Concentration:Point in time:Urine:Ordinal
C2970244|Leukocytes:Number = Count/Time:time reported elsewhere:Urine sediment:Quantitative:Microscopy.light
C2970244|WBC ?Tm UrnS Micro-nRate
C2970244|Leukocytes:NRat:XXX:Urine sed:Qn:Microscopy.light
C2970244|Leukocytes by Light microscopy in Urine sediment collected for unspecified duration
C1315296|Leukocytes [Presence] in Semen
C1315296|WBC Smn Ql
C1315296|Leukocytes:ACnc:Pt:Semen:Ord
C1315296|Leukocytes:Arbitrary Concentration:Point in time:Seminal fluid:Ordinal
C0369602|Leukocytes other
C1991551|Leukocytes &#124; bile fluid
C1991551|Leukocytes &#x7C; bile fluid
C1979503|WBC # Ur Auto
C1979503|Leukocytes [#/volume] in Urine by Automated count
C1979503|Leukocytes:NCnc:Pt:Urine:Qn:Automated count
C1979503|Leukocytes:Number Concentration (count/vol):Point in time:Urine:Quantitative:Automated count
C1991566|Leukocytes &#x7C; pleural fluid
C1991564|Leukocytes &#124; pericardial fluid
C1991564|Leukocytes &#x7C; pericardial fluid
C0803223|WBC # Ur Strip
C0803223|Leukocytes:NCnc:Pt:Urine:Qn:Test strip
C0803223|Leukocytes [#/volume] in Urine by Test strip
C0803223|Leukocytes:Number Concentration (count/vol):Point in time:Urine:Quantitative:Test strip
C1991553|Leukocytes &#x7C; blood cord
C1991575|Leukocytes &#x7C; XXX
C1991556|Leukocytes &#x7C; cerebral spinal fluid
C2969596|Leukocytes &#x7C; Blood Product unit.platelet pheresis
C1991552|Leukocytes &#x7C; bld-ser-plas
C0014467|Eosinophil
C0014467|Eosinophils
C0014467|Eosinophil, segmented
C0014467|eosinocyte
C0014467|Blood eosinophils
C0014467|Eosinophil, segmented (cell)
C0014467|Blood Eosinophil
C0014467|Eosinophilic Granulocyte
C0014467|Acidophilic Leukocyte
C0014467|Eosinophilic Leukocyte
C1991563|Leukocytes &#x7C; nose
C3172620|Leukocytes:NRat:24H:Urine sed:Qn:Microscopy
C3172620|Leukocytes in 24 hour Urine sediment by Microscopy
C3172620|Leukocytes:Number = Count/Time:24 hours:Urine sediment:Quantitative:Microscopy
C3172620|WBC 24h UrnS Micro-nRate
C1991571|Leukocytes &#124; synovial fluid
C1991571|Leukocytes &#x7C; synovial fluid
C2358190|Leukocytes &#x7C; Urethra
C3258686|Leukocytes &#x7C; Vitreous fluid
C1991559|Leukocytes &#x7C; gastric fluid
C0485041|Leukocytes [#/volume] in Semen
C0485041|WBC # Smn
C0485041|Leukocytes:NCnc:Pt:Semen:Qn
C0485041|Leukocytes:Number Concentration (count/vol):Point in time:Seminal fluid:Quantitative
C0803269|Leukocytes:ACnc:Pt:Urine sed:Ord:Microscopy.light
C0803269|Leukocytes [Presence] in Urine sediment by Light microscopy
C0803269|WBC UrnS Ql Micro
C0803269|Leukocytes:Arbitrary Concentration:Point in time:Urine sediment:Ordinal:Microscopy.light
C0803389|Leukocytes:NCnc:Pt:XXX:Qn:Automated count
C0803389|Leukocytes [#/volume] in Unspecified specimen by Automated count
C0803389|WBC # XXX Auto
C0803389|Leukocytes:Number Concentration (count/vol):Point in time:To be specified in another part of the message:Quantitative:Automated count
C0801449|Leukocytes:NRat:12H:Urine sed:Qn:Microscopy.light
C0801449|Leukocytes in 12 hour Urine sediment by Light microscopy
C0801449|Leukocytes:Number = Count/Time:12 hours:Urine sediment:Quantitative:Microscopy.light
C0801449|WBC 12h UrnS Micro-nRate
C0368036|Leukocytes:Naric:Pt:Urine sed:Qn:Microscopy.light.HPF
C0368036|Leukocytes [#/area] in Urine sediment by Microscopy high power field
C0368036|WBC #/area UrnS HPF
C0368036|Leukocytes:Number Aeric (number per area):Point in time:Urine sediment:Quantitative:Microscopy.light.HPF
C2924077|Leukocytes in 3 hour Urine sediment by Light microscopy
C2924077|Leukocytes:NRat:3H:Urine sed:Qn:Microscopy.light
C2924077|Leukocytes:Number = Count/Time:3 hours:Urine sediment:Quantitative:Microscopy.light
C2924077|WBC 3h UrnS Micro-nRate
C3484293|Basophils+Mast cells
C2598498|Leukocytes:ACnc:Pt:Urine:Ord:Visual
C2598498|Leukocytes [Presence] in Urine by Visual
C2598498|WBC Ur Ql Visual
C2598498|Leukocytes:Arbitrary Concentration:Point in time:Urine:Ordinal:Visual
C2356936|Basophils+Eosinophils+Monocytes &#x7C; Bld-Ser-Plas
C2358264|Lymphocytes+Monocytes &#x7C; Bld-Ser-Plas
C2969597|Leukocytes &#x7C; fetus
C1991555|Leukocytes &#x7C; bronchial
C2588282|Leukocytes &#x7C; Dialysis fluid
C3172621|Leukocytes:NCnc:XXX:Urine sed:Qn:Microscopy.light.HPF
C3172621|Leukocytes:Number Concentration (count/vol):time reported elsewhere:Urine sediment:Quantitative:Microscopy.light.HPF
C3172621|WBC ?Tm # UrnS HPF
C3172621|Leukocytes [#/volume] by Microscopy high power field in Urine sediment collected for unspecified duration
C3480571|Ragocytes &#x7C; Synovial fluid
C2923139|Leukocytes:NCnc:Pt:Urine:Qn:Test strip.automated
C2923139|Leukocytes [#/volume] in Urine by Automated test strip
C2923139|WBC # Ur Strip.auto
C2923139|Leukocytes:Number Concentration (count/vol):Point in time:Urine:Quantitative:Test strip.automated
C1991576|Leukocytes left shift &#x7C; bld-ser-plas
C0023172|Cell, LE
C0023172|Cells, LE
C0023172|LE Cell
C0023172|LE cell (cell)
C0023172|Lupus erythematosus (LE) cell
C0023172|Lupus erythematosus cells
C0023172|Lupus erythematosus cell
C0023172|Lupus erythematosus cell (cell)
C0023172|Lupus erythematosus (LE) cell (cell)
C0023172|L.E. cells
C0023172|L.E. cell
C0023172|Lupus erythematosus cell (morphologic abnormality)
C0023172|LE cell (body structure)
C0023172|LE Cells
C0312740|effector cell
C0312740|Effector Immune Cell
C0312740|Immune effector cell
C0312740|Immune effector cell (cell)
C0312740|Immune effector cell (body structure)
C1321301|Peripheral blood mononuclear cell (cell)
C1321301|Peripheral Blood Mononuclear Cells [Chemical/Ingredient]
C1321301|Peripheral Blood Mononuclear Cells
C1321301|PERIPHERAL BLOOD MONONUCLEAR CELL
C1321301|PBMC
C0022688|Cell, Natural Killer
C0022688|Cell, NK
C0022688|Cells, Natural Killer
C0022688|Cells, NK
C0022688|Killer Cell, Natural
C0022688|Killer Cells, Natural
C0022688|Natural Killer Cell
C0022688|NK Cell
C0022688|K lymphocyte
C0022688|Killer cell
C0022688|K cell
C0022688|NK-cell (cell)
C0022688|Natural killer (NK)-cell
C0022688|Natural killer cell (cell)
C0022688|Natural killer (NK)-cell (cell)
C0022688|NK-LGL
C0022688|NK (natural killer) cell
C0022688|Natural Killer Cells
C0022688|NK Cells
C0022688|NK-cell
C0022688|NK-cell (body structure)
C0022688|Killer Cells
C0022688|NK
C0064828|leucoagglutinins, leukocyte
C0064828|leukoagglutinins, leukocytes
C1518997|PBL
C1518997|Peripheral Blood Lymphocyte
C0004827|Basophil
C0004827|Basophils
C0004827|Basophil, segmented
C0004827|Basophil, segmented (cell)
C0004827|Basophilic Leukocyte
C0004827|Basophilic Granulocyte
C0236610|Whole Blood Band Form Leukocyte Counts
C0236601|Whole Blood Basophil Counts
C0236606|Whole Blood Blast Cell Counts
C0236602|Whole Blood Eosinophil Counts
C1254474|Whole Blood Hypersegmented Neutrophil Test
C0236609|Whole Blood Metamyelocyte Counts
C1254716|Whole Blood Mononucleated Cell Count
C0236608|Whole Blood Myelocyte Counts
C1254593|Whole Blood Myeloid Precursor Counts
C0236611|Whole Blood Neutrophil Counts
C0236600|Whole Blood Plasma Cell Counts
C1255495|Whole Blood Prolymphocyte Counts
C1255496|Whole Blood Promonocyte Counts
C0236607|Whole Blood Promyelocyte Counts
C1254480|Whole Blood Total Leukocyte Count
C0200635|Lymphocyte count
C0200635|Lymphocyte Count, Total
C0200635|Lymphocyte Counts
C0200635|Lymphocyte Counts, Total
C0200635|Total Lymphocyte Counts
C0200635|Lymphocyte Count measurement
C0200635|blood lymphocyte count
C0200635|blood lymphocyte count (lab test)
C0200635|Total lymphocyte count (procedure)
C0200635|Total lymphocyte count
C0200635|Lymphocyte count NOS
C0200635|Lymphocyte count (procedure)
C0200635|Lymphocyte count NOS (procedure)
C0200635|LYM
C0200635|Lymphocytes
C0200635|Lymphocyte Number
C0200635|Lymphocyte Numbers
C0023508|White Blood Cell Count
C0023508|Count, Leukocyte
C0023508|Counts, Leukocyte
C0023508|Leukocyte Count
C0023508|Leukocyte Counts
C0023508|Leukocyte Numbers
C0023508|Number, Leukocyte
C0023508|Numbers, Leukocyte
C0023508|White Blood Cell Count procedure
C0023508|leukocyte count (lab test)
C0023508|WBC count
C0023508|White blood cell count (procedure)
C0023508|Leukocytes
C0023508|White Blood Cells
C0023508|WBC
C0023508|White cells
C0023508|Leukocyte count NOS
C0023508|White blood cell count NOS
C0023508|White blood cell analysis
C0023508|Leucocyte count
C0023508|Leukocyte Number
C0023508|Blood Cell Count, White
C0023508|Whole Blood Leukocyte Counts
C0023508|WBC - White blood cell count
C0023508|WCC - White blood cell count
C0023508|White blood cell count - observation
C1883362|Total Basophil Count
C1883362|Basophils
C1883362|BASO
C0200638|Eosinophil count
C0200638|blood eosinophil count (lab test)
C0200638|blood eosinophil count
C0200638|Eosinophil count procedure
C0200638|Eosinophil count NOS
C0200638|Eosinophil count NOS (procedure)
C0200638|Eosinophils
C0200638|EOS
C0200638|Eosinophil count (procedure)
C0200638|Eosinophil count - observation
C0200637|Monocyte count
C0200637|blood monocyte count (lab test)
C0200637|blood monocyte count
C0200637|Monocyte count procedure
C0200637|Monocyte count (procedure)
C0200637|Monocyte count NOS (procedure)
C0200637|Monocyte count NOS
C0200637|MONO
C0200637|Monocytes
C0455285|Metamyelocyte count
C0455285|Metamyelocyte count procedure
C0455285|Metamyelocyte count (procedure)
C0455285|Metamyelocytes
C0455285|METAMY
C0455285|Metamyelocyte count procedure (procedure)
C2698887|Promonocyte Count
C2698887|Promonocytes
C2698887|PROMONO
C0455279|Promyelocyte count
C0455279|Promyelocyte count procedure
C0455279|Promyelocyte count (procedure)
C0455279|Promyelocytes
C0455279|PROMY
C0455279|Promyelocyte count procedure (procedure)
C2699318|Smudge Cell Count
C2699318|Basket Cells
C2699318|SMDGCE
C2699318|Smudge Cells
C2699318|Gumprecht Shadow Cells
C2699318|Shadow Cells
C0455284|Myelocyte count
C0455284|Myelocyte count procedure
C0455284|Myelocyte count (procedure)
C0455284|Myelocytes
C0455284|MYCY
C0455284|Myelocyte count procedure (procedure)
C2238207|neutrophils
C2238207|neutrophils as percentage of blood leukocytes (lab test)
C2238207|neutrophils as percentage of blood leukocytes
C2238207|WBC count - neutrophil % (lab test)
C2238207|WBC count - neutrophil %
C2109247|juvenile and band neutrophils as percentage of blood leukocytes (lab test)
C2109247|juvenile and band neutrophils as percentage of blood leukocytes
C2109247|juvenile and band neutrophils
C2228144|eosinophils as percentage of blood leukocytes (lab test)
C2228144|eosinophils as percentage of blood leukocytes
C2228144|eosinophils
C2237945|basophils as percentage of blood leukocytes (lab test)
C2237945|basophils as percentage of blood leukocytes
C2237945|basophils
C2200256|lymphocytes as percentage of blood leukocytes (lab test)
C2200256|lymphocytes as percentage of blood leukocytes
C2200256|lymphocytes
C2238069|blood lymphocyte count by Coulter
C2238069|blood lymphocyte count by Coulter (lab test)
C2238069|blood lymphocyte count (Coulter)
C2238069|lymphocytes (Coulter)
C0427546|leukocyte count atypical lymphocytes
C0427546|leukocyte count atypical lymphocytes (lab test)
C0427546|atypical lymphocytes
C0427546|Atypical lymphocyte observed
C0427546|Abnormal;lymphocytes
C0427546|Abnormal lymphocytes
C0427546|Abnormality of lymphocytes
C0427546|Lymphocyte abnormal
C0427546|Lymphocyte abnormality
C0427546|Lymphocyte abnormality (finding)
C2237144|monocytes as percentage of blood leukocytes
C2237144|monocytes as percentage of blood leukocytes (lab test)
C2237144|monocytes
C0948762|Absolute neutrophil count
C0948762|ANC
C0948762|blood absolute neutrophil count (ANC)
C0948762|blood absolute neutrophil count (ANC) (lab test)
C0948762|blood ANC
C0948762|blood absolute neutrophil count
C0948762|blood absolute granulocyte count
C0948762|blood ANC (absolute neutrophil count)
C0948762|blood absolute neutrophil count (lab test)
C0948762|Neutrophils
C0948762|NEUT
C0200633|Neutrophil count
C0200633|seg (blood count)
C0200633|poly count
C0200633|blood neutrophil count (lab test)
C0200633|blood neutrophil count
C0200633|Neutrophil count (procedure)
C0200633|Neutrophil count NOS (procedure)
C0200633|Neutrophil count NOS
C0200633|Neutrophil count [dup] (procedure)
C0200641|Basophil count
C0200641|blood basophil count
C0200641|blood basophil count (lab test)
C0200641|Basophil count NOS (procedure)
C0200641|Basophil count NOS
C0200641|Basophil count (procedure)
C0200641|Basophils
C0200641|Basophil count [dup] (procedure)
C1144711|automated differential WBC count
C1144711|white blood cell count with automated differential (lab test)
C1144711|WBC count with automated diff
C1144711|white blood cell count with automated differential
C1144711|automated white blood cell differential
C1144711|WBC count with automated differential
C1144711|BLOOD COUNT AUTOMATED DIFFERENTIAL WBC COUNT
C1144711|Automated differential white blood cell count
C1144711|Automated differential leukocyte (WBC) count
C1144711|Blood count; automated differential WBC count
C1144711|AUTOMATED DIFF WBC COUNT
C0523113|blood blast count
C0523113|blood blast count (lab test)
C0523113|Blast Count
C0523113|BLAST
C0523113|Blasts
C0523113|Blast cells
C0523113|Blast cells NOS
C0523113|Blast count, blood
C0523113|Blast count, blood (procedure)
C0523113|Blast count procedure
C2208800|blood granulocytes count
C2208800|blood granulocytes count (lab test)
C2097084|WBC count with manual diff
C2097084|white blood cell count with manual differential
C2097084|white blood cell count with manual differential (lab test)
C2097084|WBC count with manual differential
C2097084|Manual differential white blood cell count
C0857490|Granulocyte count
C0857490|Granulocytes
C0857490|GRAN
C0857490|Granulocyte count (procedure)
C3272948|Immature Basophil Count
C3272948|Immature Basophils
C3272948|BASOIM
C3272953|Immature Granulocyte Count
C3272953|Immature Granulocytes
C3272953|GRANIM
C0162401|Count, Differential Leukocyte
C0162401|Counts, Differential Leukocyte
C0162401|Differential Leukocyte Counts
C0162401|Leukocyte Counts, Differential
C0162401|Differential white blood cell count
C0162401|Differential Leukocyte Count
C0162401|Diff. white cell count NOS (procedure)
C0162401|Diff. white cell count NOS
C0162401|Differential white blood cell count (procedure)
C0162401|Differential WBC count
C0162401|Differential white blood cell count procedure (procedure)
C0162401|Differential white blood cell count procedure
C0162401|Leukocyte Count, Differential
C0236603|Whole Blood Monocyte Counts
C0236604|Whole Blood Atypical Lymphocyte Counts
C0236605|Whole Blood Lymphocyte Counts
C0373752|BLOOD COUNT SMEAR MCRSCP W/MNL DIFRNTL WBC COUNT
C0373752|Blood count; blood smear, microscopic examination with manual differential WBC count
C0373752|BL SMEAR W/DIFF WBC COUNT
C0373754|BLOOD COUNT MANUAL DIFRNTL WBC COUNT BUFFY COAT
C0373754|Manual differential leukocyte (WBC) count on buffy coat
C0373754|Blood count; manual differential WBC count, buffy coat
C0373754|MANUAL DIFF WBC COUNT B-COAT
C3495375|BLOOD COUNT LEUKOCYTE WBC AUTOMATED
C3495375|Automated white blood cell count
C3495375|Automated white blood cell (WBC) count
C3495375|Blood count; leukocyte (WBC), automated
C3495375|AUTOMATED LEUKOCYTE COUNT
C0427547|Total white cell count NOS
C0427547|Total white cell count NOS (procedure)
C0427547|Total white cell count measurement
C3890712|Heterophils
C3890712|Heterophil Measurement
C3890712|HETRPH
C4028024|peritoneal lavage wbc count
C4028024|peritoneal lavage wbc count (procedure)
C4064392|other leukocytes % (lab test)
C4064392|other leukocytes %
C4064392|wbc count - other leukocytes %
C1294061|Leucocyte count corrected for nucleated erythrocytes
C1294061|Leukocyte count corrected for nucleated erythrocytes (procedure)
C1294061|Leukocyte count corrected for nucleated erythrocytes
C1294062|Mononuclear cell count
C1294062|Agranulocyte count
C1294062|Mononuclear cell count (procedure)
C0580952|Myeloblast count
C0580952|Myeloblast count procedure
C0580952|Myeloblast count (procedure)
C0580952|Myeloblasts
C0580952|MYBLA
C0580952|Myeloblast count procedure (procedure)
C0427550|Reversed neutrophil/lymphocyte ratio
C0427550|Reversed neutrophil/lymphocyte ratio measurement (procedure)
C0427550|Reversed neutrophil/lymphocyte ratio measurement
C1271682|Total WBC (IMM) (procedure)
C1271682|Total WBC (IMM)
C1271681|Total white blood cell count (procedure)
C1271681|Total white blood count (procedure)
C1271681|Total white blood cell count
C1271681|Total white blood count
C0024282|Lymphocytoses
C0024282|Lymphocytosis
C0024282|lymphocytosis (diagnosis)
C0024282|Lymphocytosis [Disease/Finding]
C0024282|Disorder characterized by lymphocytosis
C0024282|Lymphocytosis (disorder)
C0024282|Lymphocytosis, NOS
C0543669|NEUTROPHILIA, HEREDITARY
C0543669|neutrophilia hereditary
C0543669|Hereditary neutrophilia (diagnosis)
C0543669|Hereditary neutrophilia
C0543669|Hereditary neutrophilia (disorder)
C0543669|Hereditary neutrophilia (finding)
C0023501|Leukemoid Reaction
C0023501|Leukemoid Reactions
C0023501|Reactions, Leukemoid
C0023501|Reaction, Leukemoid
C0023501|Leukaemoid reaction
C0023501|leukemoid reaction (diagnosis)
C0023501|Leukemoid reaction NOS
C0023501|Leukemoid Reaction [Disease/Finding]
C0023501|Reaction leukemoid
C0023501|Leukemoid reaction (disorder)
C0023501|leukemoid; reaction
C0023501|reaction; leukemoid
C0023501|Leukemoid reaction, NOS
C0023518|Leukocytoses
C0023518|Leukocytosis
C0023518|Leukocytosis, unspecified
C0023518|leukocytosis (diagnosis)
C0023518|Leukocytosis NOS
C0023518|Leukocytosis [Disease/Finding]
C0023518|Leucocytosis
C0023518|Leucocytosis (finding)
C0023518|Disorder characterized by leukocytosis
C0023518|Leucocytosis NOS
C0023518|Leukocytosis (disorder)
C0023518|Leucocytosis, NOS
C0023518|Leukocytosis, NOS
C0741439|Bandemia
C0741439|bandemia (diagnosis)
C0741439|Band neutrophil count above reference range (finding)
C0741439|Band neutrophil count above reference range
C0741439|Bandaemia
C2118400|leukocytosis secondary to steroids (diagnosis)
C2118400|leukocytosis secondary to steroids
C1853187|HOLOPROSENCEPHALY, RECURRENT INFECTIONS, AND MONOCYTOSIS
C0151857|Pleocytosis
C0151857|Pleocytosis of cerebrospinal fluid
C0151857|Pleocytoses
C0151857|Pleocytosis of CSF
C0151857|CSF pleocytosis
C0151857|Cerebrospinal fluid pleocytosis
C0151857|Pleocytosis of cerebrospinal fluid (finding)
C0398571|Other specified other white blood cell disease
C0398571|Other specified other white blood cell disease (disorder)
C3665444|Neutrophilia
C3665444|neutrophilia (diagnosis)
C3665444|Neutrophilic leukocytosis
C3665444|Neutrophilia (finding)
C3665444|Neutrophilia (disorder)
C3665444|Neutrocytosis
C3665444|Neutrophilia, NOS
C3665444|Neutrophilia (disorder) [Ambiguous]
C3665444|Nnutrophilia
C0494244|Other disorders of white blood cells
C0494244|Other white blood cell disease (disorder)
C0494244|Other white blood cell disease
C0494244|Other white blood cell disease NOS
C0494244|Other white blood cell disease NOS (disorder)
C0856808|Polymorphonuclear leucocytosis
C0856808|Polymorphonuclear leukocytosis
C3686749|Stress leukogram
C3686749|Physiologic leukocytosis (disorder)
C3686749|Physiologic leukocytosis
C3686749|Stress hemogram
C0014457|Eosinophilia
C0014457|Eosinophilias
C0014457|eosinophilic leukocytosis (diagnosis)
C0014457|eosinophilia (diagnosis)
C0014457|eosinophilic leukocytosis
C0014457|Eosinophilia [Disease/Finding]
C0014457|Eosinophilia NOS
C0014457|Eosinophilic leucocytosis
C0014457|Eosinophilia (disorder)
C0014457|Eosinophilia NOS (disorder)
C0014457|Eosinophilia, NOS
C0014457|Eosinophilia (disorder) [Ambiguous]
C0272164|Leukoerythroblastotic reaction
C0272164|Leukoerythroblastotic reaction (disorder)
C0398664|Post-splenectomy leucocytosis
C0398664|Post-splenectomy leukocytosis (disorder)
C0398664|Post-splenectomy leukocytosis
C0085702|Monocytosis
C0085702|monocytosis (diagnosis)
C0085702|Disorder characterized by monocytosis
C0085702|Monocytosis (disorder)
C0085702|Monocytosis, NOS
C0085077|Sweets Syndrome
C0085077|Syndrome, Sweet's
C0085077|Acute febrile neutrophilic dermatosis
C0085077|Febrile neutrophilic dermatosis [Sweet]
C0085077|NEUTROPHILIC DERMATOSIS, ACUTE FEBRILE
C0085077|SS
C0085077|Sweet's syndrome
C0085077|Sweet's syndrome (diagnosis)
C0085077|Syndrome, Sweet
C0085077|Sweet Syndrome
C0085077|Dermatosis, Neutrophilic, Febrile, Acute
C0085077|Sweet Syndrome [Disease/Finding]
C0085077|Disease, Gomm-Button
C0085077|Gomm-Button Disease
C0085077|Disease, Gomm Button
C0085077|Gomm Button Disease
C0085077|AFND
C0085077|Sweet disease
C0085077|Sweet's disease
C0085077|Febrile neutrophilic dermatosis
C0085077|Acute febrile neutrophilic dermatosis (disorder)
C0085077|dermatosis; febrile neutrophilic
C0085077|Sweet
C0085077|febrile neutrophilic; dermatosis
C0438221|White blood cell count normal
C0438221|White cell count normal (finding)
C0438221|White cell count normal
C0438221|Leucocyte count normal
C0438221|Leukocyte count normal
C0438221|White blood cell count normal (finding)
C0438222|Diff. white cell count normal
C0438222|Differential white cell count normal
C0438222|Diff. white cell count normal (finding)
C0438222|Differential white cell count normal (finding)
C0427542|Monocyte count normal
C0427542|Monocyte count normal (finding)
C0438223|Diff. white count abnormal
C0438223|Differential white count abnormal
C0438223|Diff. white count abnormal (finding)
C0438223|Differential white count abnormal (finding)
C0580531|White cell count abnormal
C0580531|White cell count abnormal (finding)
C0580531|Abnormal leukocyte count
C0580531|White blood cell count abnormal NOS
C0580531|White blood cell count abnormal
C0580531|Leucocyte count abnormal
C0580531|Leukocyte count abnormal
C0580531|White blood cell count abnormal (finding)
C0580319|Monocytes.abnormal
C0580319|Monocyte count abnormal
C0580319|Abnormal monocytes (finding)
C0580319|Monocyte count abnormal (finding)
C0580319|Abnormal monocytes
C0580319|Abnormal monocyte count
C0580319|Monocyte count abnormal NOS
C0580319|Monocytes abnormal
C0580550|Lymphocyte count abnormal
C0580550|Lymphocyte count abnormal (finding)
C0580550|Abnormal lymphocyte count
C0580550|Abnormal number of lymphocytes
C0580550|Abnormality of lymphocyte number
C0580550|Lymphocyte count abnormal NOS
C0580550|Abnormal lymphocyte counts
C0580550|Abnormal numbers of lymphocytes
C0023530|Leukopenia
C0023530|Leukopenias
C0023530|Leukocytopenias
C0023530|Leukopenia NOS
C0023530|Leukocytopenia, unspecified
C0023530|leukopenia (diagnosis)
C0023530|Leucopenia, NOS
C0023530|Leukopenia, NOS
C0023530|Leucocytopenia
C0023530|Leukocytopenia NOS
C0023530|Leukocytopenia
C0023530|Leukopenia [Disease/Finding]
C0023530|Leucopenia
C0023530|Leucopenia (finding)
C0023530|Leucopenia (disorder)
C0023530|Disorder characterized by neutropenia
C0023530|Leukopenia (disorder)
C0151787|Myeloid maturation arrest
C0151787|Maturation arrest myeloid
C0151787|Arrest myeloid maturation
C0024312|Lymphocytopenias
C0024312|Lymphopenia
C0024312|Lymphopenias
C0024312|Lymphocytopenia
C0024312|lymphopenia (diagnosis)
C0024312|lymphocytopenia (diagnosis)
C0024312|Decreased lymphocytes
C0024312|Lymphopenia [Disease/Finding]
C0024312|Disorder characterized by lymphopenia
C0024312|Lymphocytopenia (disorder)
C0024312|Lymphocytopenia, NOS
C1719330|Other decreased white blood cell count
C1719330|Decreased WBC count NEC
C1719725|Decreased white blood cell count, unspecified
C3687167|Decreased blood basophil number (finding)
C3687167|Decreased blood basophil number
C3670590|Leukopenia with degenerative left shift (finding)
C3670590|Leukopenia with degenerative left shift
C3687166|Decreased blood heterophil count
C3687166|Decreased blood heterophil count (finding)
C0427544|Monocytopenia
C0427544|monocytopenia (diagnosis)
C0427544|Monocytopenia (finding)
C1689996|Decreased eosinophils
C1689996|Eosinopenia
C1689996|Decreased blood eosinophil number
C1689996|Decreased blood eosinophil number (finding)
C1719331|Basophilic leukopenia
C1719331|basopenia (diagnosis)
C1719331|basopenia
C1719331|decreased basophils
C1719337|Lymphocytosis (symptomatic)
C1719337|Lymphocytosis-symptomatc
C1719340|Monocytosis (symptomatic)
C1719340|Monocytosis-symptomatic
C0085663|Plasmacytosis
C0085663|plasmacytosis (diagnosis)
C0085663|Plasmacytosis (disorder)
C0085663|Plasmocytosis
C0085663|Plasmacytosis, NOS
C1719341|Other elevated white blood cell count
C1719341|Elevated WBC count NEC
C1719336|Elevated white blood cell count, unspecified
C3686643|Increased blood heterophil number
C3686643|Increased blood heterophil number (finding)
C3686643|Heterophilia
C0427543|Monocyte count raised (finding)
C0427543|Monocyte count raised
C0427543|Monocytes increased above normal range
C0427543|Monocytosis
C0427543|Increased blood monocyte number
C0427543|Increased blood monocyte number (finding)
C0579194|Percentage differential white blood cells
C0579194|Determination of percentage differential white blood cells (procedure)
C0579194|Determination of percentage differential white blood cells
C0855357|cerebrospinal fluid leukocytes (lab test)
C0855357|cerebrospinal fluid leukocytes
C0855357|CSF cells WBC
C0855357|cerebrospinal fluid cells leukocyte
C0855357|CSF WBC cells
C0855357|CSF WBC
C0855357|Cerebrospinal fluid white blood cell count (lab test)
C0855357|CSF white blood cell count
C0855357|Cerebrospinal fluid white blood cell count NOS
C0855357|White blood cell count NOS cerebrospinal fluid
C0855357|Cerebrospinal fluid white cell count NOS
C0855357|CSF white cell count NOS
C0855357|CSF white blood cell count NOS
C0855357|Cerebrospinal fluid WBC
C0855357|White blood cell count NOS CSF
C0855357|Cerebrospinal fluid white blood cell count
C2026628|cerebrospinal fluid lymphocytes and monocytes as percentage of leukocytes
C2026628|CSF cells WBC % lymphocytes + monocyte
C2026628|cerebrospinal fluid lymphocytes and monocytes as percentage of leukocytes (lab test)
C2026628|cerebrospinal fluid cells leukocyte % lymphocytes + monocyte
C2026628|CSF lymphocytes and monocytes as percentage of leukocytes
C2026641|cerebrospinal fluid neutrophils as percentage of leukocytes
C2026641|CSF cells WBC % neutrophils
C2026641|cerebrospinal fluid neutrophils as percentage of leukocytes (lab test)
C2026641|cerebrospinal fluid cells leukocyte % neutrophils
C2026641|CSF neutrophils as percentage of leukocytes
C2026590|cerebrospinal fluid eosinophils as percentage of leukocytes (lab test)
C2026590|CSF cells WBC eosinophils
C2026590|cerebrospinal fluid cells leukocyte eosinophils
C2026590|cerebrospinal fluid eosinophils as percentage of leukocytes
C2026590|CSF eosinophils as percentage of leukocytes
C2026529|cerebrospinal fluid cells leukocyte % basophils
C2026529|cerebrospinal fluid basophils as percentage of leukocytes (lab test)
C2026529|CSF cells WBC % basophils
C2026529|cerebrospinal fluid basophils as percentage of leukocytes
C2026529|CSF basophils as percentage of leukocytes
C2026535|cerebrospinal fluid cells immature neutrophils bands (lab test)
C2026535|CSF cells WBC immature neutrophils (bands)
C2026535|cerebrospinal fluid cells immature neutrophils bands
C2026535|CSF cells immature neutrophils bands
C0523122|csf cells wbc automated count
C0523122|CSF WBC, automated count
C0523122|CSF WBC, automated count (lab test)
C0523122|White blood cell count, automated, cerebrospinal fluid
C0523122|White blood cell count, automated, cerebrospinal fluid (procedure)
C4065692|csf cells wbc manual count
C4065692|CSF WBC, manual count
C4065692|CSF WBC, manual count (lab test)
C0948695|White blood cell count low
C2135995|WBC count was abnormal
C2135995|reported abnormal white blood cell count
C2135995|reported abnormal white blood cell count (history)
C2135995|reported abnormal white cell count
C2135996|reported high white blood cell count (history)
C2135996|reported high white blood cell count
C2135996|reported high white cell count
C2186577|reported low white cell count
C2186577|reported low white blood cell count
C2186577|reported low white blood cell count (history)
C4029833|cbc with manual differential reflex
C4029833|CBC with reflex manual differential
C4029833|CBC with reflex manual differential (lab test)
C0523102|Hemogram, automated, with RBC, WBC, Hgb, Hct, indices, platelet count, and manual WBC differential
C0523102|Hemogram, automated, with red blood cells, white blood cells, hemoglobin, hematocrit, indices, platelet count, and manual white blood cell differential
C0523102|Hemogram, automated, with red blood cells, white blood cells, hemoglobin, hematocrit, indices, platelet count, and manual white blood cell differential (procedure)
C0523102|Hemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and manual WBC differential (procedure)
C0523102|Haemogram, automated, with red blood cells, white blood cells, haemoglobin, haematocrit, indices, platelet count, and manual white blood cell differential
C0523102|Haemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and manual WBC differential
C0200629|complete blood count with manual differential
C0200629|complete blood count with manual differential (lab test)
C0200629|CBC with manual differential
C0200629|Complete blood count with white cell differential, manual
C0200629|Complete blood count with white cell differential, manual (procedure)
C0200630|CBC with automated differential
C0200630|CBC with automated differential (lab test)
C0200630|Complete blood count with white cell differential, automated
C0200630|Complete blood count with white cell differential, automated (procedure)
C0523104|Hemogram, automated, with RBC, WBC, Hgb, Hct, indices, platelet count, and automated complete WBC differential
C0523104|Hemogram, automated, with red blood cells, white blood cells, hemoglobin, hematocrit, Indices, Platelet count, and automated complete white blood cell differential (procedure)
C0523104|Hemogram, automated, with red blood cells, white blood cells, hemoglobin, hematocrit, Indices, Platelet count, and automated complete white blood cell differential
C0523104|Hemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and automated complete WBC differential (procedure)
C0523104|Haemogram, automated, with red blood cells, white blood cells, haemoglobin, haematocrit, Indices, Platelet count, and automated complete white blood cell differential
C0523104|Haemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and automated complete WBC differential
C0523103|Hemogram, automated, with RBC, WBC, Hgb, Hct, indices, platelet count, and automated partial WBC differential
C0523103|Hemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and automated partial WBC differential (procedure)
C0523103|Hemogram, automated, with red blood cell, white blood cell, hemoglobin, hematocrit, Indices, Platelet count, and automated partial white blood cell differential
C0523103|Hemogram, automated, with red blood cell, white blood cell, hemoglobin, hematocrit, Indices, Platelet count, and automated partial white blood cell differential (procedure)
C0523103|Hemogram, automated, with red blood cell, white blood cell, hemoglobin, hemtocrit, Indices, Platelet count, and automated partial white blood cell differential (procedure)
C0523103|Hemogram, automated, with red blood cell, white blood cell, hemoglobin, hemtocrit, Indices, Platelet count, and automated partial white blood cell differential
C0523103|Haemogram, automated, with red blood cell, white blood cell, haemoglobin, haematocrit, Indices, Platelet count, and automated partial white blood cell differential
C0523103|Haemogram, automated, with RBC, WBC, Hgb, Hct, Indices, Platelet count, and automated partial WBC differential
C0855358|White blood cell count NOS CSF negative
C0855358|CSF WBC negative
C0855358|Cerebrospinal fluid white blood cell count NOS negative
C0855358|White blood cell count NOS cerebrospinal fluid negative
C0855358|CSF white blood cell count NOS negative
C0855358|CSF white blood cell count negative
C0855358|Cerebrospinal fluid WBC negative
C0855358|Cerebrospinal fluid white blood cell count negative
C0855359|Cerebrospinal fluid WBC positive
C0855359|CSF white blood cell count NOS positive
C0855359|Cerebrospinal fluid white blood cell count NOS positive
C0855359|White blood cell count NOS CSF positive
C0855359|CSF white blood cell count positive
C0855359|White blood cell count NOS cerebrospinal fluid positive
C0855359|CSF WBC positive
C0855359|Cerebrospinal fluid white blood cell count positive
C0857573|CSF white cell count NOS normal
C0857573|Cerebrospinal fluid white blood cell count NOS normal
C0857573|White blood cell count NOS CSF normal
C0857573|Cerebrospinal fluid white cell count NOS normal
C0857573|CSF white blood cell count NOS normal
C0857573|White blood cell count NOS cerebrospinal fluid normal
C0857792|Cerebrospinal fluid white blood cell count NOS abnormal
C0857792|Cerebrospinal fluid white cell count NOS abnormal
C0857792|White blood cell count NOS CSF abnormal
C0857792|CSF white blood cell count NOS abnormal
C0857792|CSF white cell count NOS abnormal
C0857792|White blood cell count NOS cerebrospinal fluid abnormal
C0860796|Differential white blood cell count abnormal
C0860796|Differential white blood cell count abnormal NOS
C0860796|WBC classification abnormal
C0860796|Differential WBC count abnormal
C0860796|leukocyte count differential abnormal
C0860797|Differential white blood cell count normal
C0860797|Differential WBC count normal
C0860829|CSF white blood cell count increased
C0860829|White blood cell count NOS CSF increased
C0860829|CSF WBC increased
C0860829|White blood cell count NOS cerebrospinal fluid increased
C0860829|Cerebrospinal fluid WBC increased
C0860829|Cerebrospinal fluid white blood cell count increased
C0860856|White blood cell count semen normal
C0860859|White blood cell count semen high
C1096498|CSF white blood cell count decreased
C1096498|CSF WBC decreased
C1096498|Cerebrospinal fluid WBC decreased
C1096498|Cerebrospinal fluid white blood cell count decreased
C1306872|Granulocytopenia
C1306872|Granulopenia
C1306872|Granulocyte count below reference range (finding)
C1306872|Granulocyte count below reference range
C1960456|Febrile leukopenia
C1960456|Febrile leucopenia
C1960456|Febrile leukopenia (disorder)
C0373807|Leukocyte alkaline phosphatase with count
C0373807|WBC ALKALINE PHOSPHATASE COUNT
C0373807|White blood cell alkaline phosphatase (enzyme) measurement with cell count
C0373807|Leukocyte alkaline phosphatase test with count
C0373807|WBC ALKALINE PHOSPHATASE
C1303089|B CELLS TOTAL COUNT
C1303089|Total B cell count
C1303089|Total cell count for B cells (white blood cells)
C1303089|Total B lymphocyte count (procedure)
C1303089|Total B lymphocyte count
C1303089|B cells, total count
C1504163|NK CELLS TOTAL COUNT
C1504163|NATURAL KILLER CELLS TOTAL COUNT
C1504163|Total cell count for natural killer cells (white blood cell)
C1504163|Total natural killer (NK) cell count
C1504163|Natural killer (NK) cells, total count
C2676078|WBCQ1
C2676078|WHITE BLOOD CELL COUNT QUANTITATIVE TRAIT LOCUS 1
