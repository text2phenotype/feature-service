C0555903|Total protein measurement
C1261360|Total protein result
C0036836|Serum total protein measurement
C0580563|Serum total protein normal
C0580564|Serum total protein abnormal
C0728420|Total Protein Reagent
C0805031|albumin/protein.total
C0855756|Protein total abnormal
C0855757|Protein total normal
C0855758|Protein total increased
C0859351|Serum total protein increased
C0860703|Serum total protein decreased
C0860901|Protein total decreased
C0972523|Protein Determination Reagents, Total
C1168441|total protein S assay
C1168459|Protein S total abnormal
C0555903|Total Protein Measurement
C0555903|Protein total
C0555903|Measurement of total protein
C0555903|Protein
C0555903|PROT
C0555903|Total protein
C0555903|TP - Total protein
C0555903|TPr - Total protein
C0555903|Total protein measurement (procedure)
C0428541|urine total protein measurement (lab test)
C0428541|urine total protein measurement
C0428541|urine total protein
C0428541|Measurement of total protein in urine
C0428541|Total protein level, urine
C0428541|Urine total protein (& level)
C0428541|Urine total protein (& level) (procedure)
C0428541|Urine total protein level
C0428541|Urine total protein measurement (procedure)
C2097239|serum total protein by refractometry (lab test)
C2097239|serum total protein by refractometry
C2097239|total serum protein level by refractometry
C0036836|Serum Total Protein Measurement
C0036836|total serum protein level
C0036836|serum total protein measurement (lab test)
C0036836|serum total protein
C0036836|Serum Protein Total Measurement
C0036836|Total Serum Protein Measurement
C0036836|Measurement of total protein in serum
C0036836|Serum total protein (& level) (procedure)
C0036836|Serum total protein (& level)
C0036836|Serum Total Protein Test
C0036836|Serum total protein level
C0036836|Serum total protein measurement (procedure)
C0855756|Protein total abnormal
C0855756|Protein total abnormal NOS
C0855757|Protein total normal
C0855757|Total protein normal
C0859351|Serum total protein increased
C0855758|Protein total increased
C0855758|Total protein high
C0855758|Protein total high
C0860703|Serum total protein decreased
C0860901|Protein total decreased
C0860901|Decreased total protein
C0860901|Total protein low
C1168441|total protein S assay (lab test)
C1168441|total protein S assay
C1168441|total protein S
C1168441|Assay for total protein S
C1168441|Protein S total
C1168459|Protein S total abnormal
