# HepC : Create "blacklist.bsv" for concepts that hit too many inputs
# 
# JIRA/BIOMED-118
# 
C0030705|Patient
C0037125|Silver

# JIRA/BIOMED-114
#
C1514241|Positive
C1514241|Positive Finding

# JIRA/SANDS-173
# 
C0006826|CA

# JIRA/BIOMED-118
#
C1261327|Family history: Asthma

# JIRA/BIOMED-104
#
C0032854|Poor

# JIRA/BIOMED-124
#
C0007457|Caucasoid Race 
C0043157|Caucasians


# JIRA/BIOMED-145
#
C0424670|Weight for height


# Caroyln Blose
# 
# "Page"  is not an acronym 
#
# [ ['C0013862|T059|MSH|Polyacrylamide Gel Electrophoresis|Page|29|33|positive|None
#
# C042145|DOB|Date of Birth
# C1441613|ID|Immune diffusion
# C0373675|mg|Magnesium 
# C0449201|T029|SNOMEDCT_US|PER tumor staging notation
# C0031381|PCP "Phencyclidine"

JIRA/BIOMED-236
# 
C0013146|Drugs