C0017725|Glucose
C0364479|Glucose
C0364479|Glucose:MCnc:Pt:Bld:Qn
C0337438|Glucose
C0337438|Glucose measurement
C0337438|Test;glucose
C0337438|Measurement of glucose
C0337438|Glucose measurement (procedure)
C0337438|Glucose measurement, NOS
C0337438|glucose test
C0523658|ASSAY GLUCOSE BLOOD QUANT
C0523658|Glucose; quantitative, blood (except reagent strip)
C0523658|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP
C0523658|Glucose measurement, quantitative
C0523658|Glucose measurement, quantitative (procedure)
C0202045|Glucose measurement, fasting
C0428568|Fasting blood glucose measurement
C0005802|Blood Glucose
C0005802|Sugar, Blood
C0005802|blood sugar
C0005802|Blood Glucose [Chemical/Ingredient]
C0005802|Glucose, Blood
C0005802|glycemia
C0011501|2 Deoxy D glucose
C0011501|2 Deoxyglucose
C0011501|2 Desoxy D glucose
C0011501|Deoxyglucose
C0011501|D-arabino-Hexose, 2-deoxy-
C0011501|2-deoxy-D-glucose
C0011501|2-Desoxy-D-glucose
C0011501|Deoxyglucose [Chemical/Ingredient]
C0011501|2-Deoxyglucose
C0011501|2-DG
C0011501|2DG
C0284374|glucosylglycerol
C0055893|1-O-ethyl-5,6-bis-O-(4-chlorobenzyl)-3-O-propyl-D-glucofuranoside
C0055893|clobenosid
C0055893|clobenoside
C0055893|Clobenoside (substance)
C0912322|glucosyl-ifosfamide mustard
C0912322|glufosfamide
C0912322|Beta-D-Glucosyl-Ifosfamide Mustard
C0912322|glc-IPM
C0719353|Citrate-Phos-Dex
C0719831|Dextrose (for TPN)
C0719837|Dextrose and Lactated Ringers and Potassium
C0719843|Dextrose-Heparin Sodium
C0719845|Dextrose-Magnesium Sulfate
C0719847|Dextrose-Pontocaine HCl
C0719848|Dextrose-Ritodrine Hydrochloride
C0720188|Emechek Anti-Nauseant
C0720635|Genfiber
C0720681|Glutol
C0721208|Kao Lectrolyte
C0721257|Konsyl-D
C0721786|Monojel
C0721996|Natural Vegetable Laxative
C0722001|Nausea Control
C0722002|Nausea Relief Medicine
C0723813|Travasol with Dextrose
C0724091|Uni-Laxative
C0724163|V-Lax
C0876014|Dianeal PD-2 with 3.5% Dextrose
C0306071|Emetrol
C0306071|phosphorated carbohydrate solution (Emetrol)
C0306071|carbohydrates (Emetrol)
C0306071|Emetrol for Nausea
C0306309|Glutose
C0306465|Insta-Glucose
C0596620|glucose metabolism
C0598522|O methylglucose
C0017725|D Glucose
C0017725|D-Glucose
C0017725|Dextrose
C0017725|Glucose
C0017725|Dextrose preparation
C0017725|foods dextrose
C0017725|glucose (dextrose)
C0017725|glucose (dextrose) (medication)
C0017725|foods glucose (dextrose)
C0017725|dextrose (medication)
C0017725|Glucose [Chemical/Ingredient]
C0017725|Dextrose preparation (product)
C0017725|D-glucose preparation
C0017725|Dextrose (substance)
C0017725|Glucose [endocrine]
C0017725|Glucose preparation (substance)
C0017725|D-glucopyranose monohydrate preparation
C0017725|Glucose [endocrine] (product)
C0017725|Glucose preparation
C0017725|6-(hydroxymethyl)oxane-2,3,4,5-tetrol
C0017725|DEXTROSE, UNSPECIFIED FORM
C0017725|Dextrose product
C0017725|Glucose product
C0017725|Glucose (substance)
C0017725|Glucose preparation (product)
C0017725|Glucose, NOS
C0017725|Dextrose preparation (substance)
C0017725|Glucose [endocrine] (substance)
C1276933|Glucose 50 MG/ML Irrigation Solution
C1276933|glucose 5 % Irrigation Solution
C1276933|Glucose 5% bladder irrigation (product)
C1276933|Glucose 5% bladder irrigation
C1276933|Glucose 5% bladder irrigation (substance)
C1445695|ALCOHOL/DEXTROSE
C1445695|Alcohol + dextrose (product)
C1445695|Alcohol + dextrose
C2317198|Ophthalmic form glucose (product)
C2317198|Ophthalmic form glucose
C2315494|Oral form glucose (product)
C2315494|Oral form glucose
C2364764|Navstel
C2365303|Dextrose and Electrolyte No. 75
C2586945|Aminosyn II 5% in 25% Dextrose
C2587109|Aminosyn II 3.5 % in 25 % Dextrose
C2608649|Aminosyn II 3.5 % M in 5 % Dextrose
C2608653|Aminosyn II 4.5 % M in 10 % Dextrose
C2717692|Proliferol
C2729519|Dianeal Low Calcium 3.5
C2730298|Nauzene
C1629876|Family Pharmacy brand of Glucose
C0360665|Glucose + Sodium chloride
C0360665|Glucose / Sodium Chloride
C0360665|Dextrose saline
C0360665|Dextrose saline (product)
C0360665|Dextrose saline (substance)
C1445734|DEXTROSE/THEOPHYLLINE
C1445734|Theophylline + dextrose (product)
C1445734|Theophylline + dextrose
C1445772|Milrinone + dextrose (product)
C1445772|Milrinone + dextrose
C1445773|morphine sulfate in dextrose
C1445773|morphine sulfate in dextrose (medication)
C1445773|narcotics morphine sulfate in dextrose
C1445773|Morphine sulfate + dextrose
C1445773|Morphine sulfate + dextrose (product)
C1445773|Morphine sulphate + dextrose
C1445786|Penicillin G + dextrose
C1445786|Penicillin G + dextrose (product)
C1445835|CEFOXITIN/DEXTROSE
C1445835|Cefoxitin + dextrose (product)
C1445835|Cefoxitin + dextrose
C0719849|DEXTROSE/POTASSIUM CHLORIDE/SODIUM CHLORIDE
C0719849|Glucose + Potassium chloride + Sodium chloride
C0719849|Glucose / Potassium Chloride / Sodium Chloride
C0719849|Dextrose + potassium chloride + sodium chloride
C0719849|Glucose + potassium chloride + sodium chloride (product)
C0719838|Glucose + potassium chloride
C0719838|Glucose + potassium chloride (product)
C0719838|DEXTROSE/POTASSIUM CHLORIDE
C0719838|Dextrose + Potassium chloride
C0719838|Dextrose and Potassium Chloride
C0719838|Glucose / Potassium Chloride
C0719838|Dextrose + potassium chloride (product)
C2585875|Hydroxypropyl methylcellulose + glutathione + glucose
C2585875|Hypromellose + glutathione + glucose
C2585875|Hypromellose + glutathione + glucose (product)
C2012248|glucose + vitamin C
C2012248|glucose + ascorbic acid
C2012248|foods dextrose glucose + vitamin C
C2012248|glucose + ascorbic acid (medication)
C2012248|Ascorbic Acid / Glucose
C0773380|Glucose 700 MG/ML Injectable Solution
C0773380|Dextrose 70% and Water, Dextrose 70% in Water intravenous solution
C0773380|Dextrose 70% Solution for injection
C0773380|parenteral nutrition solution Dextrose 70% in Water intravenous solution
C0773380|Dextrose Inj 70%
C0773380|DEXTROSE 70% INJ
C0773380|DEXTROSE 70% INJ [VA Product]
C0773380|DEXTROSE MONOHYDRATE 70 g in 100 mL INTRAVENOUS INJECTION, SOLUTION [Dextrose]
C0773380|dextrose 70 % Injectable Solution
C0773380|DEXTROSE 70 g in 100 mL INTRAVENOUS SOLUTION
C0773380|Glucose 70% intravenous infusion
C0773380|Glucose 70% infusion solution bag (product)
C0773380|Glucose 70% infusion solution bag
C0773380|Glucose 70% intravenous infusion (product)
C0773380|Glucose 70% intravenous infusion (substance)
C0773380|Dextrose 70% Intravenous Solution
C0976237|Glucose 50 MG/ML Injectable Solution
C0976237|Dextrose (Diagnostic Aid) Inj 5%
C0976237|Dextrose 5% and Water, Dextrose 5% in Water intravenous solution
C0976237|Dextrose 5% Solution for injection
C0976237|LVP solution Dextrose 5% in Water intravenous solution
C0976237|DEXTROSE 5% INJ BAG 50ML
C0976237|DEXTROSE 5% INJ BAG 250ML
C0976237|DEXTROSE 5% INJ BAG 100ML
C0976237|DEXTROSE 5% INJ BAG 150ML
C0976237|DEXTROSE 5% INJ BAG 1000ML
C0976237|DEXTROSE 5% INJ
C0976237|DEXTROSE 5% INJ BAG 500ML
C0976237|Dextrose Inj 5%
C0976237|DEXTROSE 5% INJ,BAG,150ML [VA Product]
C0976237|DEXTROSE 5% INJ,BAG,250ML
C0976237|DEXTROSE 5% INJ,BAG,250ML [VA Product]
C0976237|DEXTROSE 5% INJ [VA Product]
C0976237|DEXTROSE 5% INJ,BAG,1000ML
C0976237|DEXTROSE 5% INJ,BAG,50ML [VA Product]
C0976237|DEXTROSE 5% INJ,BAG,1000ML [VA Product]
C0976237|DEXTROSE 5% INJ,BAG,50ML
C0976237|DEXTROSE 5% INJ,BAG 100ML
C0976237|DEXTROSE 5% INJ,BAG 100ML [VA Product]
C0976237|DEXTROSE 5% INJ,BAG,150ML
C0976237|DEXTROSE 5% INJ,BAG,500ML [VA Product]
C0976237|DEXTROSE MONOHYDRATE 50 g in 1000 mL INTRAVENOUS INJECTION, SOLUTION [DEXTROSE]
C0976237|DEXTROSE 5% INJ,BAG,500ML
C0976237|Dextrose 5% and Water ADD-Vantage, Dextrose 5% in Water intravenous solution
C0976237|dextrose 50 MG/ML Injectable Solution
C0976237|dextrose 5 % Injectable Solution
C0976237|DEXTROSE MONOHYDRATE 50 mg in 1 mL INTRAVENOUS INJECTION, SOLUTION [Dextrose]
C0976237|DEXTROSE 5 g in 100 mL INTRAVENOUS SOLUTION
C0976237|DEXTROSE MONOHYDRATE 5 g in 100 mL INTRAVENOUS INJECTION, SOLUTION
C0976237|dextrose 5 GM per 100 ML Injectable Solution
C0976237|DEXTROSE MONOHYDRATE 5 g in 100 mL INTRAVENOUS INJECTION, SOLUTION [Dextrose]
C0976237|DEXTROSE MONOHYDRATE 50 mg in 1 mL INTRAVENOUS INJECTION, SOLUTION
C0976237|Dextrose 5% Injection Solution
C0976237|Dextrose 5g/100mL injection (product)
C0976237|Dextrose 5g/100mL injection
C0976237|DEXTROSE MONOHYDRATE 50 g in 1000 mL INTRAVENOUS INJECTION, SOLUTION [Veterinary Dextrose]
C0976237|DEXTROSE MONOHYDRATE 5 g in 100 mL INTRAVENOUS INJECTION [Dextrose]
C0976237|DEXTROSE MONOHYDRATE 5 g in 100 mL INTRAVENOUS INJECTION, SOLUTION [Veterinary 5% Dextrose]
C0976237|Glucose 5% infusion
C0976237|Dextrose 5% injection solution ampoule
C0976237|Dextrose 5% injection solution ampule (product)
C0976237|Dextrose 5% injection solution ampule
C0976237|Dextrose 5g/100mL (5%) injection solution 1000mL vial (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 1000mL vial
C0976237|Dextrose 5g/100mL (5%) injection solution 100mL vial (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 100mL vial
C0976237|Dextrose 5g/100mL (5%) injection solution 150mL bottle (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 150mL bottle
C0976237|Dextrose 5g/100mL (5%) injection solution 150mL vial (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 150mL vial
C0976237|Dextrose 5g/100mL (5%) injection solution 250mL bottle (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 250mL bottle
C0976237|Dextrose 5g/100mL (5%) injection solution 25mL vial (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 25mL vial
C0976237|Dextrose 5g/100mL (5%) injection solution 500mL vial (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 500mL vial
C0976237|Dextrose 5g/100mL (5%) injection solution 50mL vial (product)
C0976237|Dextrose 5g/100mL (5%) injection solution 50mL vial
C0976237|Glucose 5% infusion solution bottle (product)
C0976237|Glucose 5% infusion solution bottle
C0976237|Glucose 5% infusion solution 1 L bag (product)
C0976237|Glucose 5% infusion solution 1 L bag
C0976237|Glucose 5% infusion solution 100 mL bag (product)
C0976237|Glucose 5% infusion solution 100 mL bag
C0976237|Glucose 5% infusion solution 150 mL bag (product)
C0976237|Glucose 5% infusion solution 150 mL bag
C0976237|Glucose 5% infusion solution 250 mL bag (product)
C0976237|Glucose 5% infusion solution 250 mL bag
C0976237|Dextrose 5% injection solution ampoule (product)
C0976237|Glucose 5% infusion (product)
C0976237|Glucose 5% infusion (substance)
C0976237|Dextrose 5% Intravenous Solution
C0784132|Glucose 380 MG/ML Injectable Solution
C0784132|DEXTROSE 38% INJ
C0784132|DEXTROSE 38% INJ [VA Product]
C0784132|dextrose 38 % Injectable Solution
C0784132|glucose 38 % Injectable Solution
C0976216|DEXTROSE 100% PWDR
C0976216|DEXTROSE 100% PWDR [VA Product]
C0691368|Dextrose 100g/180mL Oral solution
C0691368|DEXTROSE 100GM/180ML LIQUID
C0691368|DEXTROSE 100GM/180ML [VA Product]
C0691368|DEXTROSE 100GM/180ML
C0691368|Dextrose 100 GM/180 ML Oral Solution
C0691368|glucose 100 g/180 mL oral liquid
C0976227|Glucose 0.417 MG/MG Oral Gel
C0976227|DEXTROSE 25GM/60GM SQUEEZE TUBE
C0976227|DEXTROSE 25GM/60GM SQUEEZE TUBE [VA Product]
C0976227|glucose 25 GM per 60 GM Oral Gel
C0691497|Glucose 0.4 MG/MG Oral Gel
C0691497|CVS Glucose, 40% oral gel
C0691497|Dextrose 15 GM Oral Gel/Jelly
C0691497|Glucose Gel, 40% oral gel
C0691497|DEXTROSE 15GM/45GM SQUEEZE TUBE
C0691497|Dextrose 40% Oral gel
C0691497|glucose 40% oral gel
C0691497|DEXTROSE 15GM/37.5GM SQUEEZE TUBE
C0691497|DEXTROSE 18GM/45GM SQUEEZE TUBE
C0691497|DEXTROSE 32GM/80GM SQUEEZE TUBE
C0691497|Glucose Gel 40%
C0691497|DEXTROSE 15GM/37.5GM SQUEEZE TUBE [VA Product]
C0691497|DEXTROSE 32GM/80GM SQUEEZE TUBE [VA Product]
C0691497|DEXTROSE 18GM/45GM SQUEEZE TUBE [VA Product]
C0691497|DEXTROSE 15GM/45GM SQUEEZE TUBE [VA Product]
C0691497|dextrose 40 % Oral Gel
C0691497|DEXTROSE 40% GEL,ORAL
C0691497|DEXTROSE 40% ORAL GEL (GLUCOSE)
C0691497|DEXTROSE 40% GEL,ORAL [VA Product]
C0691497|Glucose 15g Oral gel
C0691497|glucose 18 GM per 45 GM Oral Gel
C0691497|glucose 32 GM per 80 GM Oral Gel
C0691497|glucose 15 GM per 37.5 GM Oral Gel
C0691497|Dextrose 40% oral gel (product)
C0691497|Dextrose 40% oral gel (substance)
C0691497|Dextrose 40% Oral Gel/Jelly
C0982177|GLUCOSE LIQUID
C0977174|Glucose 5000 MG Chewable Tablet
C0977174|GLUCOSE 5GM CHEW TAB
C0977174|Glucose Chew Tab 5 GM
C0977174|GLUCOSE 5GM TAB,CHEW [VA Product]
C0977174|GLUCOSE 5GM TAB,CHEW
C0977174|Glucose 5g Chewable tablet
C0977174|Dextrose 5 GM Oral Tablet, Chewable [GLUTOSE]
C0977174|glucose 5 GM Chewable Tablet
C0977174|Dextrose 5 GM Oral Tablet, Chewable
C0977174|Glucose, 5 g oral tablet, chewable
C0977174|glucose 5 g oral tablet, chewable
C0977171|GLUCOSE 24GM ORAL LIQUID
C0977171|GLUCOSE 24GM LIQUID,ORAL
C0977171|GLUCOSE 24GM LIQUID,ORAL [VA Product]
C2931948|amino-acid, glucose, and electrolyte solution
C0985452|Glucose 50 MG/ML
C0985452|Dextrose 5%
C2961328|GLUCOSE 50GM/300ML ORAL LIQUID
C2961328|glucose 50 GM per 300 ML Oral Solution
C2961328|GLUCOSE 50GM/300ML LIQUID,ORAL
C2961328|GLUCOSE 50GM/300ML LIQUID,ORAL [VA Product]
C2961328|Glucose 166.7 MG/ML Oral Solution
C2962383|Enfamil Glucose
C2979326|Clinimix E 4.25/10
C2979448|Naus-Aid
C1634042|Longs Glucose
C1628288|Leader brand of glucose
C3152484|Elliotts B
C0050552|ACD solution
C0050552|acid citrate dextrose
C0050552|D-glucose, 2-hydroxy-1,2,3-propanetricarboxylate (1:1) (salt)
C0050552|Acid-Citrate-Dextrose
C0050552|ACD
C0605504|beta-D-Glucopyranosyl isothiocyanate
C0605504|beta-D-glucopyranosylisothiocyanate
C0624467|G-6-VAN
C0624467|glucose-6-vanadate
C0044547|1-O-octadecyl-2-O-methylglycerol-3-glucopyranoside
C0044547|OMGGP
C0116601|6-O-butanoyl-1,2-O-isopropylidene-alpha-D-glucofuranose
C0116601|esterbut-6
C0116601|MAG-6BUT
C0116601|monoacetone glucose 6-butyrate
C0116601|monobut-6
C0116600|3-O-butanoyl-1,2-O-isopropylidene-alpha-D-glucofuranose
C0116600|esterbut-3
C0116600|MAG-3BUT
C0116600|monoacetone glucose 3-butyrate
C0116600|monobut-3
C0116600|3n-But
C0116600|3n-butyrate
C0166821|CDP-D-glucose
C0166821|CDP-glucose
C0166821|cytidine diphosphate-glucose
C0212338|Glu-1-MePhos
C0212338|glucose-1-methylenephosphonate
C0657081|repandusinic acid A
C0660803|sarmentosine
C0660804|glucofructan
C0660981|glucose phenylosazone
C0660981|D-arabino-Hexos-2-ulose, bis(phenylhydrazone)
C0660981|glucosephenylosazone
C0662439|pedunculoside
C0257753|glucose aldonitrile pentaacetate
C0385852|2-MTAD-glucopyrano-doxaz
C0385852|2-methyl-(3,4,6-tri-O-acetyl-1,2-dideoxyglucopyrano)(2,1-d)-2-oxazoline
C0387981|3-Azi-Glc
C0387981|3-deoxy-3,3-azi-D-glucopyranose
C0387981|3-deoxy-3,3-aziglucopyranose
C0388846|N-(beta-D-glucopyranosyl)nicotinic acid
C0388846|N-glucopyranosylnicotinic acid
C0534039|dTDP-glucose
C0534039|deoxythymidine diphosphate-glucose
C0675321|dTDP-6-deoxy-4-ketoglucose
C0675321|dTDP-KDG
C0675321|TDP-4-keto-6-deoxy-D-glucose
C0759361|4,6-O-(4'-iodoethylidene)glucose
C0759361|4'-IEDG
C0759364|4,6-O-(2'-iodoethylidene)glucose
C0759364|2'-IEDG
C0767580|3,9-dibromo-12-(4-O-methylglucopyranosyl)-6,7.12,13-tetrahydroindolo(2,3-a)pyrrolo(3,4-c)carbazole-5,7-dione
C0767580|3,9-dibromo-MGTIPCD
C0768175|glucoerucin
C0768409|6-C-glucosylnalingenin
C0768410|6-C-glucosylaronadendrin
C0768878|2-(2,4,5-trihydroxyphenyl)-3,5,7-trihydroxy-6-C-glucopyranosyloxy-4H-1-benzopyran-4-one
C0768878|shamimin
C0910124|glucose-2-SNAP
C0911387|Tc-99m-thio-D-glucose
C0912160|3-O-butanoyl-1,2:5,6-di-O-isopropylidene-alpha-D-glucose
C0912160|diacetone glucose butyrate
C0912161|1,2,3,4,6-penta-O-butanoyl-alpha-D-glucose
C0912161|glucose pentabutyrate
C0967100|4,6-O-isoterchebuloyl-D-glucose
C0967100|4,6-O-isoterchebuloylglucose
C0967100|4,6-O-iso-terchebuloylglucose
C1097389|(((1,2-5,6-di-O,O-isopropylideneglucofuranos-3-yl)oxocarbonyl)methyl)cobalt tricarbonyl triphenylphosphine
C1097389|iPGlcf-ocometctpp
C1172347|3-O-benzyl-6-O-pivaloylglucopyranose 1,2,4-orthopivalate
C1172982|1-O-methyl-6-O-caffeoylglucopyranose
C1436637|N,beta-D-Glucopyranosyl vincosamide
C1436637|N-GP-VA
C1530900|TPC(m-O-Glu)(3)
C1530900|tri(glucosyloxyphenyl)chlorin
C1609691|beta-D-glucopyranosyl bismethoxyphosphoramidate
C1609691|beta-Glu-BMPA
C1700327|2,3,4,6-tetra-O-acetyl-1-thioglucopyranose
C1702259|glucopyranose spirohydantoin
C1743143|1,6-anhydro-3,4-dideoxyhex-3-enopyran-2-ulose
C2604528|FEtGlc-triazoles
C2604528|4-(2-fluoroethyl)-1-glucopyranosyl-1H-1,2,3-triazole
C2606058|6-O-octanoylglucose
C2715303|glucopyranosylidene-spiro-oxathiazole
C2932471|1,6-diferuloyl glucose
C2932910|1-benzoyl-NPGlc-TI
C2932910|1-benzoyl-4-(4-nitrophenyl)-3-glucopyranosylthiazol-2(3H)-imine
C2935358|trans-resveratrol-4'-O-beta-D-glucopyranoside
C2974270|dansyl C-glucoside
C2587130|Aminosyn II 3.5 % with Electrolytes in 25 % Dextrose with Calcium
C2587136|Aminosyn II 4.25 % with Electrolytes in 25 % Dextrose with Calcium
C1725310|Isolyte S and 5% Dextrose
C1725310|Isolyte S in 5 % Dextrose
C0722153|Normosol-R and 5% Dextrose
C0722153|Normosol-R in 5 % Dextrose
C1657070|Plasma-Lyte 148 in 5 % Dextrose
C1657070|Dextrose 5% and Plasma-Lyte 148
C2345938|Plasma-Lyte 56 in 5 % Dextrose
C2345938|Plasma-Lyte 56 and 5% Dextrose
C2346377|Plasma-Lyte M in 5 % Dextrose
C2346182|Travasol 5.5 % in Dextrose
C2346366|Plasma-Lyte R in 5 % Dextrose
C1657537|Dextrose Hydrous
C1657537|dextrose (hydrous)
C3474002|Dextrose monohydrate
C3473090|GlucoBurst
C3556165|TRUEplus Glucose
C3643617|ReliOn Glucose
C0002272|alpha Glucosidases
C0002272|alpha-Glucosidases
C0002272|Maltase Glucoamylase
C0002272|alpha glucosidase
C0002272|alpha-D-Glucoside glucohydrolases
C0002272|glucoinvertase
C0002272|glucosidosucrase
C0002272|maltase
C0002272|Alpha-glucosidase
C0002272|Maltase-Glucoamylase
C0002272|alpha-Glucosidases [Chemical/Ingredient]
C0002272|Maltases
C0002272|alpha-Glucosidase (substance)
C0002272|Alpha glucosidase (product)
C0002272|alpha-Glucosidase [dup] (substance)
C1273905|Dextrose + lidocaine hydrochloride 75mg/50mg
C1273905|Dextrose + lidocaine hydrochloride 75mg/50mg (product)
C1273905|Dextrose+lidocaine hydrochloride 75mg/50mg
C1533829|Dextrose + lidocaine hydrochloride 7.5%ww/1.5%ww injection
C1533829|Dextrose + lidocaine hydrochloride 7.5%ww/1.5%ww injection (product)
C1533820|Bupivacaine hydrochloride + dextrose 7.5mg/82.5mg injection
C1533820|Bupivacaine hydrochloride + dextrose 7.5mg/82.5mg injection (product)
C0359952|BUPIVACAINE/DEXTROSE
C0359952|local anesthetics bupivacaine in dextrose
C0359952|bupivacaine in dextrose (medication)
C0359952|bupivacaine in dextrose
C0359952|Bupivacaine + Glucose
C0359952|Bupivacaine + dextrose (product)
C0359952|Bupivacaine + dextrose
C0359952|Bupivacaine+glucose
C0359952|Bupivacaine hydrochloride+glucose
C0359952|Bupivacaine+glucose (product)
C0359952|Bupivacaine+glucose (substance)
C0773377|Glucose 600 MG/ML Injectable Solution
C0773377|Dextrose 60% and Water, Dextrose 60% in Water intravenous solution
C0773377|Dextrose 60% Solution for injection
C0773377|parenteral nutrition solution Dextrose 60% in Water intravenous solution
C0773377|DEXTROSE 60% INJ
C0773377|DEXTROSE 60% INJ [VA Product]
C0773377|dextrose 60 % Injectable Solution
C0773377|Dextrose 60g injection (product)
C0773377|Dextrose 60g injection
C0773377|Dextrose 60% in water intravenous solution 1000mL bag (product)
C0773377|Dextrose 60% in water intravenous solution 1000mL bag
C0773377|Dextrose 60% in water intravenous solution 500mL bag (product)
C0773377|Dextrose 60% in water intravenous solution 500mL bag
C0773377|Dextrose 60% Intravenous Solution
C1165353|dextrose anhydrous
C1165353|Anhydrous Dextrose
C1165353|Dextrose, Anhydrous
C1876722|Beta-D-Glucopyranose
C1876722|.BETA.-D-GLUCOPYRANOSE
C0549987|Glucose [Presence] in Urine by Test strip --4.5 hours post 75 g glucose PO
C0549987|Glucose^4.5H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0549987|Glucose^4.5 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0549987|Glucose 4.5h p 75 g Glc PO Ur Ql Strip
C0363629|Glucose [Mass/volume] in Urine --1.5 hours post 100 g glucose PO
C0363629|Glucose^1.5H post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363629|Glucose^1 1/2 hour post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363629|Glucose 1.5h p 100 g Glc PO Ur-mCnc
C0363633|Glucose [Mass/volume] in Serum or Plasma --1 hour post 0.5 g/kg glucose IV
C0363633|Glucose^1H post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363633|Glucose^1 hour post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363633|Glucose 1h p .5 g/kg Glc IV SerPl-mCnc
C0797929|Glucose [Moles/volume] in Serum or Plasma --1 hour post 50 g lactose PO
C0797929|Glucose^1H post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C0797929|Glucose^1 hour post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797929|Glucose 1h p 50 g Lac PO SerPl-sCnc
C0797936|Glucose [Moles/volume] in Serum or Plasma --30 minutes post 50 g lactose PO
C0797936|Glucose 30M p 50 g Lac PO SerPl-sCnc
C0797936|Glucose^30M post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C0797936|Glucose^30 minutes post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797944|Glucose^post CFst:SCnc:Pt:BldC:Qn:Glucometer
C0797944|Fasting glucose [Moles/volume] in Capillary blood by Glucometer
C0797944|Glucose p fast BldC Glucomtr-sCnc
C0797944|Glucose^post Calorie fast:Substance Concentration:Point in time:Blood capillary:Quantitative:Glucometer
C0549989|Glucose^45M post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0549989|Glucose [Mass/volume] in Serum or Plasma --45 minutes post 50 g lactose PO
C0549989|Glucose 45M p 50 g Lac PO SerPl-mCnc
C0549989|Glucose^45M post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549978|Glucose sp1 p chal SerPl-mCnc
C0549978|Glucose^1st specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549978|Glucose [Mass/volume] in Serum or Plasma --1st specimen post XXX challenge
C0549978|Glucose^1st specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549976|Glucose^15th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549976|Glucose [Mass/volume] in Serum or Plasma --15th specimen post XXX challenge
C0549976|Glucose sp15 p chal SerPl-mCnc
C0549976|Glucose^15th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549992|Glucose [Mass/volume] in Serum or Plasma --50 minutes post XXX challenge
C0549992|Glucose 50M p chal SerPl-mCnc
C0549992|Glucose^50M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549992|Glucose^50M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544010|Glucose [Mass/volume] in Serum or Plasma --pre XXX challenge
C1544010|Glucose pre chal SerPl-mCnc
C1544010|Glucose^pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544010|Glucose^pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544022|Glucose^12.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544022|Glucose [Mass/volume] in Serum or Plasma --12.5 hours post XXX challenge
C1544022|Glucose 12.5h p chal SerPl-mCnc
C1544022|Glucose^12.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544027|Glucose^16H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544027|Glucose 16h p chal SerPl-mCnc
C1544027|Glucose [Mass/volume] in Serum or Plasma --16 hours post XXX challenge
C1544027|Glucose^16H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544030|Glucose^18.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544030|Glucose [Mass/volume] in Serum or Plasma --18.5 hours post XXX challenge
C1544030|Glucose 18.5h p chal SerPl-mCnc
C1544030|Glucose^18.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544033|Glucose^20.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544033|Glucose [Mass/volume] in Serum or Plasma --20.5 hours post XXX challenge
C1544033|Glucose^20.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544033|Glucose 20.5h p chal SerPl-mCnc
C1544040|Glucose [Mass/volume] in Serum or Plasma --9 minutes post XXX challenge
C1544040|Glucose 9M p chal SerPl-mCnc
C1544040|Glucose^9M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544040|Glucose^9 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542932|Glucose [Mass/volume] in Serum or Plasma --31 hour post XXX challenge
C1542932|Glucose^31H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1542932|Glucose^31H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542932|Glucose 31h p chal SerPl-mCnc
C1544161|Glucose^11.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544161|Glucose [Moles/volume] in Serum or Plasma --11.5 hours post XXX challenge
C1544161|Glucose^11.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544161|Glucose 11.5h p chal SerPl-sCnc
C1544236|Glucose [Mass/volume] in Serum or Plasma --10.75 hours post XXX challenge
C1544236|Glucose^10.75H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544236|Glucose 10.75h p chal SerPl-mCnc
C1544236|Glucose^10.75H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954700|Glucose^3 AM specimen:MCnc:Pt:Ser/Plas:Qn
C1954700|Glucose [Mass/volume] in Serum or Plasma --3 AM specimen
C1954700|Glucose 3 AM SerPl-mCnc
C1954700|Glucose^3 AM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954185|Glucose Pre fructose PO SerPl-mCnc
C1954185|Glucose^pre dose fructose PO:MCnc:Pt:Ser/Plas:Qn
C1954185|Glucose [Mass/volume] in Serum or Plasma --pre dose fructose PO
C1954185|Glucose^pre dose fructose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706818|Glucose^6M post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706818|Glucose [Moles/volume] in Serum or Plasma --6 minutes post dose glucagon
C2706818|Glucose 6M p Gc SerPl-sCnc
C2706818|Glucose^6 minutes post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706903|Glucose [Moles/volume] in Serum or Plasma --6th specimen post XXX challenge
C2706903|Glucose^6th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2706903|Glucose sp6 p chal SerPl-sCnc
C2706903|Glucose^6th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924063|Glucose 3 PM SerPl-sCnc
C2924063|Glucose^3 PM specimen:SCnc:Pt:Ser/Plas:Qn
C2924063|Glucose [Moles/volume] in Serum or Plasma --3 PM specimen
C2924063|Glucose^3 PM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3533046|Glucose.serum-glucose.synv fld
C0484592|Glucose^4.5H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484592|Glucose [Mass/volume] in Serum or Plasma --4.5 hours post 100 g glucose PO
C0484592|Glucose^4.5 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484592|Glucose 4.5h p 100 g Glc PO SerPl-mCnc
C0799331|Glucose^11 AM specimen:MCnc:Pt:Ser/Plas:Qn
C0799331|Glucose 11 AM SerPl-mCnc
C0799331|Glucose [Mass/volume] in Serum or Plasma --11 AM specimen
C0799331|Glucose^11 AM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0550006|Glucose^pre dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0550006|Glucose [Mass/volume] in Serum or Plasma --pre dose lactose PO
C0550006|Glucose pre Lac PO SerPl-mCnc
C0550006|Glucose^pre dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803254|Glucose^30M post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0803254|Glucose [Mass/volume] in Serum or Plasma --30 minutes post dose glucose
C0803254|Glucose 30M p Glc SerPl-mCnc
C0803254|Glucose^30 minutes post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544031|Glucose [Mass/volume] in Serum or Plasma --19.5 hours post XXX challenge
C1544031|Glucose^19.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544031|Glucose 19.5h p chal SerPl-mCnc
C1544031|Glucose^19.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544046|Glucose^25M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544046|Glucose 25M p chal SerPl-mCnc
C1544046|Glucose [Mass/volume] in Serum or Plasma --25 minutes post XXX challenge
C1544046|Glucose^25 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544047|Glucose [Mass/volume] in Serum or Plasma --27 minutes post XXX challenge
C1544047|Glucose^27M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544047|Glucose 27M p chal SerPl-mCnc
C1544047|Glucose^27M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542934|Glucose [Mass/volume] in Serum or Plasma --2 days post XXX challenge
C1542934|Glucose^2D post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1542934|Glucose 2D p chal SerPl-mCnc
C1542934|Glucose^2 days post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544153|Glucose^50M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544153|Glucose 50M p chal SerPl-sCnc
C1544153|Glucose [Moles/volume] in Serum or Plasma --50 minutes post XXX challenge
C1544153|Glucose^50M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544154|Glucose 70M p chal SerPl-sCnc
C1544154|Glucose [Moles/volume] in Serum or Plasma --70 minutes post XXX challenge
C1544154|Glucose^70M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544154|Glucose^70M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544177|Glucose [Moles/volume] in Serum or Plasma --23.5 hours post XXX challenge
C1544177|Glucose^23.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544177|Glucose^23.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544177|Glucose 23.5h p chal SerPl-sCnc
C1544262|Glucose [Moles/volume] in Serum or Plasma --105 minutes post dose glucose
C1544262|Glucose^105M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1544262|Glucose 105M p Glc SerPl-sCnc
C1544262|Glucose^105M post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542947|Glucose [Moles/volume] in Serum or Plasma --9 minutes post XXX challenge
C1542947|Glucose^9M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542947|Glucose 9M p chal SerPl-sCnc
C1542947|Glucose^9 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544195|Glucose^29H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544195|Glucose [Moles/volume] in Serum or Plasma --29 hours post XXX challenge
C1544195|Glucose^29H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544195|Glucose 29h p chal SerPl-sCnc
C1544805|Glucose sp2 p chal Ur Strip-mCnc
C1544805|Glucose [Mass/volume] in Urine by Test strip --2nd specimen post XXX challenge
C1544805|Glucose^2nd specimen post XXX challenge:MCnc:Pt:Urine:Qn:Test strip
C1544805|Glucose^2nd specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C1644627|Glucose p fast BldC Glucomtr-mCnc
C1644627|Glucose^post CFst:MCnc:Pt:BldC:Qn:Glucometer
C1644627|Fasting glucose [Mass/volume] in Capillary blood by Glucometer
C1644627|Glucose^post Calorie fast:Mass Concentration:Point in time:Blood capillary:Quantitative:Glucometer
C1954462|Glucose [Mass/volume] in Serum or Plasma --5 hours post 50 g glucose PO
C1954462|Glucose^5H post 50 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C1954462|Glucose^5 hours post 50 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954462|Glucose 5h p 50 g Glu PO SerPl-mCnc
C2706839|Glucose^1H post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706839|Glucose [Moles/volume] in Serum or Plasma --1 hour post dose ornithine alpha-ketoglutarate
C2706839|Glucose^1 hour post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706839|Glucose 1h p OKG SerPl-sCnc
C3172453|Glucose^post CFst:MCnc:Pt:Urine:Qn
C3172453|Glucose p fast Ur-mCnc
C3172453|Glucose^post Calorie fast:Mass Concentration:Point in time:Urine:Quantitative
C3172453|Fasting glucose [Mass/volume] in Urine
C1988504|Glucose tolerance &#x7C; bld-ser-plas
C0942503|Glucose^4H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942503|Glucose [Presence] in Urine by Test strip --4 hours post dose glucose
C0942503|Glucose^4 hours post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0942503|Glucose 4h p Glc Ur Ql Strip
C0942505|Glucose^6H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942505|Glucose [Presence] in Urine by Test strip --6 hours post dose glucose
C0942505|Glucose^6 hours post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0942505|Glucose 6h p Glc Ur Ql Strip
C0941766|Glucose^45M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C0941766|Glucose [Moles/volume] in Serum or Plasma --45 minutes post XXX challenge
C0941766|Glucose 45M p chal SerPl-sCnc
C0941766|Glucose^45M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1316521|Glucose pre/p Gc SerPl-sCnc
C1316521|Glucose^pre or post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C1316521|Glucose^pre or post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1316521|Glucose [Moles/volume] in Serum or Plasma --pre or post dose glucagon
C1544049|Glucose^5.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544049|Glucose [Mass/volume] in Serum or Plasma --5.5 hours post XXX challenge
C1544049|Glucose^5.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544049|Glucose 5.5h p chal SerPl-mCnc
C1544051|Glucose^26H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544051|Glucose [Mass/volume] in Serum or Plasma --26 hours post XXX challenge
C1544051|Glucose^26H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544051|Glucose 26h p chal SerPl-mCnc
C1716428|Glucose^45M post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C1716428|Glucose [Moles/volume] in Serum or Plasma --45 minutes post dose lactose PO
C1716428|Glucose 45M p Lac PO SerPl-sCnc
C1716428|Glucose^45M post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2360466|Glucose^3H post dose fructose PO:MCnc:Pt:Ser/Plas:Qn
C2360466|Glucose [Mass/volume] in Serum or Plasma --3 hours post dose fructose PO
C2360466|Glucose^3 hours post dose fructose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2360466|Glucose 3h p fructose PO SerPl-mCnc
C2925729|Glucose [Moles/volume] in Urine by Automated test strip
C2925729|Glucose Ur Strip.auto-sCnc
C2925729|Glucose:SCnc:Pt:Urine:Qn:Test strip.automated
C2925729|Glucose:Substance Concentration:Point in time:Urine:Quantitative:Test strip.automated
C2706836|Glucose^3H post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706836|Glucose [Moles/volume] in Serum or Plasma --3 hours post dose ornithine alpha-ketoglutarate
C2706836|Glucose^3 hours post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706836|Glucose 3h p OKG SerPl-sCnc
C2706904|Glucose [Moles/volume] in Serum or Plasma --7th specimen post XXX challenge
C2706904|Glucose sp7 p chal SerPl-sCnc
C2706904|Glucose^7th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2706904|Glucose^7th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1988515|Glucose.protein bound &#x7C; bld-ser-plas
C0363664|Glucose^3H post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363664|Glucose [Mass/volume] in Urine --3 hours post 100 g glucose PO
C0363664|Glucose^3 hours post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363664|Glucose 3h p 100 g Glc PO Ur-mCnc
C0800048|Glucose p chal SerPl-mCnc
C0800048|Glucose [Mass/volume] in Serum or Plasma --post XXX challenge
C0800048|Glucose^post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0800048|Glucose^post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363631|Glucose^1.5H post dose insulin IV:MCnc:Pt:Ser/Plas:Qn
C0363631|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post dose insulin IV
C0363631|Glucose^1 1/2 hour post dose insulin Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363631|Glucose 1.5h p Ins IV SerPl-mCnc
C0797939|Glucose^3H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0797939|Glucose [Moles/volume] in Serum or Plasma --3 hours post dose glucose
C0797939|Glucose^3 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797939|Glucose 3h p Glc SerPl-sCnc
C0363687|Glucose^post CFst:MCnc:Pt:BldC:Qn
C0363687|Fasting glucose [Mass/volume] in Capillary blood
C0363687|Glucose p fast BldC-mCnc
C0363687|Glucose^post Calorie fast:Mass Concentration:Point in time:Blood capillary:Quantitative
C1114131|Glucose^3.6H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114131|Glucose [Moles/volume] in Serum or Plasma --3.6 hours post dose glucose
C1114131|Glucose^3.6 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114131|Glucose 3.6h p Glc SerPl-sCnc
C1544029|Glucose [Mass/volume] in Serum or Plasma --18 hours post XXX challenge
C1544029|Glucose^18H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544029|Glucose 18h p chal SerPl-mCnc
C1544029|Glucose^18H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544147|Glucose [Moles/volume] in Serum or Plasma --5 minutes pre XXX challenge
C1544147|Glucose^5M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544147|Glucose 5M pre chal SerPl-sCnc
C1544147|Glucose^5 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544159|Glucose^10H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544159|Glucose [Moles/volume] in Serum or Plasma --10 hours post XXX challenge
C1544159|Glucose^10H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544159|Glucose 10h p chal SerPl-sCnc
C1544184|Glucose [Moles/volume] in Serum or Plasma --2 minutes post XXX challenge
C1544184|Glucose 2M p chal SerPl-sCnc
C1544184|Glucose^2M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544184|Glucose^2 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544188|Glucose [Moles/volume] in Serum or Plasma --3.5 hours post XXX challenge
C1544188|Glucose^3.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544188|Glucose^3.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544188|Glucose 3.5h p chal SerPl-sCnc
C1544194|Glucose^28H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544194|Glucose [Moles/volume] in Serum or Plasma --28 hours post XXX challenge
C1544194|Glucose^28H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544194|Glucose 28h p chal SerPl-sCnc
C1544804|Glucose [Mass/volume] in Urine by Test strip --1st specimen post XXX challenge
C1544804|Glucose sp1 p chal Ur Strip-mCnc
C1544804|Glucose^1st specimen post XXX challenge:MCnc:Pt:Urine:Qn:Test strip
C1544804|Glucose^1st specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C1544971|Glucose [Mass/volume] in Serum or Plasma --2 hours post 50 g glucose PO
C1544971|Glucose^2H post 50 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C1544971|Glucose^2 hours post 50 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544971|Glucose 2h p 50 g Glu PO SerPl-mCnc
C1953512|Glucose 15M pre glc SerPl-sCnc
C1953512|Glucose^15M pre dose glucose:SCnc:Pt:Ser/Plas:Qn
C1953512|Glucose [Moles/volume] in Serum or Plasma --15 minutes pre dose glucose
C1953512|Glucose^15 minutes pre dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706811|Glucose^10M pre dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706811|Glucose 10M pre Gc SerPl-sCnc
C2706811|Glucose [Moles/volume] in Serum or Plasma --10 minutes pre dose glucagon
C2706811|Glucose^10 minutes pre dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706817|Glucose^5M pre dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706817|Glucose [Moles/volume] in Serum or Plasma --5 minutes pre dose glucagon
C2706817|Glucose 5M pre Gc SerPl-sCnc
C2706817|Glucose^5 minutes pre dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706820|Glucose^pre dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706820|Glucose [Moles/volume] in Serum or Plasma --pre dose insulin IV
C2706820|Glucose pre Ins IV SerPl-sCnc
C2706820|Glucose^pre dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598585|Glucose [Moles/volume] in Serum or Plasma --2.5 hours post dose betaxolol
C2598585|Glucose^2.5H post dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598585|Glucose^2 1/2 hours post dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598585|Glucose 2.5h p betaxolol SerPl-sCnc
C3533045|Glucose.serum-glucose.perition fld
C1988498|Glucose &#x7C; vitreous fluid
C1988484|Glucose &#x7C; Blood cord
C0363662|Glucose [Mass/volume] in Serum or Plasma --3 hours post 100 g glucose PO
C0363662|Glucose^3H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363662|Glucose^3 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363662|Glucose 3h p 100 g Glc PO SerPl-mCnc
C0550363|Glucose 45M p 100 g Glc PO SerPl-mCnc
C0550363|Glucose^45M post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0550363|Glucose [Mass/volume] in Serum or Plasma --45 minutes post 100 g glucose PO
C0550363|Glucose^45M post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942491|Glucose^2.5H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942491|Glucose [Presence] in Urine by Test strip --2.5 hours post dose glucose
C0942491|Glucose^2 1/2 hours post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0942491|Glucose 2.5h p Glc Ur Ql Strip
C0942498|Glucose^6H post dose glucose:MCnc:Pt:Urine:Qn
C0942498|Glucose [Mass/volume] in Urine --6 hours post dose glucose
C0942498|Glucose^6 hours post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C0942498|Glucose 6h p Glc Ur-mCnc
C1148043|Glucose [Moles/volume] in Serum or Plasma --10 minutes post dose glucose
C1148043|Glucose^10M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1148043|Glucose 10M p Glc SerPl-sCnc
C1148043|Glucose^10 minutes post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544048|Glucose [Mass/volume] in Serum or Plasma --4.5 hours post XXX challenge
C1544048|Glucose^4.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544048|Glucose^4.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544048|Glucose 4.5h p chal SerPl-mCnc
C1544145|Glucose [Moles/volume] in Serum or Plasma --15 minutes pre XXX challenge
C1544145|Glucose 15M pre chal SerPl-sCnc
C1544145|Glucose^15M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544145|Glucose^15 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544295|Glucose 30M p Triple Bolus SerPl-sCnc
C1544295|Glucose^30M post dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C1544295|Glucose [Moles/volume] in Serum or Plasma --30 minutes post dose triple bolus
C1544295|Glucose^30 minutes post dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2708582|Glucose 45M p 75 g Glc PO SerPl-sCnc
C2708582|Glucose^45M post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C2708582|Glucose [Moles/volume] in Serum or Plasma --45 minutes post 75 g glucose PO
C2708582|Glucose^45M post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706838|Glucose^45M post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706838|Glucose 45M p OKG SerPl-sCnc
C2706838|Glucose [Moles/volume] in Serum or Plasma --45 minutes post dose ornithine alpha-ketoglutarate
C2706838|Glucose^45M post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598579|Glucose pre betaxolol SerPl-sCnc
C2598579|Glucose [Moles/volume] in Serum or Plasma --pre dose betaxolol
C2598579|Glucose^pre dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598579|Glucose^pre dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484586|Glucose^2H post meal:MCnc:Pt:Bld:Qn
C0484586|Glucose [Mass/volume] in Blood --2 hours post meal
C0484586|Glucose^2 hours post meal:Mass Concentration:Point in time:Whole blood:Quantitative
C0484586|Glucose 2h p meal Bld-mCnc
C0363627|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post 0.05-0.15 U insulin/kg IV 12 hours fasting
C0363627|Glucose^1.5H post 0.05-0.15 U insulin/kg IV post 12H CFst:MCnc:Pt:Ser/Plas:Qn
C0363627|Glucose^1 1/2 hour post 0.05-0.15 U insulin/kg Intravenous post 12 hours Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363627|Glucose 1.5h p U/kg Ins IV SerPl-mCnc
C0799335|Glucose 5 PM SerPl-mCnc
C0799335|Glucose [Mass/volume] in Serum or Plasma --5 PM specimen
C0799335|Glucose^5 PM specimen:MCnc:Pt:Ser/Plas:Qn
C0799335|Glucose^5 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363632|Glucose^10M post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363632|Glucose [Mass/volume] in Serum or Plasma --10 minutes post 0.5 g/kg glucose IV
C0363632|Glucose 10M p .5 g/kg Glc IV SerPl-mCnc
C0363632|Glucose^10 minutes post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0482538|Glucose^pre 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0482538|Glucose [Mass/volume] in Serum or Plasma --pre 0.5 g/kg glucose IV
C0482538|Glucose pre .5 g/kg Glc IV SerPl-mCnc
C0482538|Glucose^pre 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0482542|Glucose pre 75 g Glc PO SerPl-mCnc
C0482542|Glucose^pre 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0482542|Glucose [Mass/volume] in Serum or Plasma --pre 75 g glucose PO
C0482542|Glucose^pre 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363645|Glucose 1M p .5 g/kg Glc IV SerPl-mCnc
C0363645|Glucose^1M post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363645|Glucose [Mass/volume] in Serum or Plasma --1 minute post 0.5 g/kg glucose IV
C0363645|Glucose^1 minute post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363655|Glucose^30M post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363655|Glucose [Mass/volume] in Serum or Plasma --30 minutes post 0.5 g/kg glucose IV
C0363655|Glucose 30M p .5 g/kg Glc IV SerPl-mCnc
C0363655|Glucose^30 minutes post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549993|Glucose sp5 p chal SerPl-mCnc
C0549993|Glucose^5th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549993|Glucose [Mass/volume] in Serum or Plasma --5th specimen post XXX challenge
C0549993|Glucose^5th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0941757|Glucose [Mass/volume] in Urine --1 hour post dose glucose
C0941757|Glucose^1H post dose glucose:MCnc:Pt:Urine:Qn
C0941757|Glucose^1 hour post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C0941757|Glucose 1h p Glc Ur-mCnc
C1316519|Glucose pre/p Arg SerPl-sCnc
C1316519|Glucose^pre or post dose arginine:SCnc:Pt:Ser/Plas:Qn
C1316519|Glucose^pre or post dose arginine:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1316519|Glucose [Moles/volume] in Serum or Plasma --pre or post dose arginine
C1114140|Glucose [Moles/volume] in Serum or Plasma --20 minutes post dose glucose
C1114140|Glucose^20M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114140|Glucose 20M p Glc SerPl-sCnc
C1114140|Glucose^20 minutes post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114882|Glucose [Moles/volume] in Serum or Plasma --1.6 hours post dose glucose
C1114882|Glucose^1.6H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114882|Glucose^1.6 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114882|Glucose 1.6h p Glc SerPl-sCnc
C1544026|Glucose^15.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544026|Glucose [Mass/volume] in Serum or Plasma --15.5 hours post XXX challenge
C1544026|Glucose 15.5h p chal SerPl-mCnc
C1544026|Glucose^15.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542946|Glucose [Moles/volume] in Serum or Plasma --8 minutes post XXX challenge
C1542946|Glucose 8M p chal SerPl-sCnc
C1542946|Glucose^8M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542946|Glucose^8 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542949|Glucose [Moles/volume] in Serum or Plasma --14 minutes post XXX challenge
C1542949|Glucose 14m p chal SerPl-sCnc
C1542949|Glucose^14M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542949|Glucose^14M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2734972|Glucose^2.17H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C2734972|Glucose^2.17H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2734972|Glucose [Mass/volume] in Serum or Plasma --2.17 hours post XXX challenge
C2734972|Glucose 2.17h p chal SerPl-mCnc
C2706812|Glucose [Moles/volume] in Serum or Plasma --15 minutes post dose glucagon
C2706812|Glucose^15M post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706812|Glucose 15M p Gc SerPl-sCnc
C2706812|Glucose^15 minutes post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598586|Glucose^15M pre dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598586|Glucose [Moles/volume] in Serum or Plasma --15 minutes pre dose betaxolol
C2598586|Glucose 15M pre betaxolol SerPl-sCnc
C2598586|Glucose^15 minutes pre dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484579|Glucose^1H post 50 g lactose PO:ACnc:Pt:Urine:Ord:Test strip
C0484579|Glucose [Presence] in Urine by Test strip --1 hour post 50 g lactose PO
C0484579|Glucose^1 hour post 50 g lactose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484579|Glucose 1h p 50 g Lac PO Ur Ql Strip
C0484585|Glucose^2H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484585|Glucose [Presence] in Urine by Test strip --2 hours post 75 g glucose PO
C0484585|Glucose^2 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484585|Glucose 2h p 75 g Glc PO Ur Ql Strip
C0484589|Glucose^30M post 50 g lactose PO:ACnc:Pt:Urine:Ord:Test strip
C0484589|Glucose [Presence] in Urine by Test strip --30 minutes post 50 g lactose PO
C0484589|Glucose 30M p 50 g Lac PO Ur Ql Strip
C0484589|Glucose^30 minutes post 50 g lactose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C1988494|Glucose &#x7C; pleural fluid
C2357654|Glucose &#x7C; Nonbiological fluid
C0363668|Glucose 45M p Ins IV SerPl-mCnc
C0363668|Glucose^45M post dose insulin IV:MCnc:Pt:Ser/Plas:Qn
C0363668|Glucose [Mass/volume] in Serum or Plasma --45 minutes post dose insulin IV
C0363668|Glucose^45M post dose insulin Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363675|Glucose^5M post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363675|Glucose [Mass/volume] in Serum or Plasma --5 minutes post 0.5 g/kg glucose IV
C0363675|Glucose 5M p .5 g/kg Glc IV SerPl-mCnc
C0363675|Glucose^5 minutes post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803252|Glucose^3H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0803252|Glucose [Mass/volume] in Serum or Plasma --3 hours post dose glucose
C0803252|Glucose^3 hours post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803252|Glucose 3h p Glc SerPl-mCnc
C0942624|Glucose [Mass/volume] in Serum or Plasma --7th specimen post XXX challenge
C0942624|Glucose^7th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0942624|Glucose sp7 p chal SerPl-mCnc
C0942624|Glucose^7th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544020|Glucose^9.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544020|Glucose [Mass/volume] in Serum or Plasma --9.5 hours post XXX challenge
C1544020|Glucose^9.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544020|Glucose 9.5h p chal SerPl-mCnc
C1544041|Glucose 12M p chal SerPl-mCnc
C1544041|Glucose [Mass/volume] in Serum or Plasma --12 minutes post XXX challenge
C1544041|Glucose^12M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544041|Glucose^12M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544187|Glucose [Moles/volume] in Serum or Plasma --6 minutes post XXX challenge
C1544187|Glucose^6M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544187|Glucose 6M p chal SerPl-sCnc
C1544187|Glucose^6 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1954697|Glucose 20M pre chal SerPl-mCnc
C1954697|Glucose [Mass/volume] in Serum or Plasma --20 minutes pre XXX challenge
C1954697|Glucose^20M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1954697|Glucose^20 minutes pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0368018|Glucose [Mass/volume] in Urine by Test strip
C0368018|Glucose Ur Strip-mCnc
C0368018|Glucose:MCnc:Pt:Urine:Qn:Test strip
C0368018|Glucose:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C2708621|Glucose^2.5H post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C2708621|Glucose [Moles/volume] in Serum or Plasma --2.5 hours post 75 g glucose PO
C2708621|Glucose^2 1/2 hours post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2708621|Glucose 2.5h p 75 g Glc PO SerPl-sCnc
C0363628|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post 100 g glucose PO
C0363628|Glucose^1.5H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363628|Glucose^1 1/2 hour post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363628|Glucose 1.5h p 100 g Glc PO SerPl-mCnc
C0363667|Glucose [Mass/volume] in Serum or Plasma --40 minutes post 0.5 g/kg glucose IV
C0363667|Glucose 40M p .5 g/kg Glc IV SerPl-mCnc
C0363667|Glucose^40M post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363667|Glucose^40M post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363671|Glucose [Mass/volume] in Serum or Plasma --4 hours post 75 g glucose PO
C0363671|Glucose^4H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363671|Glucose^4 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363671|Glucose 4h p 75 g Glc PO SerPl-mCnc
C0550000|Glucose [Mass/volume] in Serum or Plasma --7 hours post meal
C0550000|Glucose^7H post meal:MCnc:Pt:Ser/Plas:Qn
C0550000|Glucose^7 hours post meal:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0550000|Glucose 7h p meal SerPl-mCnc
C0549970|Glucose^12th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549970|Glucose sp12 p chal SerPl-mCnc
C0549970|Glucose [Mass/volume] in Serum or Plasma --12th specimen post XXX challenge
C0549970|Glucose^12th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0800972|Glucose^post 8H CFst:MCnc:Pt:Ser/Plas:Qn
C0800972|Glucose [Mass/volume] in Serum or Plasma --8 hours fasting
C0800972|Glucose^post 8 hours Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0800972|Glucose p 8h fast SerPl-mCnc
C0942493|Glucose [Mass/volume] in Urine --3 hours post dose glucose
C0942493|Glucose^3H post dose glucose:MCnc:Pt:Urine:Qn
C0942493|Glucose^3 hours post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C0942493|Glucose 3h p Glc Ur-mCnc
C1114209|Glucose^1H post 1.2 g/kg lactose PO:MCnc:Pt:Ser/Plas:Qn
C1114209|Glucose [Mass/volume] in Serum or Plasma --1 hour post 1.2 g/kg lactose PO
C1114209|Glucose^1 hour post 1.2 g/kg lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1114209|Glucose 1h p 1.2 g/kg Lac PO SerPl-mCnc
C1542929|Glucose [Mass/volume] in Serum or Plasma --28 hours post XXX challenge
C1542929|Glucose^28H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1542929|Glucose^28H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542929|Glucose 28h p chal SerPl-mCnc
C1544152|Glucose [Moles/volume] in Serum or Plasma --40 minutes post XXX challenge
C1544152|Glucose 40M p chal SerPl-sCnc
C1544152|Glucose^40M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544152|Glucose^40M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544166|Glucose^14H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544166|Glucose 14h p chal SerPl-sCnc
C1544166|Glucose [Moles/volume] in Serum or Plasma --14 hours post XXX challenge
C1544166|Glucose^14H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544294|Glucose [Moles/volume] in Serum or Plasma --15 minutes post dose triple bolus
C1544294|Glucose 15M p Triple Bolus SerPl-sCnc
C1544294|Glucose^15M post dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C1544294|Glucose^15 minutes post dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1716204|Glucose^8 AM specimen:SCnc:Pt:Ser/Plas:Qn
C1716204|Glucose [Moles/volume] in Serum or Plasma --8 AM specimen
C1716204|Glucose 8 AM SerPl-sCnc
C1716204|Glucose^8 AM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706823|Glucose^15 minutes post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706823|Glucose 15M p Ins IV SerPl-sCnc
C2706823|Glucose^15M post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706823|Glucose [Moles/volume] in Serum or Plasma --15 minutes post dose insulin IV
C2706840|Glucose [Moles/volume] in Serum or Plasma --1.5 hour post dose ornithine alpha-ketoglutarate
C2706840|Glucose^1.5H post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706840|Glucose^1 1/2 hour post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706840|Glucose 1.5h p OKG SerPl-sCnc
C2707121|Glucose sp12 p chal SerPl-sCnc
C2707121|Glucose [Moles/volume] in Serum or Plasma --12th specimen post XXX challenge
C2707121|Glucose^12th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707121|Glucose^12th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2707124|Glucose^4th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707124|Glucose sp4 p chal SerPl-sCnc
C2707124|Glucose [Moles/volume] in Serum or Plasma --4th specimen post XXX challenge
C2707124|Glucose^4th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484596|Glucose [Presence] in Urine by Test strip --5 hours post 75 g glucose PO
C0484596|Glucose^5H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484596|Glucose^5 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484596|Glucose 5h p 75 g Glc PO Ur Ql Strip
C1988482|Glucose &#x7C; blood arterial
C1988486|Glucose &#x7C; body fluid
C1316520|Glucose pre/p CLN SerPl-sCnc
C1316520|Glucose [Moles/volume] in Serum or Plasma --pre or post dose clonidine
C1316520|Glucose^pre or post dose clonidine:SCnc:Pt:Ser/Plas:Qn
C1316520|Glucose^pre or post dose clonidine:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114130|Glucose^3.3H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114130|Glucose [Moles/volume] in Serum or Plasma --3.3 hours post dose glucose
C1114130|Glucose^3.3 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114130|Glucose 3.3h p Glc SerPl-sCnc
C1544235|Glucose [Mass/volume] in Serum or Plasma --10.5 hours post XXX challenge
C1544235|Glucose^10.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544235|Glucose^10.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544235|Glucose 10.5h p chal SerPl-mCnc
C1544199|Glucose [Moles/volume] in Serum or Plasma --2 days post XXX challenge
C1544199|Glucose 2D p chal SerPl-sCnc
C1544199|Glucose^2D post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544199|Glucose^2 days post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1640470|Glucose^3H post dose lactose PO:MCnc:Pt:Urine:Qn
C1640470|Glucose [Mass/volume] in Urine --3 hours post dose lactose PO
C1640470|Glucose^3 hours post dose lactose Oral:Mass Concentration:Point in time:Urine:Quantitative
C1640470|Glucose 3h p Lac PO Ur-mCnc
C2361582|Glucose p meal SerPl-sCnc
C2361582|Glucose^post meal:SCnc:Pt:Ser/Plas:Qn
C2361582|Glucose [Moles/volume] in Serum or Plasma --post meal
C2361582|Glucose^post meal:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706826|Glucose^30 minutes post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706826|Glucose [Moles/volume] in Serum or Plasma --30 minutes post dose insulin IV
C2706826|Glucose^30M post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706826|Glucose 30M p Ins IV SerPl-sCnc
C2598589|Glucose 30M pre betaxolol SerPl-sCnc
C2598589|Glucose [Moles/volume] in Serum or Plasma --30 minutes pre dose betaxolol
C2598589|Glucose^30M pre dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598589|Glucose^30 minutes pre dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484599|Glucose^post 10H CFst:MCnc:Pt:Ser/Plas:Qn
C0484599|Glucose [Mass/volume] in Serum or Plasma --10 hours fasting
C0484599|Glucose^post 10H Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484599|Glucose p 10h fast SerPl-mCnc
C0363665|Glucose^3H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363665|Glucose [Mass/volume] in Serum or Plasma --3 hours post 75 g glucose PO
C0363665|Glucose^3 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363665|Glucose 3h p 75 g Glc PO SerPl-mCnc
C0799333|Glucose^3 PM specimen:MCnc:Pt:Ser/Plas:Qn
C0799333|Glucose 3 PM SerPl-mCnc
C0799333|Glucose [Mass/volume] in Serum or Plasma --3 PM specimen
C0799333|Glucose^3 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0799334|Glucose [Mass/volume] in Serum or Plasma --4 PM specimen
C0799334|Glucose^4 PM specimen:MCnc:Pt:Ser/Plas:Qn
C0799334|Glucose 4 PM SerPl-mCnc
C0799334|Glucose^4 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363670|Glucose [Mass/volume] in Urine --4 hours post 100 g glucose PO
C0363670|Glucose^4H post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363670|Glucose^4 hours post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363670|Glucose 4h p 100 g Glc PO Ur-mCnc
C0797943|Glucose^pre 12H CFst:SCnc:Pt:Ser/Plas:Qn
C0797943|Glucose [Moles/volume] in Serum or Plasma --pre 12 hour fast
C0797943|Glucose^pre 12 hours Calorie fast:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797943|Glucose pre 12h fast SerPl-sCnc
C0944796|Glucose [Mass/volume] in Serum or Plasma --4 hours post XXX challenge
C0944796|Glucose^4H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0944796|Glucose^4 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0944796|Glucose 4h p chal SerPl-mCnc
C0945368|Glucose^3.5H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0945368|Glucose [Presence] in Urine by Test strip --3.5 hours post dose glucose
C0945368|Glucose^3.5 hours post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0945368|Glucose 3.5h p Glc Ur Ql Strip
C0942506|Glucose [Mass/volume] in Serum or Plasma --2.5 hours post dose glucose
C0942506|Glucose^2.5H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0942506|Glucose^2 1/2 hours post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942506|Glucose 2.5h p Glc SerPl-mCnc
C0941759|Glucose^2H post dose glucose:MCnc:Pt:Urine:Qn
C0941759|Glucose [Mass/volume] in Urine --2 hours post dose glucose
C0941759|Glucose^2 hours post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C0941759|Glucose 2h p Glc Ur-mCnc
C1148005|Glucose [Moles/volume] in Serum or Plasma --4 hours post 75 g glucose PO
C1148005|Glucose^4H post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C1148005|Glucose^4 hours post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1148005|Glucose 4h p 75 g Glc PO SerPl-sCnc
C1544148|Glucose 5M p chal SerPl-sCnc
C1544148|Glucose^5M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544148|Glucose [Moles/volume] in Serum or Plasma --5 minutes post XXX challenge
C1544148|Glucose^5 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544157|Glucose [Moles/volume] in Serum or Plasma --3 hours post XXX challenge
C1544157|Glucose^3H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544157|Glucose^3 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544157|Glucose 3h p chal SerPl-sCnc
C1544172|Glucose^19.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544172|Glucose 19.5h p chal SerPl-sCnc
C1544172|Glucose [Moles/volume] in Serum or Plasma --19.5 hours post XXX challenge
C1544172|Glucose^19.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2361848|Glucose [Mass/volume] in Urine by Automated test strip
C2361848|Glucose Ur Strip.auto-mCnc
C2361848|Glucose:MCnc:Pt:Urine:Qn:Test strip.automated
C2361848|Glucose:Mass Concentration:Point in time:Urine:Quantitative:Test strip.automated
C2736395|Glucose^3H post 75 g glucose PO:MCnc:Pt:Urine:Qn
C2736395|Glucose [Mass/volume] in Urine --3 hours post 75 g glucose PO
C2736395|Glucose^3 hours post 75 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C2736395|Glucose 3h p 75 g Glc PO Ur-mCnc
C2736396|Glucose 4sp p Lact SerPl-mCnc
C2736396|Glucose^4th specimen post dose lactose:MCnc:Pt:Ser/Plas:Qn
C2736396|Glucose [Mass/volume] in Serum or Plasma --4th specimen post lactose
C2736396|Glucose^4th specimen post dose lactose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706822|Glucose^2 1/2 hours post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706822|Glucose^2.5H post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706822|Glucose [Moles/volume] in Serum or Plasma --2.5 hours post dose insulin IV
C2706822|Glucose 2.5h p Ins IV SerPl-sCnc
C2924057|Glucose [Molar concentration difference] in Serum or Plasma --3 hours post XXX challenge
C2924057|Glucose^3H post XXX challenge:SCncDiff:Pt:Ser/Plas:Qn
C2924057|Glucose^3 hours post XXX challenge:Difference in Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924057|Glucose 3h p chal SerPl-SCDiff
C2923563|Glucose [Moles/volume] in Serum or Plasma --7 AM specimen
C2923563|Glucose^7 AM specimen:SCnc:Pt:Ser/Plas:Qn
C2923563|Glucose 7 AM SerPl-sCnc
C2923563|Glucose^7 AM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1988492|Glucose &#x7C; pericardial fluid
C0363666|Glucose 3M p .5 g/kg Glc IV SerPl-mCnc
C0363666|Glucose [Mass/volume] in Serum or Plasma --3 minutes post 0.5 g/kg glucose IV
C0363666|Glucose^3M post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363666|Glucose^3 minutes post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363640|Glucose [Mass/volume] in Serum or Plasma --1 hour post 50 g lactose PO
C0363640|Glucose^1H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0363640|Glucose^1 hour post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363640|Glucose 1h p 50 g Lac PO SerPl-mCnc
C0549995|Glucose^6th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549995|Glucose sp6 p chal SerPl-mCnc
C0549995|Glucose [Mass/volume] in Serum or Plasma --6th specimen post XXX challenge
C0549995|Glucose^6th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549969|Glucose [Mass/volume] in Serum or Plasma --12 hours post XXX challenge
C0549969|Glucose^12H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549969|Glucose^12 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549969|Glucose 12h p chal SerPl-mCnc
C0550002|Glucose [Mass/volume] in Serum or Plasma --8 minutes post XXX challenge
C0550002|Glucose 8M p chal SerPl-mCnc
C0550002|Glucose^8M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0550002|Glucose^8 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942492|Glucose 45M p Glc SerPl-mCnc
C0942492|Glucose [Mass/volume] in Serum or Plasma --45 minutes post dose glucose
C0942492|Glucose^45M post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0942492|Glucose^45M post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0941756|Glucose [Moles/volume] in Serum or Plasma --15 minutes post dose glucose
C0941756|Glucose^15M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0941756|Glucose 15M p Glc SerPl-sCnc
C0941756|Glucose^15 minutes post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941760|Glucose [Moles/volume] in Serum or Plasma --2 hours post XXX challenge
C0941760|Glucose^2H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C0941760|Glucose^2 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941760|Glucose 2h p chal SerPl-sCnc
C1316522|Glucose pre/p Glc SerPl-sCnc
C1316522|Glucose^pre or post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1316522|Glucose [Moles/volume] in Serum or Plasma --pre or post dose glucose
C1316522|Glucose^pre or post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114129|Glucose [Moles/volume] in Serum or Plasma --2.6 hours post dose glucose
C1114129|Glucose^2.6H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114129|Glucose^2.6 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114129|Glucose 2.6h p Glc SerPl-sCnc
C1542986|Glucose [Moles/volume] in Serum or Plasma --8 hours post XXX challenge
C1542986|Glucose^8H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542986|Glucose^8 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542986|Glucose 8h p chal SerPl-sCnc
C1544162|Glucose [Moles/volume] in Serum or Plasma --12 hours post XXX challenge
C1544162|Glucose^12H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544162|Glucose^12 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544162|Glucose 12h p chal SerPl-sCnc
C1544176|Glucose [Moles/volume] in Serum or Plasma --22 hours post XXX challenge
C1544176|Glucose^22H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544176|Glucose^22H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544176|Glucose 22h p chal SerPl-sCnc
C1544293|Glucose pre Triple Bolus SerPl-sCnc
C1544293|Glucose [Moles/volume] in Serum or Plasma --pre dose triple bolus
C1544293|Glucose^pre dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C1544293|Glucose^pre dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542952|Glucose^22M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542952|Glucose [Moles/volume] in Serum or Plasma --22 minutes post XXX challenge
C1542952|Glucose 22M p chal SerPl-sCnc
C1542952|Glucose^22M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544193|Glucose^27H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544193|Glucose [Moles/volume] in Serum or Plasma --27 hours post XXX challenge
C1544193|Glucose^27H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544193|Glucose 27h p chal SerPl-sCnc
C1952715|Glucose [Mass/volume] in Serum or Plasma --10 minutes post dose glucose
C1952715|Glucose^10M post dose glucose:MCnc:Pt:Ser/Plas:Qn
C1952715|Glucose 10M p Glc SerPl-mCnc
C1952715|Glucose^10 minutes post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1953181|Glucose^5M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1953181|Glucose 5M p Glc SerPl-sCnc
C1953181|Glucose [Moles/volume] in Serum or Plasma --5 minutes post dose glucose
C1953181|Glucose^5 minutes post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481983|Glucose^40M post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C3481983|Glucose [Moles/volume] in Serum or Plasma --40 minutes post dose lactose PO
C3481983|Glucose^40M post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481983|Glucose 40M p Lac PO SerPl-sCnc
C0484582|Glucose^2.5H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484582|Glucose [Mass/volume] in Serum or Plasma --2.5 hours post 100 g glucose PO
C0484582|Glucose^2 1/2 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484582|Glucose 2.5h p 100 g Glc PO SerPl-mCnc
C0363639|Glucose [Mass/volume] in Urine --1 hour post 50 g glucose PO
C0363639|Glucose^1H post 50 g glucose PO:MCnc:Pt:Urine:Qn
C0363639|Glucose^1 hour post 50 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363639|Glucose 1h p 50 g Glc PO Ur-mCnc
C0482539|Glucose^pre 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0482539|Glucose [Mass/volume] in Serum or Plasma --pre 100 g glucose PO
C0482539|Glucose pre 100 g Glc PO SerPl-mCnc
C0482539|Glucose^pre 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0482543|Glucose [Mass/volume] in Serum or Plasma --pre dose insulin IV
C0482543|Glucose^pre dose insulin IV:MCnc:Pt:Ser/Plas:Qn
C0482543|Glucose pre Ins IV SerPl-mCnc
C0482543|Glucose^pre dose insulin Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0797941|Glucose [Moles/volume] in Serum or Plasma --5 hours post dose glucose
C0797941|Glucose^5H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0797941|Glucose^5 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797941|Glucose 5h p Glc SerPl-sCnc
C0549975|Glucose^15M post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0549975|Glucose 15M p Lac PO SerPl-mCnc
C0549975|Glucose [Mass/volume] in Serum or Plasma --15 minutes post dose lactose PO
C0549975|Glucose^15 minutes post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0944797|Glucose^5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0944797|Glucose [Mass/volume] in Serum or Plasma --5 hours post XXX challenge
C0944797|Glucose^5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0944797|Glucose 5h p chal SerPl-mCnc
C1315291|Glucose [Mass/volume] in Serum or Plasma --45 minutes post dose lactose PO
C1315291|Glucose^45M post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C1315291|Glucose 45M p Lac PO SerPl-mCnc
C1315291|Glucose^45M post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1148003|Glucose^30M post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C1148003|Glucose [Moles/volume] in Serum or Plasma --30 minutes post 75 g glucose PO
C1148003|Glucose 30M p 75 g Glc PO SerPl-sCnc
C1148003|Glucose^30 minutes post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544012|Glucose 15M pre chal SerPl-mCnc
C1544012|Glucose^15M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544012|Glucose [Mass/volume] in Serum or Plasma --15 minutes pre XXX challenge
C1544012|Glucose^15 minutes pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542928|Glucose^27H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1542928|Glucose [Mass/volume] in Serum or Plasma --27 hours post XXX challenge
C1542928|Glucose^27H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542928|Glucose 27h p chal SerPl-mCnc
C1544144|Glucose^30M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544144|Glucose [Moles/volume] in Serum or Plasma --30 minutes pre XXX challenge
C1544144|Glucose 30M pre chal SerPl-sCnc
C1544144|Glucose^30 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542985|Glucose [Moles/volume] in Serum or Plasma --7.5 hours post XXX challenge
C1542985|Glucose^7.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542985|Glucose^7.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542985|Glucose 7.5h p chal SerPl-sCnc
C1542988|Glucose^9H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542988|Glucose [Moles/volume] in Serum or Plasma --9 hours post XXX challenge
C1542988|Glucose^9H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542988|Glucose 9h p chal SerPl-sCnc
C1716223|Glucose^8 PM specimen:SCnc:Pt:Ser/Plas:Qn
C1716223|Glucose [Moles/volume] in Serum or Plasma --8 PM specimen
C1716223|Glucose 8 PM SerPl-sCnc
C1716223|Glucose^8 PM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1642556|Glucose^5H post dose lactose PO:MCnc:Pt:Urine:Qn
C1642556|Glucose [Mass/volume] in Urine --5 hours post dose lactose PO
C1642556|Glucose^5 hours post dose lactose Oral:Mass Concentration:Point in time:Urine:Quantitative
C1642556|Glucose 5h p Lac PO Ur-mCnc
C1979449|Glucose pre/p chal SerPl-sCnc
C1979449|Glucose^pre or post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1979449|Glucose [Moles/volume] in Serum or Plasma --pre or post XXX challenge
C1979449|Glucose^pre or post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2360467|Glucose^2H post dose fructose PO:MCnc:Pt:Ser/Plas:Qn
C2360467|Glucose [Mass/volume] in Serum or Plasma --2 hours post dose fructose PO
C2360467|Glucose^2 hours post dose fructose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2360467|Glucose 2h p fructose PO SerPl-mCnc
C2736397|Glucose [Mass/volume] in Serum or Plasma --5th specimen post lactose
C2736397|Glucose 5sp p Lact SerPl-mCnc
C2736397|Glucose^5th specimen post dose lactose:MCnc:Pt:Ser/Plas:Qn
C2736397|Glucose^5th specimen post dose lactose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706833|Glucose [Moles/volume] in Serum or Plasma --2.5 hour post dose ornithine alpha-ketoglutarate
C2706833|Glucose^2.5H post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706833|Glucose^2 1/2 hours post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706833|Glucose 2.5h p OKG SerPl-sCnc
C1988485|Glucose &#x7C; blood venous
C1988488|Glucose &#x7C; dialysis fluid
C1988493|Glucose &#124; peritoneal fluid
C1988493|Glucose &#x7C; peritoneal fluid
C1988513|Glucose.IV &#x7C; Dose
C0482541|Glucose [Mass/volume] in Serum or Plasma --pre 50 g lactose PO
C0482541|Glucose^pre 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0482541|Glucose pre 50 g Lac PO SerPl-mCnc
C0482541|Glucose^pre 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0802042|Glucose^1H post dose glucose:Imp:Pt:Ser/Plas:Nom
C0802042|Glucose^1 hour post dose glucose:Impression/interpretation of study:Point in time:Serum/Plasma:Nominal
C0802042|Glucose 1h p Glc SerPl-Imp
C0802042|Glucose [Interpretation] in Serum or Plasma--1 hour post dose glucose
C1544019|Glucose^8.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544019|Glucose [Mass/volume] in Serum or Plasma --8.5 hours post XXX challenge
C1544019|Glucose 8.5h p chal SerPl-mCnc
C1544019|Glucose^8.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544023|Glucose 13h p chal SerPl-mCnc
C1544023|Glucose [Mass/volume] in Serum or Plasma --13 hours post XXX challenge
C1544023|Glucose^13H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544023|Glucose^13H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544183|Glucose^3M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544183|Glucose [Moles/volume] in Serum or Plasma --3 minutes pre XXX challenge
C1544183|Glucose 3M pre chal SerPl-sCnc
C1544183|Glucose^3 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544253|Glucose [Moles/volume] in Serum or Plasma --1 hour post dose lactose PO
C1544253|Glucose^1H post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C1544253|Glucose^1 hour post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544253|Glucose 1h p Lac PO SerPl-sCnc
C1716342|Glucose [Mass/volume] in Urine by Test strip --4th specimen post XXX challenge
C1716342|Glucose^4th specimen post XXX challenge:MCnc:Pt:Urine:Qn:Test strip
C1716342|Glucose sp4 p chal Ur Strip-mCnc
C1716342|Glucose^4th specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C1716343|Glucose^5th specimen post XXX challenge:MCnc:Pt:Urine:Qn:Test strip
C1716343|Glucose [Mass/volume] in Urine by Test strip --5th specimen post XXX challenge
C1716343|Glucose sp5 p chal Ur Strip-mCnc
C1716343|Glucose^5th specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C2706825|Glucose [Moles/volume] in Serum or Plasma --3 hours pre dose insulin IV
C2706825|Glucose^3H pre dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706825|Glucose^3 hours pre dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706825|Glucose 3h pre Ins IV SerPl-sCnc
C0484591|Glucose^3H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484591|Glucose [Presence] in Urine by Test strip --3 hours post 75 g glucose PO
C0484591|Glucose^3 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484591|Glucose 3h p 75 g Glc PO Ur Ql Strip
C1988483|Glucose &#x7C; blood capillary
C2357655|Glucose &#x7C; Total parental nutrition
C0363643|Glucose^1H post 75 g glucose PO:MCnc:Pt:Urine:Qn
C0363643|Glucose [Mass/volume] in Urine --1 hour post 75 g glucose PO
C0363643|Glucose^1 hour post 75 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363643|Glucose 1h p 75 g Glc PO Ur-mCnc
C0797931|Glucose [Moles/volume] in Serum or Plasma --2 hours post 100 g glucose PO
C0797931|Glucose^2H post 100 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C0797931|Glucose^2 hours post 100 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797931|Glucose 2h p 100 g Glc PO SerPl-sCnc
C0797932|Glucose [Moles/volume] in Serum or Plasma --2 hours post 50 g lactose PO
C0797932|Glucose^2H post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C0797932|Glucose^2 hours post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797932|Glucose 2h p 50 g Lac PO SerPl-sCnc
C0549981|Glucose^2H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549981|Glucose [Mass/volume] in Serum or Plasma --2 hours post XXX challenge
C0549981|Glucose^2 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549981|Glucose 2h p chal SerPl-mCnc
C0942499|Glucose^1H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942499|Glucose [Presence] in Urine by Test strip --1 hour post dose glucose
C0942499|Glucose^1 hour post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0942499|Glucose 1h p Glc Ur Ql Strip
C0941770|Glucose^1.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C0941770|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post XXX challenge
C0941770|Glucose^1 1/2 hour post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941770|Glucose 1.5h p chal SerPl-sCnc
C1544011|Glucose^30M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544011|Glucose [Mass/volume] in Serum or Plasma --30 minutes pre XXX challenge
C1544011|Glucose 30M pre chal SerPl-mCnc
C1544011|Glucose^30 minutes pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544167|Glucose^15.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544167|Glucose 15.5h p chal SerPl-sCnc
C1544167|Glucose [Moles/volume] in Serum or Plasma --15.5 hours post XXX challenge
C1544167|Glucose^15.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544169|Glucose^17.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544169|Glucose [Moles/volume] in Serum or Plasma --17.5 hours post XXX challenge
C1544169|Glucose 17.5h p chal SerPl-sCnc
C1544169|Glucose^17.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1716203|Glucose 12 AM SerPl-sCnc
C1716203|Glucose^12 AM specimen:SCnc:Pt:Ser/Plas:Qn
C1716203|Glucose [Moles/volume] in Serum or Plasma --12 AM specimen
C1716203|Glucose^12 AM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1716205|Glucose^12 PM specimen:SCnc:Pt:Ser/Plas:Qn
C1716205|Glucose 12 PM SerPl-sCnc
C1716205|Glucose [Moles/volume] in Serum or Plasma --12 PM specimen
C1716205|Glucose^12 PM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706816|Glucose 4M p Gc SerPl-sCnc
C2706816|Glucose [Moles/volume] in Serum or Plasma --4 minutes post dose glucagon
C2706816|Glucose^4M post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706816|Glucose^4 minutes post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706830|Glucose^1.5H post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706830|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post dose insulin IV
C2706830|Glucose^1 1/2 hour post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706830|Glucose 1.5h p Ins IV SerPl-sCnc
C2706835|Glucose [Moles/volume] in Serum or Plasma --15 minutes pre dose ornithine alpha-ketoglutarate
C2706835|Glucose^15M pre dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706835|Glucose 15M pre OKG SerPl-sCnc
C2706835|Glucose^15 minutes pre dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598076|Glucose [Mass/volume] in Serum or Plasma --40 minutes post 50 g lactose PO
C2598076|Glucose^40M post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C2598076|Glucose 40M p 50 g lac PO SerPl-mCnc
C2598076|Glucose^40M post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2924056|Glucose [Molar concentration difference] in Serum or Plasma --2 hours post XXX challenge
C2924056|Glucose^2H post XXX challenge:SCncDiff:Pt:Ser/Plas:Qn
C2924056|Glucose^2 hours post XXX challenge:Difference in Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924056|Glucose 2h p chal SerPl-SCDiff
C0363638|Glucose [Mass/volume] in Serum or Plasma --1 hour post 50 g glucose PO
C0363638|Glucose^1H post 50 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363638|Glucose^1 hour post 50 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363638|Glucose 1h p 50 g Glc PO SerPl-mCnc
C0482540|Glucose^pre 12H CFst:MCnc:Pt:Ser/Plas:Qn
C0482540|Glucose [Mass/volume] in Serum or Plasma --pre 12 hour fast
C0482540|Glucose^pre 12 hours Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0482540|Glucose pre 12h fast SerPl-mCnc
C0797927|Glucose^1H post 100 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C0797927|Glucose [Moles/volume] in Serum or Plasma --1 hour post 100 g glucose PO
C0797927|Glucose^1 hour post 100 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797927|Glucose 1h p 100 g Glc PO SerPl-sCnc
C0797933|Glucose [Moles/volume] in Serum or Plasma --2 hours post dose glucose
C0797933|Glucose^2H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0797933|Glucose^2 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797933|Glucose 2h p Glc SerPl-sCnc
C0947224|Glucose 30M p Lac PO SerPl-mCnc
C0947224|Glucose [Mass/volume] in Serum or Plasma --30 minutes post dose lactose PO
C0947224|Glucose^30M post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0947224|Glucose^30 minutes post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0941768|Glucose^5.5H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0941768|Glucose [Moles/volume] in Serum or Plasma --5.5 hours post dose glucose
C0941768|Glucose^5.5 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941768|Glucose 5.5h p Glc SerPl-sCnc
C1542982|Glucose^6H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542982|Glucose [Moles/volume] in Serum or Plasma --6 hours post XXX challenge
C1542982|Glucose^6 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542982|Glucose 6h p chal SerPl-sCnc
C1544255|Glucose [Moles/volume] in Serum or Plasma --2 hours post dose lactose PO
C1544255|Glucose^2H post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C1544255|Glucose^2 hours post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544255|Glucose 2h p Lac PO SerPl-sCnc
C1543636|Glucose [Mass/volume] in Serum or Plasma --1st specimen post dose lactose
C1543636|Glucose^1st specimen post dose lactose:MCnc:Pt:Ser/Plas:Qn
C1543636|Glucose sp1 p Lac SerPl-mCnc
C1543636|Glucose^1st specimen post dose lactose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1716341|Glucose sp3 p chal Ur Strip-mCnc
C1716341|Glucose [Mass/volume] in Urine by Test strip --3rd specimen post XXX challenge
C1716341|Glucose^3rd specimen post XXX challenge:MCnc:Pt:Urine:Qn:Test strip
C1716341|Glucose^3rd specimen post XXX challenge:Mass Concentration:Point in time:Urine:Quantitative:Test strip
C1952717|Glucose [Mass/volume] in Serum or Plasma --8 AM specimen
C1952717|Glucose^8 AM specimen:MCnc:Pt:Ser/Plas:Qn
C1952717|Glucose 8 AM SerPl-mCnc
C1952717|Glucose^8 AM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706814|Glucose 20M p Gc SerPl-sCnc
C2706814|Glucose^20M post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706814|Glucose [Moles/volume] in Serum or Plasma --20 minutes post dose glucagon
C2706814|Glucose^20 minutes post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706829|Glucose^1.3H post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706829|Glucose [Moles/volume] in Serum or Plasma --1.3 hours post dose insulin IV
C2706829|Glucose^1.3 hours post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706829|Glucose 1.3h p Ins IV SerPl-sCnc
C2706832|Glucose [Moles/volume] in Serum or Plasma --2 hour post dose ornithine alpha-ketoglutarate
C2706832|Glucose^2H post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706832|Glucose^2 hours post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706832|Glucose 2h p OKG SerPl-sCnc
C2598075|Glucose^20M post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C2598075|Glucose [Mass/volume] in Serum or Plasma --20 minutes post 50 g lactose PO
C2598075|Glucose 20M p 50 g lac PO SerPl-mCnc
C2598075|Glucose^20 minutes post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2598580|Glucose^2H post dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598580|Glucose [Moles/volume] in Serum or Plasma --2 hours post dose betaxolol
C2598580|Glucose^2 hours post dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598580|Glucose 2h p betaxolol SerPl-sCnc
C0484597|Glucose [Mass/volume] in Serum or Plasma --6 hours post 75 g glucose PO
C0484597|Glucose^6H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484597|Glucose^6 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484597|Glucose 6h p 75 g Glc PO SerPl-mCnc
C0484600|Glucose^post CFst:ACnc:Pt:Urine:Ord:Test strip
C0484600|Fasting glucose [Presence] in Urine by Test strip
C0484600|Glucose p fast Ur Ql Strip
C0484600|Glucose^post Calorie fast:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0800042|Glucose [Presence] in Urine --5th specimen post XXX challenge
C0800042|Glucose^5th specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800042|Glucose sp5 p chal Ur Ql
C0800042|Glucose^5th specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0363634|Glucose^1H post 0.05-0.15 U insulin/kg IV post 12H CFst:MCnc:Pt:Ser/Plas:Qn
C0363634|Glucose [Mass/volume] in Serum or Plasma --1 hour post 0.05-0.15 U insulin/kg IV post 12H CFst
C0363634|Glucose^1 hour post 0.05-0.15 U insulin/kg Intravenous post 12 hours Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363634|Glucose 1h p U/kg Ins IV SerPl-mCnc
C0363677|Glucose^6H post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363677|Glucose [Mass/volume] in Urine --6 hours post 100 g glucose PO
C0363677|Glucose^6 hours post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363677|Glucose 6h p 100 g Glc PO Ur-mCnc
C0363651|Glucose^2H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363651|Glucose [Mass/volume] in Serum or Plasma --2 hours post 75 g glucose PO
C0363651|Glucose^2 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363651|Glucose 2h p 75 g Glc PO SerPl-mCnc
C0550005|Glucose [Mass/volume] in Serum or Plasma --9th specimen post XXX challenge
C0550005|Glucose^9th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0550005|Glucose sp9 p chal SerPl-mCnc
C0550005|Glucose^9th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549968|Glucose sp11 p chal SerPl-mCnc
C0549968|Glucose^11th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549968|Glucose [Mass/volume] in Serum or Plasma --11th specimen post XXX challenge
C0549968|Glucose^11th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544032|Glucose 20H p chal SerPl-mCnc
C1544032|Glucose^20H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544032|Glucose [Mass/volume] in Serum or Plasma --20 hours post XXX challenge
C1544032|Glucose^20H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542983|Glucose^6.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542983|Glucose [Moles/volume] in Serum or Plasma --6.5 hours post XXX challenge
C1542983|Glucose^6.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542983|Glucose 6.5h p chal SerPl-sCnc
C1544164|Glucose 13h p chal SerPl-sCnc
C1544164|Glucose [Moles/volume] in Serum or Plasma --13 hours post XXX challenge
C1544164|Glucose^13H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544164|Glucose^13H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544171|Glucose [Moles/volume] in Serum or Plasma --18.5 hours post XXX challenge
C1544171|Glucose^18.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544171|Glucose 18.5h p chal SerPl-sCnc
C1544171|Glucose^18.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544182|Glucose 8M pre chal SerPl-sCnc
C1544182|Glucose^8M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544182|Glucose [Moles/volume] in Serum or Plasma --8 minutes pre XXX challenge
C1544182|Glucose^8 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542950|Glucose^16M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542950|Glucose 16m p chal SerPl-sCnc
C1542950|Glucose [Moles/volume] in Serum or Plasma --16 minutes post XXX challenge
C1542950|Glucose^16M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542953|Glucose [Moles/volume] in Serum or Plasma --25 minutes post XXX challenge
C1542953|Glucose^25M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542953|Glucose 25M p chal SerPl-sCnc
C1542953|Glucose^25 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544190|Glucose [Moles/volume] in Serum or Plasma --5.5 hours post XXX challenge
C1544190|Glucose^5.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544190|Glucose^5.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544190|Glucose 5.5h p chal SerPl-sCnc
C1543638|Glucose sp3 p Lac SerPl-mCnc
C1543638|Glucose [Mass/volume] in Serum or Plasma --3rd specimen post dose lactose
C1543638|Glucose^3rd specimen post dose lactose:MCnc:Pt:Ser/Plas:Qn
C1543638|Glucose^3rd specimen post dose lactose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1716427|Glucose [Moles/volume] in Serum or Plasma --2.5 hours post 50 g lactose PO
C1716427|Glucose^2.5H post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C1716427|Glucose^2 1/2 hours post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1716427|Glucose 2.5h p 50 g Lac PO SerPl-sCnc
C1716125|Glucose^1.5H post meal:SCnc:Pt:Ser/Plas:Qn
C1716125|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post meal
C1716125|Glucose^1 1/2 hour post meal:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1716125|Glucose 1.5h p meal SerPl-sCnc
C1978755|Glucose^15M post 0.1 U/kg insulin:MCnc:Pt:Ser/Plas:Qn
C1978755|Glucose 15M p 0.1 U/kg Ins SerPl-mCnc
C1978755|Glucose [Mass/volume] in Serum or Plasma --15 minutes post 0.1 U/kg insulin
C1978755|Glucose^15 minutes post 0.1 U/kg insulin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706834|Glucose^15M post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706834|Glucose [Moles/volume] in Serum or Plasma --15 minutes post dose ornithine alpha-ketoglutarate
C2706834|Glucose 15M p OKG SerPl-sCnc
C2706834|Glucose^15 minutes post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924055|Glucose^1.5H post XXX challenge:SCncDiff:Pt:Ser/Plas:Qn
C2924055|Glucose [Molar concentration difference] in Serum or Plasma --1.5 hours post XXX challenge
C2924055|Glucose^1 1/2 hour post XXX challenge:Difference in Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924055|Glucose 1.5h p chal SerPl-SCDiff
C3699463|Glucose [Moles/volume] in Serum or Plasma --15 minutes post 50 g lactose PO
C3699463|Glucose 15M p 50 g Lac PO SerPl-sCnc
C3699463|Glucose^15 minutes post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3699463|Glucose^15M post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C0484595|Glucose [Mass/volume] in Serum or Plasma --5.5 hours post 100 g glucose PO
C0484595|Glucose^5.5H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484595|Glucose^5.5 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484595|Glucose 5.5h p 100 g Glc PO SerPl-mCnc
C1988480|Glucose &#x7C; amniotic fluid
C0800045|Glucose^8th specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800045|Glucose [Presence] in Urine --8th specimen post XXX challenge
C0800045|Glucose sp8 p chal Ur Ql
C0800045|Glucose^8th specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0363686|Glucose [Mass/volume] in Urine --12 hours fasting
C0363686|Glucose^post 12H CFst:MCnc:Pt:Urine:Qn
C0363686|Glucose^post 12 hours Calorie fast:Mass Concentration:Point in time:Urine:Quantitative
C0363686|Glucose p 12h fast Ur-mCnc
C0482536|Glucose^30M post 0.1 U/kg insulin:MCnc:Pt:Ser/Plas:Qn
C0482536|Glucose 30M p 0.1 U/kg Ins SerPl-mCnc
C0482536|Glucose [Mass/volume] in Serum or Plasma --30 minutes post 0.1 U/kg insulin
C0482536|Glucose^30 minutes post 0.1 U/kg insulin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549977|Glucose^1H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549977|Glucose [Mass/volume] in Serum or Plasma --1 hour post XXX challenge
C0549977|Glucose^1 hour post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549977|Glucose 1h p chal SerPl-mCnc
C0549998|Glucose 70M p chal SerPl-mCnc
C0549998|Glucose^70M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549998|Glucose [Mass/volume] in Serum or Plasma --70 minutes post XXX challenge
C0549998|Glucose^70M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803256|Glucose^post 50 g glucose:MCnc:Pt:Ser/Plas:Qn
C0803256|Glucose p 50 g Glc SerPl-mCnc
C0803256|Glucose [Mass/volume] in Serum or Plasma --post 50 g glucose
C0803256|Glucose^post 50 g glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0941761|Glucose^3.5H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0941761|Glucose [Moles/volume] in Serum or Plasma --3.5 hours post dose glucose
C0941761|Glucose^3.5 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941761|Glucose 3.5h p Glc SerPl-sCnc
C1316523|Glucose pre/p Ins SerPl-sCnc
C1316523|Glucose [Moles/volume] in Serum or Plasma --pre or post dose insulin
C1316523|Glucose^pre or post dose insulin:SCnc:Pt:Ser/Plas:Qn
C1316523|Glucose^pre or post dose insulin:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114141|Glucose^1.3H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114141|Glucose [Moles/volume] in Serum or Plasma --1.3 hours post dose glucose
C1114141|Glucose^1.3 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114141|Glucose 1.3h p Glc SerPl-sCnc
C1114142|Glucose^2.3H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114142|Glucose [Moles/volume] in Serum or Plasma --2.3 hours post dose glucose
C1114142|Glucose^2.3 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1114142|Glucose 2.3h p Glc SerPl-sCnc
C1114210|Glucose [Mass/volume] in Serum or Plasma --2 hours post 1.2 g/kg lactose PO
C1114210|Glucose^2H post 1.2 g/kg lactose PO:MCnc:Pt:Ser/Plas:Qn
C1114210|Glucose^2 hours post 1.2 g/kg lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1114210|Glucose 2h p 1.2 g/kg Lac PO SerPl-mCnc
C1544037|Glucose^1D post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544037|Glucose [Mass/volume] in Serum or Plasma --1 day post XXX challenge
C1544037|Glucose 1D p chal SerPl-mCnc
C1544037|Glucose^1 day post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544168|Glucose 16h p chal SerPl-sCnc
C1544168|Glucose^16H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544168|Glucose [Moles/volume] in Serum or Plasma --16 hours post XXX challenge
C1544168|Glucose^16H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544181|Glucose [Moles/volume] in Serum or Plasma --13 minutes pre XXX challenge
C1544181|Glucose 13m pre chal SerPl-sCnc
C1544181|Glucose^13M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544181|Glucose^13M pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544813|Glucose BS BldC-mCnc
C1544813|Glucose^baseline:MCnc:Pt:BldC:Qn
C1544813|Glucose [Mass/volume] in Capillary blood --baseline
C1544813|Glucose^baseline:Mass Concentration:Point in time:Blood capillary:Quantitative
C1952720|Glucose 12 PM SerPl-mCnc
C1952720|Glucose^12 PM specimen:MCnc:Pt:Ser/Plas:Qn
C1952720|Glucose [Mass/volume] in Serum or Plasma --12 PM specimen
C1952720|Glucose^12 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2708581|Glucose^1.5H post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C2708581|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post 75 g glucose PO
C2708581|Glucose^1 1/2 hour post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2708581|Glucose 1.5h p 75 g Glc PO SerPl-sCnc
C2598592|Glucose^1.5H post dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598592|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post dose betaxolol
C2598592|Glucose^1 1/2 hour post dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598592|Glucose 1.5h p betaxolol SerPl-sCnc
C2707120|Glucose^11th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707120|Glucose [Moles/volume] in Serum or Plasma --11th specimen post XXX challenge
C2707120|Glucose sp11 p chal SerPl-sCnc
C2707120|Glucose^11th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484577|Glucose^1.5H post 50 g lactose PO:ACnc:Pt:Urine:Ord:Test strip
C0484577|Glucose [Presence] in Urine by Test strip --1.5 hours post 50 g lactose PO
C0484577|Glucose^1 1/2 hour post 50 g lactose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484577|Glucose 1.5h p 50 g Lac PO Ur Ql Strip
C3655027|Glucose [Moles/volume] in Serum or Plasma --15 minutes post dose lactose PO
C3655027|Glucose 15M p Lac PO SerPl-sCnc
C3655027|Glucose^15M post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C3655027|Glucose^15 minutes post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1988496|Glucose &#x7C; synovial fluid
C0800043|Glucose sp6 p chal Ur Ql
C0800043|Glucose [Presence] in Urine --6th specimen post XXX challenge
C0800043|Glucose^6th specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800043|Glucose^6th specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0700436|Glucose [Mass/volume] in Serum or Plasma --6 hours post 100 g glucose PO
C0700436|Glucose^6H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0700436|Glucose^6 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0700436|Glucose 6h p 100 g Glc PO SerPl-mCnc
C0482544|Glucose [Mass/volume] in Serum or Plasma --post CFst
C0482544|Glucose^post CFst:MCnc:Pt:Ser/Plas:Qn
C0482544|Fasting glucose [Mass/volume] in Serum or Plasma
C0482544|Glucose p fast SerPl-mCnc
C0482544|Glucose^post Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549985|Glucose [Mass/volume] in Serum or Plasma --3.5 hours post dose lactose PO
C0549985|Glucose^3.5H post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0549985|Glucose^3.5 hours post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549985|Glucose 3.5h p Lac PO SerPl-mCnc
C0803255|Glucose^1.5H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0803255|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post dose glucose
C0803255|Glucose^1 1/2 hour post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803255|Glucose 1.5h p Glc SerPl-mCnc
C0801395|Glucose^6H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0801395|Glucose [Mass/volume] in Serum or Plasma --6 hours post 50 g lactose PO
C0801395|Glucose^6 hours post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0801395|Glucose 6h p 50 g Lac PO SerPl-mCnc
C0942494|Glucose^4H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0942494|Glucose [Mass/volume] in Serum or Plasma --4 hours post dose glucose
C0942494|Glucose^4 hours post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942494|Glucose 4h p Glc SerPl-mCnc
C0942504|Glucose [Presence] in Urine by Test strip --5 hours post dose glucose
C0942504|Glucose^5H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942504|Glucose^5 hours post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0942504|Glucose 5h p Glc Ur Ql Strip
C0945369|Glucose [Presence] in Urine by Test strip --1.5 hours post dose glucose
C0945369|Glucose^1.5H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0945369|Glucose^1 1/2 hour post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0945369|Glucose 1.5h p Glc Ur Ql Strip
C0945253|Glucose^1.5H post dose glucose:MCnc:Pt:Urine:Qn
C0945253|Glucose [Mass/volume] in Urine --1.5 hours post dose glucose
C0945253|Glucose^1 1/2 hour post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C0945253|Glucose 1.5h p Glc Ur-mCnc
C2607838|Glucose [Mass or Molecules/volume] in Serum or Plasma --post CFst
C2607838|Glucose p fast SerPl-msCnc
C2607838|Glucose^post CFst:MSCnc:Pt:Ser/Plas:Qn
C2607838|Fasting glucose [Mass or Moles/volume] in Serum or Plasma
C2607838|Glucose^post Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544016|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post XXX challenge
C1544016|Glucose^1.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544016|Glucose^1 1/2 hour post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544016|Glucose 1.5h p chal SerPl-mCnc
C1542981|Glucose [Moles/volume] in Serum or Plasma --5 hours post XXX challenge
C1542981|Glucose^5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542981|Glucose^5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542981|Glucose 5h p chal SerPl-sCnc
C1544175|Glucose [Moles/volume] in Serum or Plasma --21.5 hours post XXX challenge
C1544175|Glucose^21.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544175|Glucose^21.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544175|Glucose 21.5h p chal SerPl-sCnc
C1544297|Glucose^1H post dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C1544297|Glucose [Moles/volume] in Serum or Plasma --1 hour post dose triple bolus
C1544297|Glucose^1 hour post dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544297|Glucose 1h p Triple Bolus SerPl-sCnc
C1542948|Glucose [Moles/volume] in Serum or Plasma --12 minutes post XXX challenge
C1542948|Glucose^12M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542948|Glucose 12M p chal SerPl-sCnc
C1542948|Glucose^12M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544192|Glucose^26H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544192|Glucose [Moles/volume] in Serum or Plasma --26 hours post XXX challenge
C1544192|Glucose^26H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544192|Glucose 26h p chal SerPl-sCnc
C1641496|Glucose^4H post dose lactose PO:MCnc:Pt:Urine:Qn
C1641496|Glucose [Mass/volume] in Urine --4 hours post dose lactose PO
C1641496|Glucose^4 hours post dose lactose Oral:Mass Concentration:Point in time:Urine:Quantitative
C1641496|Glucose 4h p Lac PO Ur-mCnc
C2361581|Glucose p chal SerPl-sCnc
C2361581|Glucose^post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2361581|Glucose [Moles/volume] in Serum or Plasma --post XXX challenge
C2361581|Glucose^post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1952721|Glucose [Mass/volume] in Serum or Plasma --6 PM specimen
C1952721|Glucose^6 PM specimen:MCnc:Pt:Ser/Plas:Qn
C1952721|Glucose 6 PM SerPl-mCnc
C1952721|Glucose^6 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954699|Glucose^12 AM specimen:MCnc:Pt:Ser/Plas:Qn
C1954699|Glucose [Mass/volume] in Serum or Plasma --12 AM specimen
C1954699|Glucose 12 AM SerPl-mCnc
C1954699|Glucose^12 AM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706819|Glucose 8M p Gc SerPl-sCnc
C2706819|Glucose^8M post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706819|Glucose [Moles/volume] in Serum or Plasma --8 minutes post dose glucagon
C2706819|Glucose^8 minutes post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706827|Glucose^45M post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706827|Glucose^45M post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706827|Glucose [Moles/volume] in Serum or Plasma --45 minutes post dose insulin IV
C2706827|Glucose 45M p Ins IV SerPl-sCnc
C2598578|Glucose [Moles/volume] in Serum or Plasma --4 AM specimen
C2598578|Glucose^4 AM specimen:SCnc:Pt:Ser/Plas:Qn
C2598578|Glucose 4 AM specimen SerPl-sCnc
C2598578|Glucose^4 AM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481984|Glucose [Moles/volume] in Serum or Plasma --20 minutes post 50 g lactose PO
C3481984|Glucose^20 minutes post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481984|Glucose^20M post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C3481984|Glucose 20M p 50 g lac PO SerPl-sCnc
C3533247|Glucose.serum-glucose.plr fld
C0484587|Glucose^3.5H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484587|Glucose [Mass/volume] in Serum or Plasma --3.5 hours post 100 g glucose PO
C0484587|Glucose^3.5 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484587|Glucose 3.5h p 100 g Glc PO SerPl-mCnc
C0799332|Glucose 2 PM SerPl-mCnc
C0799332|Glucose [Mass/volume] in Serum or Plasma --2 PM specimen
C0799332|Glucose^2 PM specimen:MCnc:Pt:Ser/Plas:Qn
C0799332|Glucose^2 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363674|Glucose^5H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363674|Glucose [Mass/volume] in Serum or Plasma --5 hours post 75 g glucose PO
C0363674|Glucose^5 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363674|Glucose 5h p 75 g Glc PO SerPl-mCnc
C0363685|Glucose [Mass/volume] in Serum or Plasma --12 hours fasting
C0363685|Glucose^post 12H CFst:MCnc:Pt:Ser/Plas:Qn
C0363685|Glucose^post 12 hours Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363685|Glucose p 12h fast SerPl-mCnc
C0797934|Glucose^2H post meal:SCnc:Pt:BldC:Qn
C0797934|Glucose [Moles/volume] in Capillary blood --2 hours post meal
C0797934|Glucose^2 hours post meal:Substance Concentration:Point in time:Blood capillary:Quantitative
C0797934|Glucose 2h p meal BldC-sCnc
C0797945|Fasting glucose [Moles/volume] in Serum or Plasma
C0797945|Glucose^post CFst:SCnc:Pt:Ser/Plas:Qn
C0797945|Glucose p fast SerPl-sCnc
C0797945|Glucose^post Calorie fast:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0549999|Glucose^7H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549999|Glucose [Mass/volume] in Serum or Plasma --7 hours post XXX challenge
C0549999|Glucose^7 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549999|Glucose 7h p chal SerPl-mCnc
C0549990|Glucose [Mass/volume] in Serum or Plasma --4 minutes post XXX challenge
C0549990|Glucose^4M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549990|Glucose 4M p chal SerPl-mCnc
C0549990|Glucose^4 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803253|Glucose [Mass/volume] in Serum or Plasma --1 hour post dose glucose
C0803253|Glucose^1H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0803253|Glucose^1 hour post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803253|Glucose 1h p Glc SerPl-mCnc
C0801384|Glucose^3H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0801384|Glucose [Mass/volume] in Serum or Plasma --3 hours post XXX challenge
C0801384|Glucose^3 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0801384|Glucose 3h p chal SerPl-mCnc
C0947266|Glucose^3.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0947266|Glucose [Mass/volume] in Serum or Plasma --3.5 hours post XXX challenge
C0947266|Glucose^3.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0947266|Glucose 3.5h p chal SerPl-mCnc
C0941762|Glucose [Mass/volume] in Urine --30 minutes post dose glucose
C0941762|Glucose 30M p Glc Ur-mCnc
C0941762|Glucose^30M post dose glucose:MCnc:Pt:Urine:Qn
C0941762|Glucose^30 minutes post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C1544034|Glucose [Mass/volume] in Serum or Plasma --21.5 hours post XXX challenge
C1544034|Glucose^21.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544034|Glucose^21.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544034|Glucose 21.5h p chal SerPl-mCnc
C1544044|Glucose^19M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544044|Glucose [Mass/volume] in Serum or Plasma --19 minutes post XXX challenge
C1544044|Glucose 19M p chal SerPl-mCnc
C1544044|Glucose^19M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544160|Glucose [Moles/volume] in Serum or Plasma --10.75 hours post XXX challenge
C1544160|Glucose 10.75h p chal SerPl-sCnc
C1544160|Glucose^10.75H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544160|Glucose^10.75H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544174|Glucose^20.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544174|Glucose [Moles/volume] in Serum or Plasma --20.5 hours post XXX challenge
C1544174|Glucose^20.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544174|Glucose 20.5h p chal SerPl-sCnc
C1544237|Glucose 13m pre chal SerPl-mCnc
C1544237|Glucose^13M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544237|Glucose [Mass/volume] in Serum or Plasma --13 minutes pre XXX challenge
C1544237|Glucose^13M pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706828|Glucose^1 hour post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706828|Glucose^1H post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706828|Glucose [Moles/volume] in Serum or Plasma --1 hour post dose insulin IV
C2706828|Glucose 1h p Ins IV SerPl-sCnc
C2598588|Glucose [Moles/volume] in Serum or Plasma --30 minutes post dose betaxolol
C2598588|Glucose 30M p betaxolol SerPl-sCnc
C2598588|Glucose^30M post dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598588|Glucose^30 minutes post dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924054|Glucose^1H post XXX challenge:SCncDiff:Pt:Ser/Plas:Qn
C2924054|Glucose [Molar concentration difference] in Serum or Plasma --1 hour post XXX challenge
C2924054|Glucose^1 hour post XXX challenge:Difference in Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924054|Glucose 1h p chal SerPl-SCDiff
C2923561|Glucose^11 AM specimen:SCnc:Pt:Ser/Plas:Qn
C2923561|Glucose [Moles/volume] in Serum or Plasma --11 AM specimen
C2923561|Glucose 11 AM SerPl-sCnc
C2923561|Glucose^11 AM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2970600|Glucose^baseline:MCnc:Pt:Dial fld prt:Qn
C2970600|Glucose BS DiafP-mCnc
C2970600|Glucose [Mass/volume] in Peritoneal dialysis fluid --baseline
C2970600|Glucose^baseline:Mass Concentration:Point in time:Peritoneal dialysis fluid:Quantitative
C1988481|Glucose &#x7C; bld-ser-plas
C1988490|Glucose &#x7C; gastric fluid
C0482534|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post 75 g glucose PO
C0482534|Glucose^1.5H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0482534|Glucose^1 1/2 hour post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0482534|Glucose 1.5h p 75 g Glc PO SerPl-mCnc
C0363646|Glucose^20M post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363646|Glucose [Mass/volume] in Serum or Plasma --20 minutes post 0.5 g/kg glucose IV
C0363646|Glucose 20M p .5 g/kg Glc IV SerPl-mCnc
C0363646|Glucose^20 minutes post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942500|Glucose^2H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942500|Glucose [Presence] in Urine by Test strip --2 hours post dose glucose
C0942500|Glucose^2 hours post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0942500|Glucose 2h p Glc Ur Ql Strip
C0942723|Glucose [Mass/volume] in Serum or Plasma --11 hour post XXX challenge
C0942723|Glucose^11H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0942723|Glucose^11H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942723|Glucose 11h p chal SerPl-mCnc
C0941767|Glucose^4H post dose glucose:MCnc:Pt:Urine:Qn
C0941767|Glucose [Mass/volume] in Urine --4 hours post dose glucose
C0941767|Glucose^4 hours post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C0941767|Glucose 4h p Glc Ur-mCnc
C1315495|Glucose [Mass/volume] in Serum or Plasma --30 minutes post 1.2 g/kg lactose PO
C1315495|Glucose^30M post 1.2 g/kg lactose PO:MCnc:Pt:Ser/Plas:Qn
C1315495|Glucose 30M p 1.2 g/kg Lac PO SerPl-mCnc
C1315495|Glucose^30 minutes post 1.2 g/kg lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1114881|Glucose^40M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1114881|Glucose [Moles/volume] in Serum or Plasma --40 minutes post dose glucose
C1114881|Glucose 40M p Glc SerPl-sCnc
C1114881|Glucose^40M post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544017|Glucose [Mass/volume] in Serum or Plasma --100 minutes post XXX challenge
C1544017|Glucose^100M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544017|Glucose 100M p chal SerPl-mCnc
C1544017|Glucose^100M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544018|Glucose^110M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544018|Glucose [Mass/volume] in Serum or Plasma --110 minutes post XXX challenge
C1544018|Glucose 110m p chal SerPl-mCnc
C1544018|Glucose^110M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544185|Glucose 3M p chal SerPl-sCnc
C1544185|Glucose^3M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544185|Glucose [Moles/volume] in Serum or Plasma --3 minutes post XXX challenge
C1544185|Glucose^3 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544186|Glucose 4M p chal SerPl-sCnc
C1544186|Glucose^4M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544186|Glucose [Moles/volume] in Serum or Plasma --4 minutes post XXX challenge
C1544186|Glucose^4 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1641493|Glucose [Mass/volume] in Urine --1 hour post dose lactose PO
C1641493|Glucose^1H post dose lactose PO:MCnc:Pt:Urine:Qn
C1641493|Glucose^1 hour post dose lactose Oral:Mass Concentration:Point in time:Urine:Quantitative
C1641493|Glucose 1h p Lac PO Ur-mCnc
C0484583|Glucose^2.5H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484583|Glucose [Mass/volume] in Serum or Plasma --2.5 hours post 75 g glucose PO
C0484583|Glucose^2 1/2 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484583|Glucose 2.5h p 75 g Glc PO SerPl-mCnc
C1988487|Glucose &#x7C; cerebral spinal fluid
C1988514|Glucose.PO &#x7C; Dose
C0363669|Glucose^4H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363669|Glucose [Mass/volume] in Serum or Plasma --4 hours post 100 g glucose PO
C0363669|Glucose^4 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363669|Glucose 4h p 100 g Glc PO SerPl-mCnc
C0797938|Glucose^3H post 100 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C0797938|Glucose [Moles/volume] in Serum or Plasma --3 hours post 100 g glucose PO
C0797938|Glucose^3 hours post 100 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797938|Glucose 3h p 100 g Glc PO SerPl-sCnc
C0363650|Glucose^2H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0363650|Glucose [Mass/volume] in Serum or Plasma --2 hours post 50 g lactose PO
C0363650|Glucose^2 hours post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363650|Glucose 2h p 50 g Lac PO SerPl-mCnc
C0363656|Glucose 30M p U/kg Ins IV SerPl-mCnc
C0363656|Glucose [Mass/volume] in Serum or Plasma --30 minutes post 0.05-0.15 U insulin/kg IV post 12H CFst
C0363656|Glucose^30M post 0.05-0.15 U insulin/kg IV post 12H CFst:MCnc:Pt:Ser/Plas:Qn
C0363656|Glucose^30 minutes post 0.05-0.15 U insulin/kg Intravenous post 12 hours Calorie fast:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549982|Glucose [Mass/volume] in Serum or Plasma --2 minutes post XXX challenge
C0549982|Glucose 2M p chal SerPl-mCnc
C0549982|Glucose^2M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549982|Glucose^2 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0804102|Glucose 105M p chal SerPl-mCnc
C0804102|Glucose [Mass/volume] in Serum or Plasma --105 minutes post XXX challenge
C0804102|Glucose^105M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0804102|Glucose^105M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1148004|Glucose^3H post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C1148004|Glucose [Moles/volume] in Serum or Plasma --3 hours post 75 g glucose PO
C1148004|Glucose^3 hours post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1148004|Glucose 3h p 75 g Glc PO SerPl-sCnc
C1544013|Glucose^5M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544013|Glucose 5M pre chal SerPl-mCnc
C1544013|Glucose [Mass/volume] in Serum or Plasma --5 minutes pre XXX challenge
C1544013|Glucose^5 minutes pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544043|Glucose [Mass/volume] in Serum or Plasma --16 minutes post XXX challenge
C1544043|Glucose^16M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544043|Glucose 16m p chal SerPl-mCnc
C1544043|Glucose^16M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544045|Glucose 22M p chal SerPl-mCnc
C1544045|Glucose^22M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544045|Glucose [Mass/volume] in Serum or Plasma --22 minutes post XXX challenge
C1544045|Glucose^22M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542933|Glucose^36H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1542933|Glucose [Mass/volume] in Serum or Plasma --36 hours post XXX challenge
C1542933|Glucose^36H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542933|Glucose 36h p chal SerPl-mCnc
C1544197|Glucose [Moles/volume] in Serum or Plasma --31 hour post XXX challenge
C1544197|Glucose^31H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544197|Glucose^31H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544197|Glucose 31h p chal SerPl-sCnc
C1642055|Glucose [Mass/volume] in Urine --2 hours post dose lactose PO
C1642055|Glucose^2H post dose lactose PO:MCnc:Pt:Urine:Qn
C1642055|Glucose^2 hours post dose lactose Oral:Mass Concentration:Point in time:Urine:Quantitative
C1642055|Glucose 2h p Lac PO Ur-mCnc
C2707122|Glucose^2nd specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707122|Glucose [Moles/volume] in Serum or Plasma --2nd specimen post XXX challenge
C2707122|Glucose sp2 p chal SerPl-sCnc
C2707122|Glucose^2nd specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481982|Glucose^20M post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C3481982|Glucose [Moles/volume] in Serum or Plasma --20 minutes post dose lactose PO
C3481982|Glucose^20 minutes post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481982|Glucose 20M p Lac PO SerPl-sCnc
C0549973|Glucose 15M p 50 g Lac PO SerPl-mCnc
C0549973|Glucose [Mass/volume] in Serum or Plasma --15 minutes post 50 g lactose PO
C0549973|Glucose^15M post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0549973|Glucose^15 minutes post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0797940|Glucose^4H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0797940|Glucose [Moles/volume] in Serum or Plasma --4 hours post dose glucose
C0797940|Glucose^4 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797940|Glucose 4h p Glc SerPl-sCnc
C0942693|Glucose [Mass/volume] in Serum or Plasma --2 hours post dose lactose PO
C0942693|Glucose^2H post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0942693|Glucose^2 hours post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942693|Glucose 2h p Lac PO SerPl-mCnc
C0941771|Glucose [Moles/volume] in Serum or Plasma --pre 50 g glucose PO
C0941771|Glucose^pre 50 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C0941771|Glucose pre 50 g Glc PO SerPl-sCnc
C0941771|Glucose^pre 50 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544163|Glucose 12.5h p chal SerPl-sCnc
C1544163|Glucose^12.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544163|Glucose [Moles/volume] in Serum or Plasma --12.5 hours post XXX challenge
C1544163|Glucose^12.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544173|Glucose [Moles/volume] in Serum or Plasma --20 hours post XXX challenge
C1544173|Glucose 20H p chal SerPl-sCnc
C1544173|Glucose^20H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544173|Glucose^20H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1647453|Glucose^30M post dose lactose PO:MCnc:Pt:Urine:Qn
C1647453|Glucose [Mass/volume] in Urine --30 minutes post dose lactose PO
C1647453|Glucose 30M p Lac PO Ur-mCnc
C1647453|Glucose^30 minutes post dose lactose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0549979|Glucose^2.5H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0549979|Glucose [Presence] in Urine by Test strip --2.5 hours post 75 g glucose PO
C0549979|Glucose^2 1/2 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0549979|Glucose 2.5h p 75 g Glc PO Ur Ql Strip
C0549984|Glucose^3.5H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0549984|Glucose [Presence] in Urine by Test strip --3.5 hours post 75 g glucose PO
C0549984|Glucose^3.5 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0549984|Glucose 3.5h p 75 g Glc PO Ur Ql Strip
C0363625|Glucose 30M p 100 g Glc PO Ur-mCnc
C0363625|Glucose [Mass/volume] in Urine --30 minutes post 100 g glucose PO
C0363625|Glucose^30M post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363625|Glucose^30 minutes post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0800038|Glucose sp1 p chal Ur Ql
C0800038|Glucose [Presence] in Urine --1st specimen post XXX challenge
C0800038|Glucose^1st specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800038|Glucose^1st specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0363644|Glucose^1 hour post dose insulin Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363644|Glucose [Mass/volume] in Serum or Plasma --1 hour post dose insulin IV
C0363644|Glucose^1H post dose insulin IV:MCnc:Pt:Ser/Plas:Qn
C0363644|Glucose 1h p Ins IV SerPl-mCnc
C0797928|Glucose^1H post 50 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C0797928|Glucose [Moles/volume] in Serum or Plasma --1 hour post 50 g glucose PO
C0797928|Glucose^1 hour post 50 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797928|Glucose 1h p 50 g Glc PO SerPl-sCnc
C0550004|Glucose [Mass/volume] in Serum or Plasma --9 hours post XXX challenge
C0550004|Glucose^9H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0550004|Glucose^9H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0550004|Glucose 9h p chal SerPl-mCnc
C0801342|Glucose p Glc SerPl-Imp
C0801342|Glucose^post dose glucose:Imp:Pt:Ser/Plas:Nom
C0801342|Glucose^post dose glucose:Impression/interpretation of study:Point in time:Serum/Plasma:Nominal
C0801342|Glucose [Interpretation] in Serum or Plasma--post dose glucose
C0942751|Glucose [Units/volume] in Serum or Plasma --7th specimen post XXX challenge
C0942751|Glucose^7th specimen post XXX challenge:ACnc:Pt:Ser/Plas:Qn
C0942751|Glucose sp7 p chal SerPl-aCnc
C0942751|Glucose^7th specimen post XXX challenge:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C0941758|Glucose [Moles/volume] in Serum or Plasma --1 hour post XXX challenge
C0941758|Glucose^1H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C0941758|Glucose^1 hour post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941758|Glucose 1h p chal SerPl-sCnc
C0941763|Glucose 30M p chal SerPl-sCnc
C0941763|Glucose^30M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C0941763|Glucose [Moles/volume] in Serum or Plasma --30 minutes post XXX challenge
C0941763|Glucose^30 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544015|Glucose 80M p chal SerPl-mCnc
C1544015|Glucose [Mass/volume] in Serum or Plasma --80 minutes post XXX challenge
C1544015|Glucose^80M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544015|Glucose^80M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544028|Glucose 17.5h p chal SerPl-mCnc
C1544028|Glucose [Mass/volume] in Serum or Plasma --17.5 hours post XXX challenge
C1544028|Glucose^17.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544028|Glucose^17.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544038|Glucose^3M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544038|Glucose [Mass/volume] in Serum or Plasma --3 minutes post XXX challenge
C1544038|Glucose 3M p chal SerPl-mCnc
C1544038|Glucose^3 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544050|Glucose^25H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544050|Glucose [Mass/volume] in Serum or Plasma --25 hours post XXX challenge
C1544050|Glucose^25H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544050|Glucose 25h p chal SerPl-mCnc
C1544158|Glucose [Moles/volume] in Serum or Plasma --9.5 hours post XXX challenge
C1544158|Glucose^9.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544158|Glucose^9.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544158|Glucose 9.5h p chal SerPl-sCnc
C1544178|Glucose 1D p chal SerPl-sCnc
C1544178|Glucose [Moles/volume] in Serum or Plasma --1 day post XXX challenge
C1544178|Glucose^1D post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544178|Glucose^1 day post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542951|Glucose [Moles/volume] in Serum or Plasma --19 minutes post XXX challenge
C1542951|Glucose 19M p chal SerPl-sCnc
C1542951|Glucose^19M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542951|Glucose^19M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542954|Glucose^27M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542954|Glucose 27M p chal SerPl-sCnc
C1542954|Glucose [Moles/volume] in Serum or Plasma --27 minutes post XXX challenge
C1542954|Glucose^27M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1714484|Glucose^2H post meal:MCnc:Pt:Milk:Qn
C1714484|Glucose [Mass/volume] in Milk --2 hours post meal
C1714484|Glucose^2 hours post meal:Mass Concentration:Point in time:Milk:Quantitative
C1714484|Glucose 2h p meal Mlk-mCnc
C2360464|Glucose [Mass/volume] in Serum or Plasma --2.5 hours post dose fructose PO
C2360464|Glucose^2.5H post dose fructose PO:MCnc:Pt:Ser/Plas:Qn
C2360464|Glucose^2 1/2 hours post dose fructose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2360464|Glucose 2.5h p fructose PO SerPl-mCnc
C1952722|Glucose 8 PM SerPl-mCnc
C1952722|Glucose [Mass/volume] in Serum or Plasma --8 PM specimen
C1952722|Glucose^8 PM specimen:MCnc:Pt:Ser/Plas:Qn
C1952722|Glucose^8 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954698|Glucose 10 PM SerPl-mCnc
C1954698|Glucose^10 PM specimen:MCnc:Pt:Ser/Plas:Qn
C1954698|Glucose [Mass/volume] in Serum or Plasma --10 PM specimen
C1954698|Glucose^10 PM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954184|Glucose [Mass/volume] in Serum or Plasma --1 hour post dose fructose PO
C1954184|Glucose^1H post dose fructose PO:MCnc:Pt:Ser/Plas:Qn
C1954184|Glucose^1 hour post dose fructose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954184|Glucose 1h p fructose PO SerPl-mCnc
C1954186|Glucose 30M p fructose PO SerPl-mCnc
C1954186|Glucose^30M post dose fructose PO:MCnc:Pt:Ser/Plas:Qn
C1954186|Glucose [Mass/volume] in Serum or Plasma --30 minutes post dose fructose PO
C1954186|Glucose^30 minutes post dose fructose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2598590|Glucose [Moles/volume] in Serum or Plasma --45 minutes post dose betaxolol
C2598590|Glucose 45M p betaxolol SerPl-sCnc
C2598590|Glucose^45M post dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598590|Glucose^45M post dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706905|Glucose^8th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2706905|Glucose sp8 p chal SerPl-sCnc
C2706905|Glucose [Moles/volume] in Serum or Plasma --8th specimen post XXX challenge
C2706905|Glucose^8th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484580|Glucose [Presence] in Urine by Test strip --1 hour post 75 g glucose PO
C0484580|Glucose^1H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484580|Glucose^1 hour post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484580|Glucose 1h p 75 g Glc PO Ur Ql Strip
C0363626|Glucose^1.5H post 0.5 g/kg glucose IV:MCnc:Pt:Ser/Plas:Qn
C0363626|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post 0.5 g/kg glucose IV
C0363626|Glucose^1 1/2 hour post 0.5 g/kg glucose Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363626|Glucose 1.5h p .5 g/kg Glc IV SerPl-mCnc
C0549980|Glucose [Mass/volume] in Serum or Plasma --20 minutes post XXX challenge
C0549980|Glucose 20M p chal SerPl-mCnc
C0549980|Glucose^20M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549980|Glucose^20 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0804103|Glucose^45M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0804103|Glucose 45M p chal SerPl-mCnc
C0804103|Glucose [Mass/volume] in Serum or Plasma --45 minutes post XXX challenge
C0804103|Glucose^45M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942495|Glucose [Mass/volume] in Urine --5 hours post dose glucose
C0942495|Glucose^5H post dose glucose:MCnc:Pt:Urine:Qn
C0942495|Glucose^5 hours post dose glucose:Mass Concentration:Point in time:Urine:Quantitative
C0942495|Glucose 5h p Glc Ur-mCnc
C0942497|Glucose^6H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0942497|Glucose [Mass/volume] in Serum or Plasma --6 hours post dose glucose
C0942497|Glucose^6 hours post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942497|Glucose 6h p Glc SerPl-mCnc
C0941769|Glucose^6H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0941769|Glucose [Moles/volume] in Serum or Plasma --6 hours post dose glucose
C0941769|Glucose^6 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941769|Glucose 6h p Glc SerPl-sCnc
C1542980|Glucose^4H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542980|Glucose [Moles/volume] in Serum or Plasma --4 hours post XXX challenge
C1542980|Glucose^4 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542980|Glucose 4h p chal SerPl-sCnc
C1544180|Glucose^20M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544180|Glucose [Moles/volume] in Serum or Plasma --20 minutes pre XXX challenge
C1544180|Glucose 20M pre chal SerPl-sCnc
C1544180|Glucose^20 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544256|Glucose [Moles/volume] in Serum or Plasma --3 hours post dose lactose PO
C1544256|Glucose^3H post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C1544256|Glucose^3 hours post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544256|Glucose 3h p Lac PO SerPl-sCnc
C1716206|Glucose^4 PM specimen:SCnc:Pt:Ser/Plas:Qn
C1716206|Glucose [Moles/volume] in Serum or Plasma --4 PM specimen
C1716206|Glucose 4 PM SerPl-sCnc
C1716206|Glucose^4 PM specimen:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706824|Glucose^15M pre dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706824|Glucose [Moles/volume] in Serum or Plasma --15 minutes pre dose insulin IV
C2706824|Glucose 15M pre Ins IV SerPl-sCnc
C2706824|Glucose^15 minutes pre dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484590|Glucose 30M p 75 g Glc PO Ur Ql Strip
C0484590|Glucose^30M post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484590|Glucose [Presence] in Urine by Test strip --30 minutes post 75 g glucose PO
C0484590|Glucose^30 minutes post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484594|Glucose [Presence] in Urine by Test strip --4 hours post 75 g glucose PO
C0484594|Glucose^4H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484594|Glucose^4 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484594|Glucose 4h p 75 g Glc PO Ur Ql Strip
C3482270|Glucose^pre 100 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3482270|Glucose^pre 100 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C3482270|Glucose pre 100 g Glc PO SerPl-sCnc
C3482270|Glucose [Moles/volume] in Serum or Plasma --pre 100 g glucose PO
C1988489|Glucose &#x7C; dialysis fluid peritoneal
C0363635|Glucose [Mass/volume] in Serum or Plasma --1 hour post 100 g glucose PO
C0363635|Glucose^1H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363635|Glucose^1 hour post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363635|Glucose 1h p 100 g Glc PO SerPl-mCnc
C0363678|Glucose [Mass/volume] in Serum or Plasma --baseline
C0363678|Glucose^baseline:MCnc:Pt:Ser/Plas:Qn
C0363678|Glucose BS SerPl-mCnc
C0363678|Glucose^baseline:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549967|Glucose [Mass/volume] in Serum or Plasma --10th specimen post XXX challenge
C0549967|Glucose^10th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549967|Glucose sp10 p chal SerPl-mCnc
C0549967|Glucose^10th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549971|Glucose^13th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549971|Glucose [Mass/volume] in Serum or Plasma --13th specimen post XXX challenge
C0549971|Glucose sp13 p chal SerPl-mCnc
C0549971|Glucose^13th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549997|Glucose [Mass/volume] in Serum or Plasma --7.5 hours post XXX challenge
C0549997|Glucose^7.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549997|Glucose^7.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549997|Glucose 7.5h p chal SerPl-mCnc
C0942507|Glucose [Mass/volume] in Serum or Plasma --3.5 hours post dose glucose
C0942507|Glucose^3.5H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0942507|Glucose^3.5 hours post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942507|Glucose 3.5h p Glc SerPl-mCnc
C0941765|Glucose^45M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0941765|Glucose 45M p Glc SerPl-sCnc
C0941765|Glucose [Moles/volume] in Serum or Plasma --45 minutes post dose glucose
C0941765|Glucose^45M post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544021|Glucose^11.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544021|Glucose [Mass/volume] in Serum or Plasma --11.5 hours post XXX challenge
C1544021|Glucose^11.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544021|Glucose 11.5h p chal SerPl-mCnc
C1544261|Glucose [Moles/volume] in Serum or Plasma --75 minutes post dose glucose
C1544261|Glucose 75M p Glc SerPl-sCnc
C1544261|Glucose^75M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C1544261|Glucose^75M post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544299|Glucose [Moles/volume] in Serum or Plasma --3 hours post dose triple bolus
C1544299|Glucose^3H post dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C1544299|Glucose^3 hours post dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544299|Glucose 3h p Triple Bolus SerPl-sCnc
C2360465|Glucose^1.5H post dose fructose PO:MCnc:Pt:Ser/Plas:Qn
C2360465|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post dose fructose PO
C2360465|Glucose^1 1/2 hour post dose fructose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2360465|Glucose 1.5h p fructose PO SerPl-mCnc
C1952856|Glucose [Moles/volume] in Serum or Plasma --pre dose glucose
C1952856|Glucose pre Glc SerPl-sCnc
C1952856|Glucose^pre dose glucose:SCnc:Pt:Ser/Plas:Qn
C1952856|Glucose^pre dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706821|Glucose^2 hours post dose insulin Intravenous:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706821|Glucose^2H post dose insulin IV:SCnc:Pt:Ser/Plas:Qn
C2706821|Glucose [Moles/volume] in Serum or Plasma --2 hours post dose insulin IV
C2706821|Glucose 2h p Ins IV SerPl-sCnc
C1988497|Glucose &#x7C; urine
C0482537|Glucose [Mass/volume] in Serum or Plasma --30 minutes post 75 g glucose PO
C0482537|Glucose 30M p 75 g Glc PO SerPl-mCnc
C0482537|Glucose^30M post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0482537|Glucose^30 minutes post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363637|Glucose^1H post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363637|Glucose [Mass/volume] in Urine --1 hour post 100 g glucose PO
C0363637|Glucose^1 hour post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363637|Glucose 1h p 100 g Glc PO Ur-mCnc
C0363641|Glucose^1H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363641|Glucose [Mass/volume] in Serum or Plasma --1 hour post 75 g glucose PO
C0363641|Glucose^1 hour post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363641|Glucose 1h p 75 g Glc PO SerPl-mCnc
C0363653|Glucose^2H post 75 g glucose PO:MCnc:Pt:Urine:Qn
C0363653|Glucose [Mass/volume] in Urine --2 hours post 75 g glucose PO
C0363653|Glucose^2 hours post 75 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363653|Glucose 2h p 75 g Glc PO Ur-mCnc
C0482535|Glucose^2H post meal:MCnc:Pt:Ser/Plas:Qn
C0482535|Glucose [Mass/volume] in Serum or Plasma --2 hours post meal
C0482535|Glucose^2 hours post meal:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0482535|Glucose 2h p meal SerPl-mCnc
C0796798|Glucose^4H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0796798|Glucose [Mass/volume] in Serum or Plasma --4 hours post 50 g lactose PO
C0796798|Glucose^4 hours post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0796798|Glucose 4h p 50 g Lac PO SerPl-mCnc
C0549986|Glucose [Mass/volume] in Serum or Plasma --3rd specimen post XXX challenge
C0549986|Glucose sp3 p chal SerPl-mCnc
C0549986|Glucose^3rd specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549986|Glucose^3rd specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549972|Glucose^14th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549972|Glucose sp14 p chal SerPl-mCnc
C0549972|Glucose [Mass/volume] in Serum or Plasma --14th specimen post XXX challenge
C0549972|Glucose^14th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0550003|Glucose sp8 p chal DiafP-mCnc
C0550003|Glucose^8th specimen post XXX challenge:MCnc:Pt:Dial fld prt:Qn
C0550003|Glucose [Mass/volume] in Peritoneal dialysis fluid --8th specimen post XXX challenge
C0550003|Glucose^8th specimen post XXX challenge:Mass Concentration:Point in time:Peritoneal dialysis fluid:Quantitative
C0549965|Glucose [Mass/volume] in Serum or Plasma --10 minutes post XXX challenge
C0549965|Glucose 10M p chal SerPl-mCnc
C0549965|Glucose^10M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549965|Glucose^10 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803251|Glucose^2H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0803251|Glucose [Mass/volume] in Serum or Plasma --2 hours post dose glucose
C0803251|Glucose^2 hours post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0803251|Glucose 2h p Glc SerPl-mCnc
C0802043|Glucose^3H post dose glucose:Imp:Pt:Ser/Plas:Nom
C0802043|Glucose^3 hours post dose glucose:Impression/interpretation of study:Point in time:Serum/Plasma:Nominal
C0802043|Glucose 3h p Glc SerPl-Imp
C0802043|Glucose [Interpretation] in Serum or Plasma--3 hours post dose glucose
C0942692|Glucose^1H post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0942692|Glucose [Mass/volume] in Serum or Plasma --1 hour post dose lactose PO
C0942692|Glucose^1 hour post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942692|Glucose 1h p Lac PO SerPl-mCnc
C0945404|Glucose^4H post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0945404|Glucose [Mass/volume] in Serum or Plasma --4 hours post dose lactose PO
C0945404|Glucose^4 hours post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0945404|Glucose 4h p Lac PO SerPl-mCnc
C0942694|Glucose^5H post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0942694|Glucose [Mass/volume] in Serum or Plasma --5 hours post dose lactose PO
C0942694|Glucose^5 hours post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942694|Glucose 5h p Lac PO SerPl-mCnc
C1542930|Glucose^29H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1542930|Glucose [Mass/volume] in Serum or Plasma --29 hours post XXX challenge
C1542930|Glucose^29H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1542930|Glucose 29h p chal SerPl-mCnc
C1544170|Glucose [Moles/volume] in Serum or Plasma --18 hours post XXX challenge
C1544170|Glucose^18H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544170|Glucose 18h p chal SerPl-sCnc
C1544170|Glucose^18H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544238|Glucose [Mass/volume] in Serum or Plasma --3 minutes pre XXX challenge
C1544238|Glucose 3M pre chal SerPl-mCnc
C1544238|Glucose^3M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544238|Glucose^3 minutes pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954898|Glucose^2H post dose glucose:MCnc:Pt:Bld:Qn
C1954898|Glucose [Mass/volume] in Blood --2 hours post dose glucose
C1954898|Glucose^2 hours post dose glucose:Mass Concentration:Point in time:Whole blood:Quantitative
C1954898|Glucose 2h p Glc Bld-mCnc
C2598591|Glucose^1H post dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598591|Glucose [Moles/volume] in Serum or Plasma --1 hour post dose betaxolol
C2598591|Glucose^1 hour post dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598591|Glucose 1h p betaxolol SerPl-sCnc
C0484588|Glucose^3.5H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484588|Glucose [Mass/volume] in Serum or Plasma --3.5 hours post 75 g glucose PO
C0484588|Glucose^3.5 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484588|Glucose 3.5h p 75 g Glc PO SerPl-mCnc
C0484576|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post 50 g lactose PO
C0484576|Glucose^1.5H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0484576|Glucose^1 1/2 hour post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484576|Glucose 1.5h p 50 g Lac PO SerPl-mCnc
C3533248|Glucose.serum-glucose.pericard fld
C1988499|Glucose &#x7C; XXX
C0363658|Glucose [Mass/volume] in Serum or Plasma --30 minutes post 100 g glucose PO
C0363658|Glucose 30M p 100 g Glc PO SerPl-mCnc
C0363658|Glucose^30M post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363658|Glucose^30 minutes post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363661|Glucose^30 minutes post dose insulin Intravenous:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363661|Glucose^30M post dose insulin IV:MCnc:Pt:Ser/Plas:Qn
C0363661|Glucose [Mass/volume] in Serum or Plasma --30 minutes post dose insulin IV
C0363661|Glucose 30M p Ins IV SerPl-mCnc
C0800039|Glucose [Presence] in Urine --2nd specimen post XXX challenge
C0800039|Glucose sp2 p chal Ur Ql
C0800039|Glucose^2nd specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800039|Glucose^2nd specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0800041|Glucose [Presence] in Urine --4th specimen post XXX challenge
C0800041|Glucose^4th specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800041|Glucose sp4 p chal Ur Ql
C0800041|Glucose^4th specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0800044|Glucose^7th specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800044|Glucose sp7 p chal Ur Ql
C0800044|Glucose [Presence] in Urine --7th specimen post XXX challenge
C0800044|Glucose^7th specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0363673|Glucose [Mass/volume] in Urine --5 hours post 100 g glucose PO
C0363673|Glucose^5H post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363673|Glucose^5 hours post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363673|Glucose 5h p 100 g Glc PO Ur-mCnc
C0797930|Glucose^1H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0797930|Glucose [Moles/volume] in Serum or Plasma --1 hour post dose glucose
C0797930|Glucose^1 hour post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797930|Glucose 1h p Glc SerPl-sCnc
C0796797|Glucose^3H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0796797|Glucose [Mass/volume] in Serum or Plasma --3 hours post 50 g lactose PO
C0796797|Glucose^3 hours post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0796797|Glucose 3h p 50 g Lac PO SerPl-mCnc
C0797323|Glucose^5.5H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0797323|Glucose [Mass/volume] in Serum or Plasma --5.5 hours post 75 g glucose PO
C0797323|Glucose^5.5 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0797323|Glucose 5.5h p 75 g Glc PO SerPl-mCnc
C0549983|Glucose [Mass/volume] in Serum or Plasma --2nd specimen post XXX challenge
C0549983|Glucose^2nd specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549983|Glucose sp2 p chal SerPl-mCnc
C0549983|Glucose^2nd specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549964|Glucose^10H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549964|Glucose [Mass/volume] in Serum or Plasma --10 hours post XXX challenge
C0549964|Glucose^10H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549964|Glucose 10h p chal SerPl-mCnc
C0550357|Glucose [Mass/volume] in Serum or Plasma --15 minutes post 100 g glucose PO
C0550357|Glucose^15M post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0550357|Glucose 15M p 100 g Glc PO SerPl-mCnc
C0550357|Glucose^15 minutes post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0880214|Glucose [Moles/volume] in Urine by Test strip
C0880214|Glucose:SCnc:Pt:Urine:Qn:Test strip
C0880214|Glucose Ur Strip-sCnc
C0880214|Glucose:Substance Concentration:Point in time:Urine:Quantitative:Test strip
C0945746|Glucose^6H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0945746|Glucose [Mass/volume] in Serum or Plasma --6 hours post XXX challenge
C0945746|Glucose^6 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0945746|Glucose 6h p chal SerPl-mCnc
C0945403|Glucose^1.5H post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0945403|Glucose [Mass/volume] in Serum or Plasma --1.5 hours post dose lactose PO
C0945403|Glucose^1 1/2 hour post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0945403|Glucose 1.5h p Lac PO SerPl-mCnc
C0941572|Glucose [Presence] in Urine by Test strip
C0941572|Glucose Ur Ql Strip
C0941572|Glucose:ACnc:Pt:Urine:Ord:Test strip
C0941572|Glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C1544149|Glucose 10M p chal SerPl-sCnc
C1544149|Glucose [Moles/volume] in Serum or Plasma --10 minutes post XXX challenge
C1544149|Glucose^10M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544149|Glucose^10 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544150|Glucose [Moles/volume] in Serum or Plasma --15 minutes post XXX challenge
C1544150|Glucose^15M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544150|Glucose 15M p chal SerPl-sCnc
C1544150|Glucose^15 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544196|Glucose^30H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544196|Glucose [Moles/volume] in Serum or Plasma --30 hours post XXX challenge
C1544196|Glucose 30H p chal SerPl-sCnc
C1544196|Glucose^30H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544198|Glucose^36H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544198|Glucose [Moles/volume] in Serum or Plasma --36 hours post XXX challenge
C1544198|Glucose^36H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544198|Glucose 36h p chal SerPl-sCnc
C2361537|Glucose [Mass/volume] in Serum or Plasma --pre-meal
C2361537|Glucose^pre-meal:MCnc:Pt:Ser/Plas:Qn
C2361537|Glucose pre-meal SerPl-mCnc
C2361537|Glucose^pre-meal:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1978482|Glucose [Presence] in Urine by Automated test strip
C1978482|Glucose:ACnc:Pt:Urine:Ord:Test strip.automated
C1978482|Glucose Ur Ql Strip.auto
C1978482|Glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip.automated
C2707125|Glucose sp9 p chal SerPl-sCnc
C2707125|Glucose^9th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707125|Glucose [Moles/volume] in Serum or Plasma --9th specimen post XXX challenge
C2707125|Glucose^9th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481985|Glucose [Moles/volume] in Serum or Plasma --40 minutes post 50 g lactose PO
C3481985|Glucose^40M post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C3481985|Glucose^40M post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3481985|Glucose 40M p 50 g lac PO SerPl-sCnc
C0363672|Glucose [Mass/volume] in Serum or Plasma --5 hours post 100 g glucose PO
C0363672|Glucose^5H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363672|Glucose^5 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363672|Glucose 5h p 100 g Glc PO SerPl-mCnc
C0797925|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post 50 g lactose PO
C0797925|Glucose^1.5H post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C0797925|Glucose^1 1/2 hour post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797925|Glucose 1.5h p 50 g Lac PO SerPl-sCnc
C0549991|Glucose sp4 p chal SerPl-mCnc
C0549991|Glucose [Mass/volume] in Serum or Plasma --4th specimen post XXX challenge
C0549991|Glucose^4th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549991|Glucose^4th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549996|Glucose sp6 p Lac SerPl-mCnc
C0549996|Glucose [Mass/volume] in Serum or Plasma --6th specimen post dose lactose
C0549996|Glucose^6th specimen post dose lactose:MCnc:Pt:Ser/Plas:Qn
C0549996|Glucose^6th specimen post dose lactose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0944798|Glucose^2.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0944798|Glucose [Mass/volume] in Serum or Plasma --2.5 hours post XXX challenge
C0944798|Glucose^2 1/2 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0944798|Glucose 2.5h p chal SerPl-mCnc
C0942502|Glucose^3H post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942502|Glucose [Presence] in Urine by Test strip --3 hours post dose glucose
C0942502|Glucose^3 hours post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0942502|Glucose 3h p Glc Ur Ql Strip
C0945506|Glucose^8th specimen post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0945506|Glucose sp8 p chal SerPl-mCnc
C0945506|Glucose [Mass/volume] in Serum or Plasma --8th specimen post XXX challenge
C0945506|Glucose^8th specimen post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0945252|Glucose^2.5H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0945252|Glucose [Moles/volume] in Serum or Plasma --2.5 hours post dose glucose
C0945252|Glucose^2 1/2 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0945252|Glucose 2.5h p Glc SerPl-sCnc
C1544146|Glucose [Moles/volume] in Serum or Plasma --10 minutes pre XXX challenge
C1544146|Glucose^10M pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544146|Glucose 10M pre chal SerPl-sCnc
C1544146|Glucose^10 minutes pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544155|Glucose 75M p chal SerPl-sCnc
C1544155|Glucose^75M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544155|Glucose [Moles/volume] in Serum or Plasma --75 minutes post XXX challenge
C1544155|Glucose^75M post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542984|Glucose^7H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542984|Glucose [Moles/volume] in Serum or Plasma --7 hours post XXX challenge
C1542984|Glucose^7 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1542984|Glucose 7h p chal SerPl-sCnc
C1542987|Glucose [Moles/volume] in Serum or Plasma --8.5 hours post XXX challenge
C1542987|Glucose^8.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1542987|Glucose 8.5h p chal SerPl-sCnc
C1542987|Glucose^8.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544298|Glucose^2H post dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C1544298|Glucose [Moles/volume] in Serum or Plasma --2 hours post dose triple bolus
C1544298|Glucose^2 hours post dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544298|Glucose 2h p Triple Bolus SerPl-sCnc
C1544191|Glucose [Moles/volume] in Serum or Plasma --25 hours post XXX challenge
C1544191|Glucose^25H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544191|Glucose^25H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544191|Glucose 25h p chal SerPl-sCnc
C1642554|Glucose^6H post dose lactose PO:MCnc:Pt:Urine:Qn
C1642554|Glucose [Mass/volume] in Urine --6 hours post dose lactose PO
C1642554|Glucose^6 hours post dose lactose Oral:Mass Concentration:Point in time:Urine:Quantitative
C1642554|Glucose 6h p Lac PO Ur-mCnc
C2361597|Glucose^post CFst:SCnc:Pt:Urine:Qn
C2361597|Fasting glucose [Moles/volume] in Urine
C2361597|Glucose p fast Ur-sCnc
C2361597|Glucose^post Calorie fast:Substance Concentration:Point in time:Urine:Quantitative
C2735752|Glucose^1M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C2735752|Glucose [Mass/volume] in Serum or Plasma --1 minute post XXX challenge
C2735752|Glucose 1M p chal SerPl-mCnc
C2735752|Glucose^1 minute post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706813|Glucose [Moles/volume] in Serum or Plasma --15 minutes pre dose glucagon
C2706813|Glucose 15M pre Gc SerPl-sCnc
C2706813|Glucose^15M pre dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706813|Glucose^15 minutes pre dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706837|Glucose^30M post dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706837|Glucose [Moles/volume] in Serum or Plasma --30 minutes post dose ornithine alpha-ketoglutarate
C2706837|Glucose 30M p OKG SerPl-sCnc
C2706837|Glucose^30 minutes post dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484584|Glucose^2H post 50 g lactose PO:ACnc:Pt:Urine:Ord:Test strip
C0484584|Glucose [Presence] in Urine by Test strip --2 hours post 50 g lactose PO
C0484584|Glucose^2 hours post 50 g lactose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484584|Glucose 2h p 50 g Lac PO Ur Ql Strip
C2923562|Glucose^7 AM specimen:SCnc:Pt:BldC:Qn:Glucometer
C2923562|Glucose [Moles/volume] in Capillary blood by Glucometer --7 AM specimen
C2923562|Glucose 7 AM BldC Glucomtr-sCnc
C2923562|Glucose^7 AM specimen:Substance Concentration:Point in time:Blood capillary:Quantitative:Glucometer
C3655028|Glucose 2.5h p Lac PO SerPl-sCnc
C3655028|Glucose^2 1/2 hours post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3655028|Glucose^2.5H post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C3655028|Glucose [Moles/volume] in Serum or Plasma --2.5 hours post dose lactose PO
C1988495|Glucose &#x7C; Stool
C0484581|Glucose^1H post meal:MCnc:Pt:Ser/Plas:Qn
C0484581|Glucose [Mass/volume] in Serum or Plasma --1 hour post meal
C0484581|Glucose^1 hour post meal:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484581|Glucose 1h p meal SerPl-mCnc
C0799330|Glucose [Mass/volume] in Serum or Plasma --10 AM specimen
C0799330|Glucose 10 AM SerPl-mCnc
C0799330|Glucose^10 AM specimen:MCnc:Pt:Ser/Plas:Qn
C0799330|Glucose^10 AM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0798169|Glucose^pre 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C0798169|Glucose pre 75 g Glc PO SerPl-sCnc
C0798169|Glucose [Moles/volume] in Serum or Plasma --pre 75 g glucose PO
C0798169|Glucose^pre 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797937|Glucose [Moles/volume] in Serum or Plasma --30 minutes post dose glucose
C0797937|Glucose^30M post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0797937|Glucose 30M p Glc SerPl-sCnc
C0797937|Glucose^30 minutes post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0549974|Glucose^15M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549974|Glucose 15M p chal SerPl-mCnc
C0549974|Glucose [Mass/volume] in Serum or Plasma --15 minutes post XXX challenge
C0549974|Glucose^15 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0550001|Glucose^8H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0550001|Glucose [Mass/volume] in Serum or Plasma --8 hours post XXX challenge
C0550001|Glucose^8 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0550001|Glucose 8h p chal SerPl-mCnc
C0941764|Glucose^4.5H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0941764|Glucose [Moles/volume] in Serum or Plasma --4.5 hours post dose glucose
C0941764|Glucose^4.5 hours post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0941764|Glucose 4.5h p Glc SerPl-sCnc
C1114892|Glucose [Mass/volume] in Serum or Plasma --3 hours post 1.2 g/kg lactose PO
C1114892|Glucose^3H post 1.2 g/kg lactose PO:MCnc:Pt:Ser/Plas:Qn
C1114892|Glucose^3 hours post 1.2 g/kg lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1114892|Glucose 3h p 1.2 g/kg Lac PO SerPl-mCnc
C1544025|Glucose 14h p chal SerPl-mCnc
C1544025|Glucose [Mass/volume] in Serum or Plasma --14 hours post XXX challenge
C1544025|Glucose^14H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544025|Glucose^14H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544039|Glucose [Mass/volume] in Serum or Plasma --6 minutes post XXX challenge
C1544039|Glucose 6M p chal SerPl-mCnc
C1544039|Glucose^6 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544039|Glucose^wapost XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544039|Glucose^ 6M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544252|Glucose^30M post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C1544252|Glucose [Moles/volume] in Serum or Plasma --30 minutes post dose lactose PO
C1544252|Glucose 30M p Lac PO SerPl-sCnc
C1544252|Glucose^30 minutes post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2707123|Glucose [Moles/volume] in Serum or Plasma --3rd specimen post XXX challenge
C2707123|Glucose^3rd specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707123|Glucose sp3 p chal SerPl-sCnc
C2707123|Glucose^3rd specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924058|Glucose^4H post XXX challenge:SCncDiff:Pt:Ser/Plas:Qn
C2924058|Glucose [Molar concentration difference] in Serum or Plasma --4 hours post XXX challenge
C2924058|Glucose^4 hours post XXX challenge:Difference in Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924058|Glucose 4h p chal SerPl-SCDiff
C2703882|Glucose &#x7C; Water
C0797926|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post dose glucose
C0797926|Glucose^1.5H post dose glucose:SCnc:Pt:Ser/Plas:Qn
C0797926|Glucose^1 1/2 hour post dose glucose:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797926|Glucose 1.5h p Glc SerPl-sCnc
C0797935|Glucose^2H post meal:SCnc:Pt:Ser/Plas:Qn
C0797935|Glucose [Moles/volume] in Serum or Plasma --2 hours post meal
C0797935|Glucose^2 hours post meal:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0797935|Glucose 2h p meal SerPl-sCnc
C0797942|Glucose BS SerPl-sCnc
C0797942|Glucose^baseline:SCnc:Pt:Ser/Plas:Qn
C0797942|Glucose [Moles/volume] in Serum or Plasma --baseline
C0797942|Glucose^baseline:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0942752|Glucose^8th specimen post XXX challenge:ACnc:Pt:Ser/Plas:Qn
C0942752|Glucose [Units/volume] in Serum or Plasma --8th specimen post XXX challenge
C0942752|Glucose sp8 p chal SerPl-aCnc
C0942752|Glucose^8th specimen post XXX challenge:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative
C1148006|Glucose^5H post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C1148006|Glucose [Moles/volume] in Serum or Plasma --5 hours post 75 g glucose PO
C1148006|Glucose^5 hours post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1148006|Glucose 5h p 75 g Glc PO SerPl-sCnc
C1544014|Glucose^5M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544014|Glucose 5M p chal SerPl-mCnc
C1544014|Glucose [Mass/volume] in Serum or Plasma --5 minutes post XXX challenge
C1544014|Glucose^5 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544024|Glucose [Mass/volume] in Serum or Plasma --13.5 hours post XXX challenge
C1544024|Glucose 13.5h p chal SerPl-mCnc
C1544024|Glucose^13.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544024|Glucose^13.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544035|Glucose^22H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544035|Glucose [Mass/volume] in Serum or Plasma --22 hours post XXX challenge
C1544035|Glucose^22H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544035|Glucose 22h p chal SerPl-mCnc
C1544165|Glucose [Moles/volume] in Serum or Plasma --13.5 hours post XXX challenge
C1544165|Glucose 13.5h p chal SerPl-sCnc
C1544165|Glucose^13.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544165|Glucose^13.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544254|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post dose lactose PO
C1544254|Glucose^1.5H post dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C1544254|Glucose^1 1/2 hour post dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544254|Glucose 1.5h p Lac PO SerPl-sCnc
C1544263|Glucose^1H post meal:SCnc:Pt:Ser/Plas:Qn
C1544263|Glucose [Moles/volume] in Serum or Plasma --1 hour post meal
C1544263|Glucose^1 hour post meal:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544263|Glucose 1h p meal SerPl-sCnc
C2734078|Glucose^1H post meal:MCnc:Pt:Urine:Qn
C2734078|Glucose [Mass/volume] in Urine --1 hour post meal
C2734078|Glucose^1 hour post meal:Mass Concentration:Point in time:Urine:Quantitative
C2734078|Glucose 1h p meal Ur-mCnc
C2706831|Glucose pre OKG SerPl-sCnc
C2706831|Glucose [Moles/volume] in Serum or Plasma --pre dose ornithine alpha-ketoglutarate
C2706831|Glucose^pre dose ornithine alpha-ketoglutarate:SCnc:Pt:Ser/Plas:Qn
C2706831|Glucose^pre dose ornithine alpha-ketoglutarate:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598587|Glucose^3H post dose betaxolol:SCnc:Pt:Ser/Plas:Qn
C2598587|Glucose [Moles/volume] in Serum or Plasma --3 hours post dose betaxolol
C2598587|Glucose^3 hours post dose betaxolol:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2598587|Glucose 3h p betaxolol SerPl-sCnc
C2707118|Glucose [Moles/volume] in Serum or Plasma --1st specimen post XXX challenge
C2707118|Glucose sp1 p chal SerPl-sCnc
C2707118|Glucose^1st specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707118|Glucose^1st specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2707119|Glucose sp10 p chal SerPl-sCnc
C2707119|Glucose [Moles/volume] in Serum or Plasma --10th specimen post XXX challenge
C2707119|Glucose^10th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2707119|Glucose^10th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2707127|Glucose 10M p Gc SerPl-sCnc
C2707127|Glucose^10M post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2707127|Glucose [Moles/volume] in Serum or Plasma --10 minutes post dose glucagon
C2707127|Glucose^10 minutes post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484593|Glucose^4.5H post 75 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0484593|Glucose [Mass/volume] in Serum or Plasma --4.5 hours post 75 g glucose PO
C0484593|Glucose^4.5 hours post 75 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0484593|Glucose 4.5h p 75 g Glc PO SerPl-mCnc
C0363659|Glucose^30M post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0363659|Glucose 30M p 50 g Lac PO SerPl-mCnc
C0363659|Glucose [Mass/volume] in Serum or Plasma --30 minutes post 50 g lactose PO
C0363659|Glucose^30 minutes post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0800049|Glucose^post meal:MCnc:Pt:Ser/Plas:Qn
C0800049|Glucose p meal SerPl-mCnc
C0800049|Glucose [Mass/volume] in Serum or Plasma --post meal
C0800049|Glucose^post meal:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363647|Glucose^2H post 100 g glucose PO:MCnc:Pt:Ser/Plas:Qn
C0363647|Glucose [Mass/volume] in Serum or Plasma --2 hours post 100 g glucose PO
C0363647|Glucose^2 hours post 100 g glucose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0363647|Glucose 2h p 100 g Glc PO SerPl-mCnc
C0363649|Glucose^2H post 100 g glucose PO:MCnc:Pt:Urine:Qn
C0363649|Glucose [Mass/volume] in Urine --2 hours post 100 g glucose PO
C0363649|Glucose^2 hours post 100 g glucose Oral:Mass Concentration:Point in time:Urine:Quantitative
C0363649|Glucose 2h p 100 g Glc PO Ur-mCnc
C0363688|Glucose^post CFst:MCnc:Pt:BldV:Qn
C0363688|Glucose p fast BldV-mCnc
C0363688|Fasting glucose [Mass/volume] in Venous blood
C0363688|Glucose^post Calorie fast:Mass Concentration:Point in time:Blood venous:Quantitative
C0549966|Glucose 10M pre chal SerPl-mCnc
C0549966|Glucose [Mass/volume] in Serum or Plasma --10 minutes pre XXX challenge
C0549966|Glucose^10M pre XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549966|Glucose^10 minutes pre XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0804104|Glucose^75M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0804104|Glucose 75M p chal SerPl-mCnc
C0804104|Glucose [Mass/volume] in Serum or Plasma --75 minutes post XXX challenge
C0804104|Glucose^75M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942501|Glucose [Presence] in Urine by Test strip --30 minutes post dose glucose
C0942501|Glucose^30M post dose glucose:ACnc:Pt:Urine:Ord:Test strip
C0942501|Glucose 30M p Glc Ur Ql Strip
C0942501|Glucose^30 minutes post dose glucose:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0947225|Glucose [Mass/volume] in Serum or Plasma --3 hours post dose lactose PO
C0947225|Glucose^3H post dose lactose PO:MCnc:Pt:Ser/Plas:Qn
C0947225|Glucose^3 hours post dose lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0947225|Glucose 3h p Lac PO SerPl-mCnc
C1542931|Glucose^30H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1542931|Glucose 30H p chal SerPl-mCnc
C1542931|Glucose [Mass/volume] in Serum or Plasma --30 hours post XXX challenge
C1542931|Glucose^30H post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544151|Glucose^20M post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544151|Glucose [Moles/volume] in Serum or Plasma --20 minutes post XXX challenge
C1544151|Glucose 20M p chal SerPl-sCnc
C1544151|Glucose^20 minutes post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544179|Glucose [Moles/volume] in Serum or Plasma --pre-meal
C1544179|Glucose pre-meal SerPl-sCnc
C1544179|Glucose^pre-meal:SCnc:Pt:Ser/Plas:Qn
C1544179|Glucose^pre-meal:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544239|Glucose^30M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544239|Glucose [Mass/volume] in Serum or Plasma --30 minutes post XXX challenge
C1544239|Glucose 30M p chal SerPl-mCnc
C1544239|Glucose^30 minutes post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1543637|Glucose [Mass/volume] in Serum or Plasma --2nd specimen post dose lactose
C1543637|Glucose^2nd specimen post dose lactose:MCnc:Pt:Ser/Plas:Qn
C1543637|Glucose sp2 p Lac SerPl-mCnc
C1543637|Glucose^2nd specimen post dose lactose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1954701|Glucose 6 AM SerPl-mCnc
C1954701|Glucose [Mass/volume] in Serum or Plasma --6 AM specimen
C1954701|Glucose^6 AM specimen:MCnc:Pt:Ser/Plas:Qn
C1954701|Glucose^6 AM specimen:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2925730|Glucose^pre dose lactose PO:SCnc:Pt:Ser/Plas:Qn
C2925730|Glucose [Moles/volume] in Serum or Plasma --pre dose lactose PO
C2925730|Glucose pre Lac PO SerPl-sCnc
C2925730|Glucose^pre dose lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2707126|Glucose pre Gc SerPl-sCnc
C2707126|Glucose^pre dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2707126|Glucose [Moles/volume] in Serum or Plasma --pre dose glucagon
C2707126|Glucose^pre dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0484598|Glucose^6H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484598|Glucose [Presence] in Urine by Test strip --6 hours post 75 g glucose PO
C0484598|Glucose^6 hours post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484598|Glucose 6h p 75 g Glc PO Ur Ql Strip
C0484578|Glucose^1.5H post 75 g glucose PO:ACnc:Pt:Urine:Ord:Test strip
C0484578|Glucose [Presence] in Urine by Test strip --1.5 hours post 75 g glucose PO
C0484578|Glucose^1 1/2 hour post 75 g glucose Oral:Arbitrary Concentration:Point in time:Urine:Ordinal:Test strip
C0484578|Glucose 1.5h p 75 g Glc PO Ur Ql Strip
C2924053|Glucose [Molar concentration difference] in Serum or Plasma --30 minutes post XXX challenge
C2924053|Glucose^30M post XXX challenge:SCncDiff:Pt:Ser/Plas:Qn
C2924053|Glucose^30 minutes post XXX challenge:Difference in Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924053|Glucose 30M p chal SerPl-SCDiff
C0800040|Glucose^3rd specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800040|Glucose [Presence] in Urine --3rd specimen post XXX challenge
C0800040|Glucose sp3 p chal Ur Ql
C0800040|Glucose^3rd specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0800046|Glucose^9th specimen post XXX challenge:ACnc:Pt:Urine:Ord
C0800046|Glucose sp9 p chal Ur Ql
C0800046|Glucose [Presence] in Urine --9th specimen post XXX challenge
C0800046|Glucose^9th specimen post XXX challenge:Arbitrary Concentration:Point in time:Urine:Ordinal
C0800047|Glucose p fast Ur Ql
C0800047|Glucose^post CFst:ACnc:Pt:Urine:Ord
C0800047|Fasting glucose [Presence] in Urine
C0800047|Glucose^post Calorie fast:Arbitrary Concentration:Point in time:Urine:Ordinal
C0798168|Glucose [Moles/volume] in Serum or Plasma --2 hours post 75 g glucose PO
C0798168|Glucose^2H post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C0798168|Glucose^2 hours post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C0798168|Glucose 2h p 75 g Glc PO SerPl-sCnc
C0797054|Glucose^2.5H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0797054|Glucose [Mass/volume] in Serum or Plasma --2.5 hours post 50 g lactose PO
C0797054|Glucose^2 1/2 hours post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0797054|Glucose 2.5h p 50 g Lac PO SerPl-mCnc
C0797055|Glucose [Mass/volume] in Serum or Plasma --5 hours post 50 g lactose PO
C0797055|Glucose^5H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0797055|Glucose^5 hours post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0797055|Glucose 5h p 50 g Lac PO SerPl-mCnc
C0549994|Glucose [Mass/volume] in Serum or Plasma --6.5 hours post XXX challenge
C0549994|Glucose^6.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549994|Glucose^6.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0549994|Glucose 6.5h p chal SerPl-mCnc
C0549988|Glucose [Mass/volume] in Serum or Plasma --40 minutes post XXX challenge
C0549988|Glucose^40M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C0549988|Glucose 40M p chal SerPl-mCnc
C0549988|Glucose^40M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0801396|Glucose [Mass/volume] in Serum or Plasma --12 hours post 50 g lactose PO
C0801396|Glucose^12H post 50 g lactose PO:MCnc:Pt:Ser/Plas:Qn
C0801396|Glucose^12 hours post 50 g lactose Oral:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0801396|Glucose 12h p 50 g Lac PO SerPl-mCnc
C0942496|Glucose^5H post dose glucose:MCnc:Pt:Ser/Plas:Qn
C0942496|Glucose [Mass/volume] in Serum or Plasma --5 hours post dose glucose
C0942496|Glucose^5 hours post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C0942496|Glucose 5h p Glc SerPl-mCnc
C1544036|Glucose^23.5H post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544036|Glucose [Mass/volume] in Serum or Plasma --23.5 hours post XXX challenge
C1544036|Glucose^23.5 hours post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544036|Glucose 23.5h p chal SerPl-mCnc
C1544042|Glucose [Mass/volume] in Serum or Plasma --14 minutes post XXX challenge
C1544042|Glucose^14M post XXX challenge:MCnc:Pt:Ser/Plas:Qn
C1544042|Glucose 14m p chal SerPl-mCnc
C1544042|Glucose^14M post XXX challenge:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C1544143|Glucose [Moles/volume] in Serum or Plasma --pre XXX challenge
C1544143|Glucose pre chal SerPl-sCnc
C1544143|Glucose^pre XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544143|Glucose^pre XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544156|Glucose [Moles/volume] in Serum or Plasma --2.5 hours post XXX challenge
C1544156|Glucose^2.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544156|Glucose^2 1/2 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544156|Glucose 2.5h p chal SerPl-sCnc
C1544296|Glucose^45M post dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C1544296|Glucose 45M p Triple Bolus SerPl-sCnc
C1544296|Glucose [Moles/volume] in Serum or Plasma --45 minutes post dose triple bolus
C1544296|Glucose^45M post dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544189|Glucose [Moles/volume] in Serum or Plasma --4.5 hours post XXX challenge
C1544189|Glucose^4.5H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C1544189|Glucose^4.5 hours post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C1544189|Glucose 4.5h p chal SerPl-sCnc
C2360270|Glucose^1H post 75 g glucose PO:SCnc:Pt:Ser/Plas:Qn
C2360270|Glucose [Moles/volume] in Serum or Plasma --1 hour post 75 g glucose PO
C2360270|Glucose^1 hour post 75 g glucose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2360270|Glucose 1h p 75 g Glc PO SerPl-sCnc
C1952716|Glucose [Mass/volume] in Serum or Plasma --20 minutes post dose glucose
C1952716|Glucose 20M p Glc SerPl-mCnc
C1952716|Glucose^20M post dose glucose:MCnc:Pt:Ser/Plas:Qn
C1952716|Glucose^20 minutes post dose glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C2706815|Glucose [Moles/volume] in Serum or Plasma --2 minutes post dose glucagon
C2706815|Glucose 2M p Gc SerPl-sCnc
C2706815|Glucose^2M post dose glucagon:SCnc:Pt:Ser/Plas:Qn
C2706815|Glucose^2 minutes post dose glucagon:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2706902|Glucose sp5 p chal SerPl-sCnc
C2706902|Glucose [Moles/volume] in Serum or Plasma --5th specimen post XXX challenge
C2706902|Glucose^5th specimen post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C2706902|Glucose^5th specimen post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924059|Glucose [Molar concentration difference] in Serum or Plasma --5 hours post XXX challenge
C2924059|Glucose^5H post XXX challenge:SCncDiff:Pt:Ser/Plas:Qn
C2924059|Glucose^5 hours post XXX challenge:Difference in Substance Concentration:Point in time:Serum/Plasma:Quantitative
C2924059|Glucose 5h p chal SerPl-SCDiff
C2602566|Estimated average glucose &#x7C; Bld-Ser-Plas
C1506098|IPX 750
C1506098|IPX-750
C1506098|IPX750
C3711206|ethanone-1-C-beta-D-glucopyranoside
C3711206|3,7-anhydro-1-deoxyglycero-gulo-2-octulose
C0533572|1,2-5,6-di-O-isopropylidene-alpha-D-glucofuranosyl (-)-(S)-propanesulfinate
C0533572|1,2-5,6-di-O-isopropylideneglucofuranosyl propanesulfinate
C0533572|DIPrGluco propanesulfinate
C1615567|gem-difluorocarba-D-glucose
C2354010|2,3,4,6-tetra-O-acetylglucopyranosyl bromide
C0630418|3,5-O-benzylidene-1,2-O-isopropylidene-alpha-D-glucofuranose
C0630418|3,5-O-benzylidene-1,2-O-isopropylideneglucofuranose
C0630418|3,5-BIGD
C0049237|5-hydroxymethyl-1,2,3,4-cyclohexanetetrol
C0049237|pseudo-DL-glucose
C0049237|5a-carba-aldohexopyranose
C0049237|5a-carba-glucopyranose
C3660097|1,5-anhydro-2-deoxy-D-ribo-hex-1-enitol
C1098606|4,6-O-B-D-G
C1098606|4,6-O-benzylidene-D-glucopyranose
C0756246|D-glucose,O-beta-D-glucopyranosyl
C0756246|D-glucose, O-D-glucopyranosyl
C0061427|alpha-D-glucopyranosyl fluoride
C0061427|glucosyl fluoride
C1699869|2-epsilon-lysino-2-deoxy-6-phosphoglucose
C1699869|glucoselysine-6-phosphate
C0043756|1,2,3,6-tetragalloylglucose
C0043756|1,2,3,6-TGG
C2974622|4-deoxy-4-fluoro-beta-D-glucopyranose
C0537801|Y-ART 3
C0537801|Y-ART-3
C0620373|4,6-pyruvylated D-glucose
C0620373|4,6-pyruvylated glucose
C0620373|4,6-PYDGLC
C0538894|SQ-1-O-DHA
C0538894|sulfoquinovosyl-1-O-dihydroxyacetone
C0163570|monoacetone-glucose
C0163570|1,2-O-isopropylidene-D-glucofuranose
C1122647|N-benzoyl-N'-glucopyranosylurea
C2745802|TAMAGF cpd
C2745802|3,5,6-triacetyl-1,2-O-isopropylidene-alpha-D-glucofuranose
C1569487|1-O-galloyl-6-O-luteoyl-alpha-D-glucose
C1569487|GLAG cpd
C0759542|UDP-4-keto-6-deoxyglucose
C0249652|3-O-(2-iodoethyl)-D-glucose
C0249652|3-O-(2-iodoethyl)glucose
C0140293|retinoyl beta-glucose
C0140293|retinoylglucose
C0608761|zinc thioglucose
C0630420|1,2,3,4-tetraacetoxy-5-(acetoxymethyl)cyclohexane
C0630420|1,2,3,4-TAMC
C1741296|hexos-4-ulose
C1741296|4-ketoglucose
C0763300|glucose valproate
C0045319|2,3,4,5,6-pentagalloylglucose
C0045319|3-O-digalloyl-1,2,6-trigalloylglucose
C0045319|D-Glucose, 2,3,4,5,6-pentakis(3,4,5-trihydroxybenzoate)
C0649280|pseudo-laminarabiose
C1098234|1-O-methyl-2,3-di-O-galloylglucose
C0617236|alpha-D-Glucofuranose, cyclic 1,2:3,5-bis(butylboronate) 6-acetate
C0617236|D-glucofuranose cyclic 1,2-3,5 bis(butylboronate)-6-acetate
C0617236|glucose BBA
C0061402|D-Glucose, 6-ester with arsenic acid (H3AsO4)
C0061402|glucose 6-arsenate
C1099047|5-fluoroglucopyranosyl fluoride
C1099047|5FGlcF cpd
C0059829|ethylidene glucose
C0059829|4,6-O-ethylidene glucose
C0646794|2,4,6-tri-O-galloyl-D-glucose
C0646794|2,4,6-tri-O-galloylglucose
C0646794|2,4,6-TGDG
C0643789|M-2,3,4-AAGlu
C0643789|methyl 2,3,4-tri-O-acetyl-alpha-D-glucopyranoside
C0643789|methyl 2,3,4-tri-O-acetylglucopyranoside
C1311599|1,3,6-tri-O-galloylglucose
C2717224|1,2,6-tri-O-galloyl-beta-D-allose
C0043771|1,2-5,6-di-O-isopropylidene-D-glucofuranose
C0043771|diacetone glucose
C0658269|3,6-anhydro-D-glucose
C0658269|3,6-anhydroglucose
C1259059|2-D-HBA-G
C1259059|2-deoxy-2-(3-hydroxybutyramido)-glucose
C1620154|1,6-di-O-galloyl-beta-D-glucose
C1122646|N-acetyl-N'-glucopyranosylurea
C0380377|beta-D-Glc-IPM
C0380377|beta-D-glucosylisophosphoramide mustard
C0380377|beta-D-glucosyl-ifosfamide mustard
C1098236|1,2,3-TGG
C1098236|1,2,3-tri-O-galloylglucose
C0533218|3,6-dideoxy-3-((R)-3-hydroxybutyramido)-D-glucose
C0533218|3,6-dideoxy-3-(3-hydroxybutyramido)glucose
C0533218|Qui3NAcyl
C0660802|2-O-carboxymethylglucose
C0244541|3-deoxy-3-iodo-D-glucose
C0053308|4,6-benzylidene-D-glucose
C0053308|alpha-D-Glucopyranose, 4,6-O-(phenylmethylene)-
C0053308|benzylidene glucopyranose
C0053308|benzylidene glucose
C0537306|glucose pentaacetate
C0537306|penta-O-acetyl-alpha-D-glucopyranose
C0537306|penta-O-acetylglucopyranose
C0044632|1-thioglucose
C0049366|5-thio-D-glucose
C3712805|1-O-galloyl-6-O-vanilloyl-beta-glucose
C0251796|D-glucose-L-cysteine
C0251796|glucose-Cys
C0251796|glucose-cysteine
C0044042|1,6-anhydro-beta-D-glucopyranose
C0044042|1,6-anhydro-beta-glucopyranose
C0044042|levoglucosan
C0061437|glucosyl urea
C0061437|glucosylurea
C0061437|glucoseureide
C0061437|glucose-ureide
C0648562|1-fluoroglucopyranosyl fluoride
C0632958|beta-D-Glucopyranose, 1,2,6-tris(3-nitropropanoate)
C0632958|karakin
C0632958|karakine
C3501161|AS-3 solution
C3501161|AS3 solution
C2198636|5% dextrose infusion
C2198636|5% dextrose infusion (medication)
C3847687|Glucose challenge &#x7C; Exhaled gas
C3851301|3,6-O-(o-xylylene)glucopyranosyl fluoride
C3870240|Glucose 45M p 50 g Lac PO SerPl-sCnc
C3870240|Glucose^45M post 50 g lactose Oral:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3870240|Glucose [Moles/volume] in Serum or Plasma --45 minutes post 50 g lactose PO
C3870240|Glucose^45M post 50 g lactose PO:SCnc:Pt:Ser/Plas:Qn
C3870547|Glucose^1 1/2 hour post dose triple bolus:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C3870547|Glucose [Moles/volume] in Serum or Plasma --1.5 hours post dose triple bolus
C3870547|Glucose^1.5H post dose triple bolus:SCnc:Pt:Ser/Plas:Qn
C3870547|Glucose 1.5h p Triple Bolus SerPl-sCnc
C3853667|glucose 24 g/31 g oral gel
C3853667|Glucose 24g Oral gel
C3853667|DEXTROSE 24GM/31GM SQUEEZE TUBE [VA Product]
C3853667|DEXTROSE 24GM/31GM SQUEEZE TUBE
C3853667|dextrose 77.4 % Oral Gel
C3853667|Glucose 0.774 MG/MG Oral Gel
C0011795|Dextran 70
C0011795|plasma expanders dextran hm
C0011795|dextran-70
C0011795|dextran HM
C0011795|plasma expanders dextran-70
C0011795|dextran HM (medication)
C0011795|dextran-70 (medication)
C0011795|Dextran-HM
C0011795|Dextran 70 [Chemical/Ingredient]
C0011795|Dextran M 70
C0011795|Dextran 70 (product)
C0011795|Dextran 70 (substance)
C4036718|Glucose^2H post meal:SCnc:Pt:Ser/Plas/Bld:Qn
C4036718|Glucose^2 hours post meal:Substance Concentration:Point in time:Serum/Plasma/Whole blood:Quantitative
C4036718|Glucose [Moles/volume] in Serum, Plasma or Blood --2 hours post meal
C4036718|Glucose 2h p meal SerPlBld-sCnc
C4036714|Glucose^11H post XXX challenge:SCnc:Pt:Ser/Plas:Qn
C4036714|Glucose 11h p chal SerPl-sCnc
C4036714|Glucose [Moles/volume] in Serum or Plasma --11 hour post XXX challenge
C4036714|Glucose^11H post XXX challenge:Substance Concentration:Point in time:Serum/Plasma:Quantitative
C4040089|Protein-bound glucose (substance)
C4040089|Protein-bound glucose
C4042478|(99m)Tc-2-((3-carboxy-1-oxopropyl)amino)-2-deoxy-D-glucose
C4042478|(99m)Tc-CPADG
C4044340|Somah
C2684476|Glucose 254 MG/ML Oral Solution
C2684476|Glucose Oral Liquid 15 GM/59ML
C2684476|glucose 25% oral liquid
C2684476|Dextrose 25% Oral Solution
C2684476|Glucose 15g Oral solution
C2684476|dextrose 25 % Oral Solution
C2684476|glucose 15 GM / 59 ML Oral Solution
C2684476|glucose 15 GM / 60 ML Oral Solution
C2684476|Glucose 15g/59mL Oral solution
C2684476|DEXTROSE 15GM/59ML ORAL LIQUID
C2684476|DEXTROSE 15GM/59ML LIQUID,ORAL
C2684476|DEXTROSE 15GM/59ML LIQUID,ORAL [VA Product]
C2684476|CVS Glucose 15g Liquid Shot (Grape)
C4070392|Glucose^45M post dose arginine+insulin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C4070392|Glucose [Mass/volume] in Serum or Plasma --45 minutes post dose arginine+insulin
C4070392|Glucose^45M post dose arginine+insulin:MCnc:Pt:Ser/Plas:Qn
C4070392|Glucose 45M p Arg+Ins SerPl-mCnc
C4070394|Glucose [Mass/volume] in Serum or Plasma --15 minutes post dose arginine+insulin
C4070394|Glucose^15 minutes post dose arginine+insulin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C4070394|Glucose 15M p Arg+Ins SerPl-mCnc
C4070394|Glucose^15M post dose arginine+insulin:MCnc:Pt:Ser/Plas:Qn
C4070393|Glucose^30 minutes post dose arginine+insulin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C4070393|Glucose [Mass/volume] in Serum or Plasma --30 minutes post dose arginine+insulin
C4070393|Glucose 30M p Arg+Ins SerPl-mCnc
C4070393|Glucose^30M post dose arginine+insulin:MCnc:Pt:Ser/Plas:Qn
C4070391|Glucose^1 hour post dose arginine+insulin:Mass Concentration:Point in time:Serum/Plasma:Quantitative
C4070391|Glucose^1H post dose arginine+insulin:MCnc:Pt:Ser/Plas:Qn
C4070391|Glucose [Mass/volume] in Serum or Plasma --1 hour post dose arginine+insulin
C4070391|Glucose 1h p Arg+Ins SerPl-mCnc
C4050442|Glucose [Moles/volume] in Peritoneal dialysis fluid --overnight dwell
C4050442|Glucose^overnight dwell:SCnc:Pt:Dial fld prt:Qn
C4050442|Glucose DiafP-sCnc
C4050442|Glucose^overnight dwell:Substance Concentration:Point in time:Peritoneal dialysis fluid:Quantitative
C0538727|icodextrin
C0538727|icodextrin [Chemical/Ingredient]
C0538727|Icodextran
C0538727|Icodextrin (product)
C0538727|Icodextran (product)
C0538727|Icodextrin (substance)
C0063739|invert sugar
C0063739|invertose
C0063739|foods invert sugar (discontinued)
C0063739|invert sugar (discontinued)
C0063739|invert sugar (discontinued) (medication)
C0063739|invert sugar [Chemical/Ingredient]
C0063739|MAIZE INVERT SUGAR
C0063739|Sugar, Invert
C0063739|Corn Invert Sugar
C0063739|Maize Inver Sugar
C1298380|Dextrose 25% solution (product)
C1298380|Dextrose 25% solution
C1302925|10 ML Glucose 50 MG/ML Prefilled Syringe
C1302925|10 ML dextrose 5 % Prefilled Syringe
C1302925|Dextrose 5g/100mL (5%) injection solution 10mL syringe (product)
C1302925|Dextrose 5g/100mL (5%) injection solution 10mL syringe
C0357164|Parenteral glucose
C0357164|Intravenous glucose
C0357164|Parenteral form glucose (product)
C0357164|Parenteral form glucose
C0357164|Parenteral glucose (product)
C0357164|Parenteral glucose (substance)
C0719832|Dextrose 2.5%
C1443653|Dextrose 10% solution (product)
C1443653|Dextrose 10% solution
C1443654|Dextrose 20% solution (product)
C1443654|Dextrose 20% solution
C1443655|Dextrose 30% solution (product)
C1443655|Dextrose 30% solution
C1443656|Dextrose 40% solution (product)
C1443656|Dextrose 40% solution
C0308817|Glucose 500 MG/ML Oral Solution
C0308817|DEXTROSE 50% SOLUTION (product)
C0308817|DEXTROSE 50% SOLUTION
C0308817|DEXTROSE MONOHYDRATE 50 g in 100 mL ORAL LIQUID [Dextrose 50%]
C0308817|Glutol 100g/180ml Solution
C0308817|DEXTROSE 50% SOLUTION (substance)
C0308817|Dextrose 50% Oral Solution
C1443657|Dextrose 60% solution (product)
C1443657|Dextrose 60% solution
C1443658|Dextrose 70% solution (product)
C1443658|Dextrose 70% solution
C1445749|Lactated Ringer solution + dextrose
C1445749|Lactated Ringer's solution + dextrose (product)
C1445749|Lactated Ringer's solution + dextrose
C0887283|Glucose, (alpha-D)-Isomer
C0887284|Glucose, (beta-D)-Isomer
C0887285|Glucose, (DL)-Isomer
C0017734|Monohydrate, Glucose
C0017734|Glucose Monohydrate
C0359954|Dextrose-Lidocaine Hydrochloride
C0359954|Lidocaine Hydrochloride with Dextrose
C0359954|Lignocaine hydrochloride+glucose
C0359954|Lidocaine hydrochloride+glucose (product)
C0359954|Lidocaine hydrochloride+glucose
C0359954|Lignocaine hydrochloride+glucose (product)
C0359954|Lignocaine hydrochloride+glucose (substance)
C0360655|Potassium+dextrose infusion
C0360655|Potassium+dextrose infusion (product)
C0360655|Potassium+dextrose infusion (substance)
C0718770|B-D Glucose
C1613037|CPDA-1 Anticoagulant
C1657066|Delflex A Low Ca Low Mg with 2.5% Dextrose
C1650394|Dextran in Dextrose
C1654896|Steriflex No.6
C0051220|allose
C0601729|popiodol suspension
C0055816|citrate phosphate dextrose
C0055816|citroglucophosphate
C0055816|D-Glucose, mixt. with 2-hydroxy-1,2,3-propanetricarboxylic acid and phosphoric acid
C0055816|ANTICOAGULANT CITRATE DEXTROSE PHOSPHATE
C0055816|citrate phosphate dextrose (medication)
C0055816|CPD
C0603338|hithiol
C0604308|polyketoacidomycin
C0082716|glucose 6-(hydrogen sulfate)
C0082716|glucose sulfate
C0049418|6,6-dideuteroglucose
C0061420|GIK solution
C0061420|GIKCS
C0061420|glucose-insulin-potassium cardioplegic solution
C0061420|glucose-insulin-potassium substrate
C0207603|S-MA(2)
C0207603|S-MA2 solution
C0056450|CPDA solutions
C0163839|Darrow's solution
C0163839|Darrows solution
C0050888|ADSOL
C0050888|AS-1 preservative solution
C0054039|Bretschneider cardioplegic solution
C0054039|HTK solution
C0054039|Custodiol solution
C0054039|histidine-tryptophan-ketoglutarate solution
C0054039|HTK solution of Bretschneider
C0054039|Bretschneider solution
C0058329|Dioralyte
C0078516|rehydration solution, oral, WHO
C0078516|WHO-ORS
C0078516|World Health Organization oral rehydration solution
C0360675|dextrolyte
C0360675|Dextrolyte (product)
C0360675|Dextrolyte (substance)
C0075156|Stanford cardioplegic solution
C0075156|Stanford solution
C0526083|Hicaliq
C0069944|PAGGS-sorbit
C0069944|PAGGS-sorbitol solution
C0635934|PIGPA solution
C0052462|AS-3 preservative solution
C0073555|Roe cardioplegic solution
C0640586|regidrone
C0640586|Rehydron
C0640586|Rehydrone
C0646235|Sweetrex
C0646657|Glc-Spheron
C0167250|Krebs-Henseleit solution
C0167250|KHB solution
C0167250|Krebs-Henseleit buffer
C0174598|TES-Tris buffer
C0174598|TEST yolk buffer
C0174598|TES-Tris yolk buffer
C0220292|LPDG solution
C0220292|low potassium dextran glucose solution
C0254356|Ep4 solution
C0257665|glucose-glycine-formate
C0257665|glucose-glycine-formiate
C0257665|medikhronal
C0257665|medichronal
C0292649|CP 11EB
C0292649|CP-11EB
C0299071|dextrose albumin solution
C0391004|isosal
C0391253|MBS solution
C0531138|STHGAL solution
C0676371|PentaLyte
C0759569|2-deoxy-D-glucose tetraacetate
C0759569|2-deoxy-glucose tetraacetate
C0759569|2-DOG TA
C0759880|fattiviracin A1
C0759880|fattiviracin-A1
C0760344|4'-dehydroxyphlorizin
C0967642|PAGGS-M solution
C1657532|Dex4
C1657532|Dex4 Mango Twist
C1657532|Dex4 Grape
C1657532|Dex4 Assorted Fruit
C1657532|Dex4 Fruit Punch
C1657532|Dex4 Orange
C1657532|Dex4 Raspberry
C1657532|Dex4 Berry Twist
C1657532|Dex4 Citrus Punch
C1657532|Dex4 Natural Orange
C1827843|Glucose + treacle
C1827843|Glucose + treacle (product)
C1827175|caffeine + dextrose (medication)
C1827175|caffeine + dextrose
C1827175|Caffeine / Glucose
C1827175|Caffeine+glucose (product)
C1827175|Caffeine+glucose
C1827175|Caffeine + glucose (product)
C1827175|Caffeine + glucose
C1337358|iso-osmotic dextrose
C2344965|Dianeal PD-2/4.25
C2344988|Aminosyn II 3.5% in 5% Dextrose
C2344992|Dianeal PD-2/2.5
C2345003|Dianeal PD-2/1.5
C2345010|Dianeal Low Calcium 1.5
C2345012|Dianeal Low Calcium 4.25
C2345039|Aminosyn II 4.25% in 10% Dextrose
C2345043|Aminosyn II 4.25% in 20% Dextrose
C2345047|Dianeal Low Calcium 2.5
C2345053|Aminosyn II 4.25/25
C2345281|Clinimix E 4.25/5
C2345299|Clinimix 2.75/5
C2345303|Clinimix 4.25/10
C2345307|Clinimix 4.25/20
C2345311|Clinimix 4.25/25
C2345315|Clinimix 4.25/5
C2345332|Clinimix 5/15
C2345337|Clinimix 5/20
C2345341|Clinimix 5/25
C2345347|Clinimix E 2.75/5
C2345353|Clinimix E 2.75/10
C2345358|Clinimix E 4.25/25
C2345366|Clinimix E 5/15
C2345376|Clinimix E 5/20
C2345378|Clinimix E 5/25
C2345402|Clinimix E 5/35
C2345480|Ionosol-B
C2345490|Ionosol-MB
C2345499|Ionosol-T
C2345519|Isolyte H
C2345602|Isolyte M
C2345614|Isolyte P
C2345761|Normosol-M
C2346032|Travasol 2.75
C2346078|Travasol 2.75/5
C2346120|Travasol 4.25/10
C2346124|Travasol 4.25/25
C2346128|Travasol 4.25/5
C2346361|Dianeal PD-2/3.5
C0364479|Glucose:MCnc:Pt:Bld:Qn
C0364479|Glucose [Mass/volume] in Blood
C0364479|Glucose Bld-mCnc
C0364479|Glucose:Mass Concentration:Point in time:Whole blood:Quantitative
C0523660|Glucose measurement, post glucose dose
C0523660|Glucose measurement, post glucose dose (procedure)
C0337438|Glucose
C0337438|Glucose measurement
C0337438|Test;glucose
C0337438|Measurement of glucose
C0337438|GLUC
C0337438|Glucose measurement (procedure)
C0337438|Glucose measurement, NOS
C0337438|glucose test
C0392201|Blood glucose
C0392201|blood glucose tests (lab test)
C0392201|blood glucose tests
C0392201|Blood glucose measurement
C0392201|blood glucose level
C0392201|blood glucose measurement (lab test)
C0392201|Blood glucose (sugar) level
C0392201|Measurement of glucose in blood
C0392201|Blood Sugar
C0392201|Glucose Measurement, Blood
C0392201|Blood sugar level
C0392201|BS - Blood glucose level
C0392201|Glucose measurement, blood (procedure)
C0202048|Glucose measurement by monitoring device
C0202048|Glucose measurement by monitoring device (procedure)
C0202048|Glucose measurement by monitoring device (procedure) [Ambiguous]
C2732668|Urea, electrolytes and glucose measurement
C2732668|Measurement of urea, sodium, potassium, chloride, bicarbonate and glucose (procedure)
C2732668|Measurement of urea, sodium, potassium, chloride, bicarbonate and glucose
C2732640|Calculation of estimated average glucose based on hemoglobin A1c (procedure)
C2732640|Calculation of estimated average glucose based on hemoglobin A1c
C2732640|Estimated average glucose measurement
C2732640|Calculation of estimated average glucose based on haemoglobin A1c
C0204885|Ward glucometer test
C0204885|Ward glucometer test (procedure)
C0202040|cerebrospinal fluid glucose (lab test)
C0202040|cerebrospinal fluid glucose
C0202040|CSF glucose
C0202040|Glucose CSF
C0202040|Glucose measurement, cerebrospinal fluid
C0202040|Glucose measurement, cerebrospinal fluid (procedure)
C0202040|Glucose measurement, CSF (procedure)
C0202040|CSF Glucose Test
C0202040|Glucose measurement, CSF
C1271625|Urine clinitest
C1271625|Urine clinitest (procedure)
C0202041|serum glucose
C0202041|Serum Glucose Measurement
C0202041|Serum Glucose Test
C0202041|Glucose measurement, serum
C0202041|Glucose measurement, serum (procedure)
C0202042|Plasma Glucose Measurement
C0202042|plasma glucose measurement (lab test)
C0202042|plasma glucose
C0202042|Plasma glucose level
C0202042|Plasma glucose level (procedure)
C0202042|Glucose measurement, plasma
C0202042|Glucose measurement, plasma (procedure)
C0523655|Glucose cerebrospinal fluid/glucose plasma ratio measurement (procedure)
C0523655|Glucose cerebrospinal fluid/glucose plasma ratio measurement
C0523655|Glucose CSF/glucose plasma ratio measurement (procedure)
C0523655|Glucose CSF/glucose plasma ratio measurement
C0004076|urine glucose
C0004076|Glucose measurement, urine
C0004076|urine glucose measurement (lab test)
C0004076|urine glucose measurement
C0004076|Glucose urine
C0004076|Urine screen for sugar (& [glucose]) (procedure)
C0004076|Sugar - urine test (& glucose)
C0004076|Urine glucose test NOS
C0004076|Urine glucose test NOS (procedure)
C0004076|Sugar - urine test (& glucose) (procedure)
C0004076|Urine test for glucose (procedure)
C0004076|Urine screen for sugar (& [glucose])
C0004076|Urine test for glucose
C0004076|Glucose - urine test
C0004076|Sugar - urine test
C0004076|Urine Glucose Test
C0004076|Glucose measurement, urine (procedure)
C0373621|Glucose test; post glucose dose (includes glucose)
C0373621|Glucose; post glucose dose (includes glucose)
C0373621|GLUCOSE POST GLUCOSE DOSE
C0373621|Blood glucose (sugar) level after receiving dose of glucose
C0373621|Measurement of glucose after glucose dose
C0373621|GLUCOSE TEST
C0523658|ASSAY GLUCOSE BLOOD QUANT
C0523658|Glucose; quantitative, blood (except reagent strip)
C0523658|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP
C0523658|Glucose measurement, quantitative
C0523658|Glucose measurement, quantitative (procedure)
C0373622|Glucose; tolerance test (GTT), 3 specimens (includes glucose)
C0373622|GLUCOSE TOLERANCE TEST GTT 3 SPECIMENS
C0373622|Glucose tolerance test (gtt)
C0373623|GLUCOSE TOLERANCE EA ADDL BEYOND 3 SPECIMENS
C0373623|Glucose; tolerance test, each additional beyond 3 specimens (List separately in addition to code for primary procedure)
C0373623|Gtt-added samples
C0373620|Glucose; blood, reagent strip
C0373620|blood glucose determination by reagent strip (lab test)
C0373620|blood glucose determination by reagent strip
C0373620|blood glucose level by reagent strip
C0373620|GLUCOSE BLOOD REAGENT STRIP
C0373620|Blood glucose (sugar) measurement using reagent strip
C0373620|Measurement of glucose in blood using reagent strip
C0373620|REAGENT STRIP/BLOOD GLUCOSE
C4064987|glucose in serum or plasma (lab test)
C4064987|glucose in serum or plasma
C0202045|Glucose measurement, fasting
C0202045|Glucose measurement, fasting (procedure)
C0202045|fasting glucose test
C0202045|Test;glucose;fasting
C0202046|Glucose measurement, random
C0202046|Glucose measurement, random (procedure)
C0202046|random glucose test
C0202046|Test;glucose;random
C0017741|Glucose Tolerance Test
C0017741|Glucose Tolerance Tests
C0017741|Test;glucose tolerance
C0017741|Glucose tolerance test (GTT)
C0017741|Blood glucose (sugar) tolerance test
C0017741|Glucose tolerance test NOS
C0017741|Glucose tolerance test NOS (procedure)
C0017741|GTT
C0017741|GTT - Glucose tolerance test
C0017741|OGTT - Oral glucose tolerance test
C0017741|Glucose challenge test
C0017741|Glucose tolerance test (procedure)
C0017741|Glucose tolerance test, NOS
C0523657|Glucose measurement, tolbutamide tolerance test
C0523657|Glucose measurement, tolbutamide tolerance test (procedure)
C1272314|Fecal clinitest (procedure)
C1272314|Faecal clinitest (procedure)
C1272314|Faecal clinitest
C1272314|Fecal clinitest
C0427743|Glucose concentration
C0427743|Glucose concentration, test strip measurement (procedure)
C0427743|Glucose concentration, test strip measurement
C1295145|Glucose measurement estimated from glycated haemoglobin
C1295145|Glucose measurement estimated from glycated hemoglobin (procedure)
C1295145|Glucose measurement estimated from glycated hemoglobin
C0428549|Fluid sample glucose measurement
C0428549|body fluid glucose measurement (lab test)
C0428549|body fluid glucose
C0428549|body fluid glucose measurement
C0428549|Measurement of glucose in body fluid
C0428549|Body Fluid Glucose Test
C0428549|Fluid sample glucose level
C0428549|Fluid sample glucose measurement (procedure)
C0428549|Glucose measurement, body fluid
C1319276|Faecal glucose level
C1319276|Faecal glucose measurement
C1319276|Fecal glucose level (procedure)
C1319276|Fecal glucose level
C1319276|Fecal glucose measurement
C2732844|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 120 minutes after 75 gram oral glucose challenge (procedure)
C2732844|Quantitative measurement of glucose in serum or plasma specimen 120 minutes after 75 gram oral glucose challenge
C2732844|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 120 minutes after 75 gram oral glucose challenge
C2733143|Quantitative measurement of substance rate of glucose excretion in urine specimen
C2733143|Quantitative measurement of substance rate of glucose excretion in urine
C2733143|Quantitative measurement of substance rate of glucose excretion in urine specimen (procedure)
C2732700|Quantitative measurement of mass concentration of glucose in pericardial fluid specimen (procedure)
C2732700|Quantitative measurement of mass concentration of glucose in pericardial fluid specimen
C2732700|Quantitative measurement of glucose in pericardial fluid specimen
C2732794|Quantitative measurement of mass concentration of glucose in 1 hour postprandial urine specimen (procedure)
C2732794|Quantitative measurement of mass concentration of glucose in 1 hour postprandial urine specimen
C2732794|Quantitative measurement of glucose in 1 hour postprandial urine specimen
C2732897|Quantitative measurement of glucose in peritoneal dialysis fluid specimen
C2732897|Quantitative measurement of mass concentration of glucose in peritoneal dialysis fluid specimen
C2732897|Quantitative measurement of mass concentration of glucose in peritoneal dialysis fluid specimen (procedure)
C2732804|Quantitative measurement of mass concentration of glucose in synovial fluid specimen
C2732804|Quantitative measurement of glucose in synovial fluid specimen
C2732804|Quantitative measurement of mass concentration of glucose in synovial fluid specimen (procedure)
C2733070|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 6 hours after glucose challenge
C2733070|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 6 hours after glucose challenge (procedure)
C2733070|Quantitative measurement of glucose in serum or plasma specimen 6 hours after glucose challenge
C2732796|Quantitative measurement of mass rate of excretion of glucose in 24 hour urine specimen
C2732796|Quantitative measurement of mass rate of excretion of glucose in 24 hour urine specimen (procedure)
C2732796|Quantitative measurement of glucose in 24 hour urine specimen
C2732716|Quantitative measurement of mass concentration of glucose in postcalorie fasting serum or plasma specimen
C2732716|Quantitative measurement of mass concentration of glucose in postcalorie fasting serum or plasma
C2732716|Quantitative measurement of mass concentration of glucose in postcalorie fasting serum or plasma specimen (procedure)
C2732249|Quantitative measurement of mass concentration of glucose in pleural fluid specimen (procedure)
C2732249|Quantitative measurement of mass concentration of glucose in pleural fluid specimen
C2732249|Quantitative measurement of glucose in pleural fluid specimen
C2711175|Measurement of fasting glucose in urine specimen using dipstick
C2711175|Measurement of fasting glucose in urine specimen using dipstick (procedure)
C2188672|urine fasting glucose measurement
C2188672|urine fasting glucose measurement (lab test)
C2188672|urine glucose fasting
C2188672|glucose, fasting, urine
C2188672|urine fasting glucose
C0428568|fasting blood glucose measurement (lab test)
C0428568|fasting blood glucose measurement
C0428568|blood glucose fasting
C0428568|fasting blood glucose
C0428568|Fasting blood glucose (& level)
C0428568|Fasting blood glucose (& level) (procedure)
C0428568|Fasting blood glucose level
C0428568|Fasting blood glucose level (procedure)
C0428568|FBS - Fasting blood sugar
C0428568|FBG - Fasting blood glucose
C0428568|Fasting blood glucose measurement (procedure)
C2238123|fasting whole blood glucose measurement
C2238123|fasting whole blood glucose measurement (lab test)
C2238123|glucose, fasting, whole blood
C2238123|fasting whole blood glucose
C2238123|whole blood fasting glucose
C2317664|fasting fingerstick blood glucose
C2317664|fasting fingerstick blood glucose measurement
C2317664|fingerstick blood glucose fasting
C2317664|fasting fingerstick blood glucose measurement (lab test)
C4028983|footstick blood glucose fasting (lab test)
C4028983|footstick blood glucose fasting
