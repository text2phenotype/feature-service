C0419735|patient immune to hepatitis A
C0419735|patient immune to Hep A
C0419735|patient vaccinated for Hep A
C1170008|hepatitis A and hepatitis B vaccine                                                                            
C0419735|Hepatitis A immunization (SNOMED:243789007)
C3644200|Hepatitis A immune globulin                                                                                
C3526526|hepatitis A vaccine, adult dosage                                                                             
C0694731|hepatitis A vaccine, pediatric dosage, unspecified formulation                                                               
C1548491|hepatitis A vaccine, pediatric/adolescent dosage, 2 dose schedule                                                             
C1548492|hepatitis A vaccine, pediatric/adolescent dosage, 3 dose schedule                                                             
C3644157|hepatitis A vaccine, unspecified formulation
C3526526|Hep A, adult                                                                                        
C3644200|Hep A, IG                                                                                         
C1548491|Hep A, ped/adol, 2 dose                                                                                  
C1548492|Hep A, ped/adol, 3 dose                                   
C0694731|Hep A, pediatric, unspecified formulation                                                                         
C3644157|Hep A, unspecified formulation
C1170008|Hep A-Hep B
C0730242|combined hepatitis a & hepatitis b vaccination
C0730242|combined hepatitis A and hepatitis B vaccination (medication)
C0730242|combined hepatitis A and hepatitis B vaccination
C0730242|Combined hepatitis A and B vaccination
C0730242|Combined hepatitis A and B vaccination (procedure)
C1281986|Hepatitis A and typhoid vaccination (procedure)
C1281986|Hepatitis A and typhoid vaccination
C0419735|Immunisation;hepatitis A
C0419735|Hepatitis A immunization
C0419735|Hepatitis A immunisation
C0419735|Hepatitis A immunisation (procedure)
C0419735|hepatitis a vaccine administration (medication)
C0419735|hepatitis a vaccine administration
C0419735|Hepatitis A vaccination
C0419735|Hepatitis A vaccination, unspecified
C0419735|Hepatitis A immunization (procedure)
C0419735|Immunization;hepatitis A
C0419736|First hepatitis A vaccination (procedure)
C0419736|First hepatitis A vaccination
C0419736|First hepatitis A vaccination (medication)
C0419736|hepatitis a vaccines first vaccination
C0419736|1st hepatitis A vaccination
C0419737|Second hepatitis A vaccination
C0419737|Second hepatitis A vaccination (procedure)
C0419737|Second hepatitis A vaccination (medication)
C0419737|hepatitis a vaccines second vaccination
C0419737|2nd hepatitis A vaccination
C0419739|Booster hepatitis A vaccination
C0419739|Booster hepatitis A vaccination (procedure)
C0419738|Third hepatitis A vaccination
C0419738|Third hepatitis A vaccination (procedure)
C0419738|3rd hepatitis A vaccination
C1170689|Twinrix Junior
C1170008|Hepatitis A and hepatitis B vaccine
C1170008|Hep A-Hep B
C1170008|hepatitis A-hepatitis B vaccine
C3644200|Hep A, IG
C3644200|Hepatitis A immune globulin
C3526526|Hepatitis A vaccine, adult dosage
C3526526|Hep A, adult
C0694731|Hep A, pediatric, unspecified formulation
C0694731|hepatitis A vaccine, pediatric dosage, unspecified formulation
C0694731|Hep A, pediatric, NOS
C1548491|Hep A, ped/adol, 2 dose
C1548491|hepatitis A vaccine, pediatric/adolescent dosage, 2 dose schedule
C1548492|hepatitis A vaccine, pediatric/adolescent dosage, 3 dose schedule
C1548492|Hep A, ped/adol, 3 dose
C3644157|Hep A, unspecified formulation
C3644157|hepatitis A vaccine, unspecified formulation
