C1399448|Birth to an HCV-infected mother
C1399448|Born with HCV
C1399448|Mother has HCV
C1399448|Mother had HCV
C1399448|maternal; hepatitis, affecting fetus
C1399448|hepatitis; maternal, affecting fetus
C1399448|maternal; hepatitis, affecting fetus
