C0030705|T101|Patient|
C0030705|T101|Patients|
C0030705|T101|PT|
C0030705|T101|*^patient|
C0030705|T101|^Patient|
C0030705|T101|LAY USER/PATIENT|
C0030705|T101|Patient (person)|
C0037125|T196|Silver|
C0037125|T196|Ag|
C0037125|T196|Silver [Chemical/Ingredient]|
C0037125|T196|Ag element|
C0037125|T196|Ag - Silver|
C0037125|T196|Silver (substance)|
C0037125|T196|Silver, NOS|
C1514241|T033|Positive|
C1514241|T033|Positive Finding|
C0006826|T191|Cancer|
C0006826|T191|Cancers|
C0006826|T191|Malignant neoplasm without specification of site|
C0006826|T191|Malignant Neoplasms|
C0006826|T191|CA|
C0006826|T191|Malignant neoplastic disease|
C0006826|T191|malignant neoplasm|
C0006826|T191|unspecified malignant neoplasm|
C0006826|T191|malignant neoplasm (diagnosis)|
C0006826|T191|cancer, NOS|
C0006826|T191|unspecified malignant neoplasm (diagnosis)|
C0006826|T191|Cancer NOS|
C0006826|T191|Malignancy|
C0006826|T191|neoplasm/cancer|
C0006826|T191|CA - Cancer|
C0006826|T191|Malignant neoplasm of unspecified site NOS (disorder)|
C0006826|T191|Malignant neoplasm of unspecified site|
C0006826|T191|Malignant tumor|
C0006826|T191|Malignant neoplasm of unspecified site (disorder)|
C0006826|T191|Malignant tumour|
C0006826|T191|Ca - unspecified site NOS|
C0006826|T191|Ca - unspecified site|
C0006826|T191|[X]Malignant neoplasm without specification of site|
C0006826|T191|Malignant neoplasm NOS|
C0006826|T191|Ca - unspecified site NOS (disorder)|
C0006826|T191|(Neoplasms) or (cancers) (disorder)|
C0006826|T191|Neoplasms - malignant|
C0006826|T191|[X]Malignant neoplasm without specification of site (disorder)|
C0006826|T191|Malignant tumour (disorder)|
C0006826|T191|(Neoplasms) or (cancers)|
C0006826|T191|Malignant neoplasm of unspecified site NOS|
C0006826|T191|NEOPLASM, MALIGNANT|
C0006826|T191|Malignant Growth|
C0006826|T191|Neoplasm malignant|
C0006826|T191|Cancer (NOS)|
C0006826|T191|Med: Malignant neoplastic disease|
C0006826|T191|Malignant neoplastic disease (disorder)|
C0006826|T191|tumor; malignant, unclassified|
C0006826|T191|tumor; unclassified, malignant|
C0006826|T191|Malignant tumor (disorder)|
C0006826|T191|Cancer, unspecified site|
C0006826|T191|Malignancy, unspecified site|
C1261327|T033|Family history: Asthma (context-dependent category)|
C1261327|T033|Family history: Asthma (situation)|
C1261327|T033|Family history: Asthma|
C1261327|T033|FH: Asthma (situation)|
C1261327|T033|FH: Asthma|
C1261327|T033|Family history of asthma|
C1261327|T033|family history; asthma|
C1261327|T033|history; family, with asthma|
C0032854|T102|Poverty|
C0032854|T102|Poverty status|
C0032854|T102|Low Income|
C0032854|T102|Poor|
C0032854|T102|Financially poor|
C0032854|T102|Financially poor (finding)|
C0032854|T102|Social problem - poverty|
C0032854|T102|Economic deprivation|
C0032854|T102|Pauper|
C0032854|T102|Severe lack of money|
C0032854|T102|Living in poverty|
C0007457|T098|Caucasoid Race|
C0007457|T098|white race|
C0007457|T098|racial background Caucasian|
C0007457|T098|racial background Caucasian (history)|
C0007457|T098|Race: Caucasian|
C0007457|T098|Caucasian race|
C0007457|T098|Race: Caucasian (racial group)|
C0007457|T098|Race: Caucasian (finding)|
C0007457|T098|Race: White|
C0007457|T098|Caucasoid|
C0007457|T098|WHITE|
C0007457|T098|Caucasian Races|
C0007457|T098|Caucasoid Races|
C0007457|T098|Race, Caucasian|
C0007457|T098|Race, Caucasoid|
C0007457|T098|Races, Caucasian|
C0007457|T098|Races, Caucasoid|
C0007457|T098|Caucasian|
C0007457|T098|Whites|
C0007457|T098|Caucasians|
C0007457|T098|Occidental|
C0007457|T098|Caucasian (racial group)|
C0043157|T098|Caucasians|
C0043157|T098|caucasian|
C0043157|T098|RaceWhite|
C0043157|T098|Caucasian (living organism) (ethnic group)|
C0043157|T098|White - ethnic group (ethnic group)|
C0043157|T098|White - ethnic group|
C0043157|T098|White|
C0043157|T098|White/Caucasian|
C0043157|T098|Whites|
C0043157|T098|Caucasoid|
C0043157|T098|Caucasian (ethnic group)|
C0043157|T098|Caucasian, NOS|
C0043157|T098|Caucasian (living organism)|
C0424670|T033|Weight for height|
C0424670|T033|Weight for height (observable entity)|
C0424670|T033|Ponderal index|
C0013146|T048|Abuse, Drug|
C0013146|T048|drug abuse|
C0013146|T048|Recreational drug use|
C0013146|T048|rndx drug abuse|
C0013146|T048|rndx drug abuse (diagnosis)|
C0013146|T048|Abuse;drug(s)|
C0013146|T048|Medication abuse|
C0013146|T048|substance abuse drug|
C0013146|T048|drug abuse (diagnosis)|
C0013146|T048|Drugs of abuse|
C0013146|T048|Drug abuse NOS|
C0013146|T048|Drug abuse (disorder)|
C0013146|T048|disorder, drug abuse|
C0013146|T048|abuse; drugs|
C0013146|T048|Drug abuse, NOS|