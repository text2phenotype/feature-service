C0002059|Alkaline Phosphatase
C0201850|Alkaline phosphatase measurement
C0050528|acetylphosphatase
C0073127|retinyl phosphatase
C0061565|beta-glycerophosphatase
C0061565|glycerol-2-phosphatase
C0061565|Glycerol 2-phosphatase
C0061565|Glycerol 2-phosphatase (substance)
C0061952|guanidinodeoxy-scyllo-inositol-4-phosphatase
C0061952|Guanidinodeoxy-scyllo-inositol-4-phosphatase (substance)
C0065665|mannitol-1-phosphatase
C0065665|Mannitol-1-phosphatase (substance)
C0070862|phosphoglycerate phosphatase
C0070862|Phosphoglycerate phosphatase (substance)
C0070943|phosphoserine phosphatase
C0070943|Choline phosphatase
C0070943|L-3-phosphoserine-phosphatase
C0070943|Phosphoserine phosphatase (substance)
C0072710|pyridoxal-5-phosphatase
C0075313|streptomycin-6-phosphatase
C0075313|Streptomycin-6-phosphatase (substance)
C0076406|thiamine monophosphatase
C0077558|tyrosine phosphate hydrolase
C0065687|mannose-6-phosphatase
C0070891|phosphonate esterase
C0062678|hexose phosphatase
C0060773|Fructose-2,6-bisphosphatase
C0060773|FRUCTOSE BISPHOSPHATASE 02 06
C0060773|fructose-2,6-diphosphatase
C0060773|Fructose 2,6-bisphosphatase
C0060773|Fructose-2,6-bisphosphate 2-phosphatase
C0060773|Fructose-2,6-bisphosphatase (substance)
C0060774|fructose-6-phosphatase
C0061563|glycerol-1-phosphatase
C0061563|Glycerol-1-phosphatase (substance)
C0284786|capping enzyme, Artemia salina
C0070941|phosphorylphosphatase
C0070946|phosphothreonine phosphatase
C0136841|phosphocholine phosphatase
C0245367|glyceraldehyde 3-phosphate phosphatase
C0171000|lysophosphatidic acid phosphatase
C0251880|glucose-3-phosphatase
C0259479|polyphosphoinositide phosphatase
C0060776|PHOSPHOFRUCTOKINASE FRUCTOSE BISPHOSPHATASE 002 006
C0060776|Fru-kinase-Fru-bisphosphatase
C0060776|F Kinase-F-bisphosphatase
C0060776|6-Phosphofructo 2-kinase-fructose 2,6-bisphosphatase
C0060776|Fructose-6-phosphate,2-kinase-fructose-2,6-bisphosphatase
C0060776|6-PF-2-K-Fru-2,6-P(2)ase
C0060776|6-Phosphofructo-2-kinase-fructose-2,6-bisphosphatase
C0384935|phosphonoacetate hydrolase
C0384935|Phosphonoacetate hydrolase (substance)
C0384935|phnA protein
C0385927|synaptojanin
C0385927|synaptojanin-1
C0385927|synaptojanin1
C0536328|glucosylglycerol-phosphate phosphatase
C0443450|Alk. phos. - bile isoenzyme
C0443450|Alkaline phosphatase biliary isoenzyme
C0443450|Alkaline phosphatase biliary isoenzyme (substance)
C0061401|Glc-1,6-P(2) phosphatase
C0061401|glucose 1,6-bisphosphatase
C0061401|glucose 1,6-diphosphate phosphatase
C0061401|glucose bisphosphatase
C0070830|PDMase
C0070830|phosphodiesterase-phosphomonoesterase
C0070830|PDM phosphatase
C0106564|bisphosphoglycerate synthase-phosphatase
C0053804|bisphosphoglycerate phosphatase
C0053804|diphosphoglycerate phosphatase
C0053804|glycerate-2,3-P2 phosphatase
C0053804|Bisphosphoglycerate phosphatase (substance)
C0119666|glycerate-2,3-P2 synthase
C0140297|retinyl monophosphate phosphatase
C0163342|1L-myo-inositol-1-phosphatase
C0163342|1L-myo-inositol-1-phosphate phosphohydrolase
C0163342|inositol phosphatase
C0163342|inositol-1-phosphate phosphohydrolase
C0163342|myo-inositol monophosphatase
C0163342|myo-inositol-1-phosphatase
C0163342|inositol monophosphatase
C0163342|myo-inositol-1 (or 4)-monophosphatase
C0163342|1L-myo-Inositol-1-phosphatase (substance)
C0163342|inositol monophosphate phosphatase impA
C0121682|hexose-6-phosphate phosphohydrolase
C0145597|thiamine phosphate phosphatase
C0243811|phosphatidyl-inositol-bisphosphate phosphatase
C0243811|phosphatidylinositol 4,5-bisphosphate phosphomonoesterase
C0243811|triphosphoinositide phosphatase
C0243811|Phosphatidylinositol-bisphosphatase
C0243811|type IV 5-phosphatase
C0243811|phosphoinositide 5-phosphatase
C0243811|phospholipid-specific inositol polyphosphate 5-phosphatase
C0243811|inositol polyphosphate 5-phosphatase type IV
C0243811|ptdIns(4,5)P2 5-phosphatase
C0243811|phosphatidylinositol-4,5-bisphosphate-5-phosphatase
C0243811|Phosphatidylinositol-bisphosphatase (substance)
C0076951|trehalose-6-phosphate phosphatase
C0076951|trehalose-6-phosphate phosphohydrolase
C0076951|trehalose-phosphatase
C0076951|Trehalose-phosphatase (substance)
C0147378|tyrosine-o-phosphate phosphatase
C0077893|UMPase
C0077893|uridine monophosphatase
C0147902|uridine monophosphatase-2
C0243858|2-keto-3-deoxyoctonate-8-phosphate phosphatase
C0243858|3-deoxy-D-manno-octulosonate 8-phosphate phosphatase
C0243858|KDO-8-phosphatase
C0243858|3-deoxy-manno-octulosonate-8-phosphatase
C0243858|3-Deoxy-manno-octulosonate-8-phosphatase (substance)
C0070792|PGPase
C0070792|phosphatidylglycerolphosphate phosphatase
C0070792|phosphatidylglycerophosphatase
C0070792|Phosphatidylglycerophosphatase (substance)
C0072718|pyridoxal phosphate phosphatase
C0072718|pyridoxal-P hydrolase
C0072718|pyridoxamine phosphate phosphatase
C0072718|pyridoxamine-P hydrolase
C0072718|pyridoxine phosphate phosphatase
C0072718|vitamin B(6)-phosphate phosphatase
C0046855|3'-phosphoadenosine-5'-phosphosulfate phosphohydrolase
C0046855|PAPS phosphohydrolase
C0148536|VITF-A
C0126638|m-RNA guanylyltransferase.RNA (guanine-7) methyltransferase
C0129120|mRNA capping enzyme, Shope Fibroma virus
C0063589|inositol triphosphate phosphatase
C0063589|inositol triphosphate phosphomonoesterase
C0063589|INTP esterase
C0063589|triphosphoinositide phosphomonoesterase
C0119679|glycerol-3-phosphatase
C0067046|I-P3ase
C0067046|inositol 1,4,5-triphosphate phosphatase
C0067046|myo-inositol 1,4,5-triphosphate phosphatase
C0134093|organophosphate hydrolase
C0244922|1-alkyl-2-acetyl-sn-glycero-3-phosphate phosphohydrolase
C0244922|alkylacetyl-GP phosphohydrolase
C0244922|alkylacetylglycerophosphatase
C0244922|Alkylacetylglycerophosphatase (substance)
C0088353|1,4,5-triphosphate-1,2,4,5-tetrakisphosphate 5-phosphatase
C0088353|inositol-polyphosphate 5-phosphatase
C0088353|inositol polyphosphate 5-phosphatase
C0088353|inositol 5-phosphatase
C0088353|IP3-5-phosphatase
C0088353|inositol-1,4,5-trisphosphate 5-phosphatase
C0088353|inositol triphosphatase
C0088353|myoinositol trisphosphatase
C0088353|inositol-1,4,5-trisphosphate 5'-phosphatase
C0088353|Ins(1,4,5)P3 5'-phosphatase
C0088353|Inpp5f protein, mouse
C0088353|inositol triphosphate 5-phosphatase
C0083008|inositol 1,3,4,5-tetrakisphosphate 3-phosphomonoesterase
C0083008|Ins(1,3,4,5)P4 3-phosphatase
C0083008|inositol 1,3,4,5-polyphosphate 5-phosphatase
C0083008|inositol 1,3,4,5-tetrakisphosphate 3-phosphatase
C0083008|inositol tetrakisphosphate phosphomonoesterase
C0083008|inositol 1,3,4,5-tetrakisphosphate phosphomonoesterase
C0083008|Ins(1,3,4,5)P4 phosphomonoesterase
C0083008|multiple inositol-polyphosphate phosphatase
C0083008|Ins(1,3,4,5)P4 5-phosphatase
C0083008|Inositol-1,3,4,5-tetrakisphosphate 3-phosphatase (substance)
C0083008|Inositol-1,3,4,5-tetrakisphosphate 3-phosphatase
C0083008|MIPP enzyme
C0083008|multiple inositol polyphosphate phosphatase
C0066978|mutT protein, E coli
C0208628|D-myo-inositol (1,4)-bisphosphate 1-phosphatase
C0208628|inositol bisphosphatase
C0208628|inositol polyphosphate 1-phosphatase
C0208628|inositol-1,4-bisphosphate-1-phosphatase
C0208628|IP2 1-phosphatase
C0208628|myoinositol diphosphatase
C0208628|inositol-1,4-bisphosphate 1-phosphatase
C0208628|Inositol-1,4-bisphosphate 1-phosphatase (substance)
C0063566|inositol 1,3,4-triphosphate 4-phosphatase
C0063566|INTP 4-phosphatase
C0063566|phosphatidylinositol-3,4-bisphosphate 4-phosphatase
C0063566|PtdIns(3,4)P2 4-phosphatase
C0063566|PTDINS-4P-phosphatase
C0063566|phosphatidylinositol 4-phosphatase
C0063566|inositol polyphosphate 4-phosphatase
C0063566|Ins polyP 4-phosphatase
C0063566|ptdIns4P monoesterase
C0063566|phosphatidylinositol-4-phosphate monoesterase
C0063566|inositol 1,3,4-trisphosphate 4-phosphatase
C0063566|phosphatidylinositol 4-phosphate phosphatase
C0057631|dGTPase
C0057631|Deoxy-GTPase
C0057631|dGTPase (substance)
C0245366|GLPH phosphatase
C0638832|INTP 3-phosphatase
C0638832|inositol polyphosphate 3-phosphatase
C0638832|phosphatidylinositol 3-phosphatase
C0638832|phosphatidylinositol-3-phosphatase
C0638832|Phosphatidylinositol-3-phosphatase (substance)
C0061413|Glucose-1-phosphatase
C0061413|glucose 1 phosphatase
C0061413|agp protein, E coli
C0061413|glucose-1-phosphatase, E coli
C0061413|Glucose-1-phosphatase (substance)
C0123583|1,3,4,5,6-InsP5-1-3-phosphatase
C0123583|inositol 1,3,4,5,6-pentakisphosphate-1-3-phosphatase
C0210507|8-oxo-deoxy-GTPase
C0210507|8-oxodGTPase
C0210507|8-oxo-dGTPase
C0210507|8-oxo-7,8-dihydroguanosine triphosphatase
C0210507|7,8-Dihydro-8-Oxoguanine Triphosphatase
C0210507|Nucleoside Diphosphate-Linked Moiety X Motif 1
C0210507|Nudix Motif 1
C0210507|8-oxo-2'-deoxyguanosine 5'-triphosphate pyrophosphohydrolase
C0210507|2-Hydroxy-dATP Diphosphatase
C0210507|EC 3.6.1.56
C0210507|EC 3.6.1.55
C0247876|Cer-1-P phosphatase
C0247876|ceramide-1-phosphate phosphatase
C0251087|FDP 6-phosphatase
C0251087|Fru(2,6)P2 6-phosphatase
C0251087|fructose-2,6-bisphosphate 6-phosphatase
C0251087|Fructose-2,6-bisphosphate 6-phosphatase (substance)
C1430004|MutX protein, Streptococcus pneumoniae
C0259478|PPI phosphatase
C0295334|NPtase
C0295334|Staphylococcal NPtase
C0295334|Staphylococcal neutral phosphatase
C0295334|NPase, S. aureus
C0295334|neutral phosphatase, S. aureus
C0297587|2-deoxyglucose-6-phosphate phosphatase
C0297587|2-deoxyglucose-6-phosphatase
C0297587|2-deoxyglucose-6-phosphatase (substance)
C0300570|2-keto-3-deoxyoctulosonate-activated 4'-phosphatase
C0300570|KDO-activated lipid A 4'-phosphatase
C0300570|lipid A 4'-phosphatase
C0382361|PI(3,4,5)P3 5-Pase
C0382361|PtdIns(3,4,5)P3 5-phosphatase
C0382361|phosphatidylinositol-3,4,5-trisphosphate 5-phosphatase
C0388055|SHIP2 protein, human
C0388055|inositol polyphosphate phosphatase-like 1 protein, human
C0388055|INPPL1 protein, human
C0390960|2-carboxyarabinitol 1-phosphate phosphatase
C0390960|CA1P phosphatase
C0390960|CA1Pase
C0528468|PIP(2) phosphatase
C0528937|PHON1protein, Shigella flexneri
C0301810|Alkaline phosphatase isoenzymes
C0301810|Alkaline phosphatase isoenzyme
C0301810|Alkaline phosphatase isoenzyme (substance)
C0301810|Alkaline phosphatase isoenzyme, NOS
C0134983|Intestine Alkaline Phosphatase
C0312399|Alkaline phosphatase isoenzyme, bone fraction
C0312399|Alkaline phosphatase.bone
C0312399|Bone Specific Alkaline Phosphatase
C0312399|Bone Alkaline Phosphatase
C0312399|Bone-Specific Alkaline Phosphatase
C0312399|BSAP
C0312399|BAP
C0312399|Alkaline Phosphatase, Bone Specific
C0312399|bALP
C0312399|Alkaline phosphatase bone isoenzyme
C0312399|Alkaline phosphatase isoenzyme, bone fraction (substance)
C0312398|Alkaline phosphatase.liver
C0312398|Alk. phos. - liver isoenzyme
C0312398|Liver Alkaline Phosphatase
C0312398|Alkaline phosphatase isoenzyme, liver fraction
C0312398|Alkaline phosphatase liver isoenzyme
C0312398|Alkaline phosphatase isoenzyme, liver fraction (substance)
C0002059|Alkaline Phosphatase
C0002059|Orthophosphoric-monoester phosphohydrolase (alkaline optimum)
C0002059|AP
C0002059|alkaline phosphomonoesterase
C0002059|glycerophosphatase
C0002059|Alkaline Phosphatase [Chemical/Ingredient]
C0002059|Phosphomonoesterase
C0002059|ALP - Alkaline phosphatase
C0002059|AP - Alkaline phosphatase
C0002059|Alkaline phosphatase (substance)
C0740201|alkaline phosphatase Regan isoenzyme
C0740201|placental-like Regan isoenzyme
C0740201|Regan isoenzyme
C0740201|ALPP
C0740201|Alkaline phosphatase.regan
C0740201|alkaline phosphatase, placental
C0740201|placental alkaline phosphatase isoenzyme
C0740201|Reagan isoenzyme
C0740201|Regan isoenzyme (substance)
C2932888|ALPL protein, human
C2932888|alkaline phosphatase, liver-bone-kidney, human
C2932888|TNSALP protein, human
C2932888|TNAP phosphatase, human
C2932888|tissue-non specific alkaline phosphatase, human
C2932888|Liver/Bone/Kidney-Type Alkaline Phosphatase
C2932888|Glycerophosphatase
C2932888|Alkaline Phosphatase, Tissue-Nonspecific Isozyme
C2932888|Tissue-Nonspecific ALP
C2932888|EC 3.1.3.1
C2932888|Alkaline Phosphomonoesterase
C2932890|ALPPL2 protein, human
C2932890|alkaline phosphatase Nagao isozyme, human
C2932890|alkaline phosphatase, placental-like, human
C1318717|Alkaline phosphatase
C1318717|Alkaline phosphatase stain (substance)
C1318717|Alkaline phosphatase stain
C1980989|Alkaline phosphatase &#124; peritoneal fluid
C1980989|Alkaline phosphatase &#x7C; peritoneal fluid
C1980987|Alkaline phosphatase &#x7C; body fluid
C1980991|Alkaline phosphatase &#x7C; urine
C1980986|Alkaline phosphatase &#x7C; bld-ser-plas
C2703301|Alkaline phosphatase &#x7C; Amniotic Fluid
C2737363|Alkaline phosphatase &#x7C; Blood cord
C2924679|Alkaline phosphatase &#x7C; Dialysis fluid
C1980990|Alkaline phosphatase &#x7C; Tissue and Smears
C3490795|asfotase alfa
C3490795|asfotase alfa (medication)
C3490795|enzyme replenishers asfotase alfa
C2930591|ALPP protein, human
C2930591|alkaline phosphatase, placental (Regan isozyme), human
C2930591|Alkaline phosphatase Regan isozyme, human
C2930591|Alkaline Phosphomonoesterase
C2930591|Alkaline Phosphatase Regan Isozyme
C2930591|EC 3.1.3.1
C2930591|Alkaline Phosphatase, Placental Type
C2930591|PLAP-1
C2930591|Placental Alkaline Phosphatase 1
C2930591|Regan Isozyme
C1307712|alkaline protease AprP, Pseudomonas
C1307712|AprP protease, Pseudomonas
C1148297|Alkaline phosphatase.heat stable
C1148297|Heat stable alkaline phosphatase (substance)
C1148297|Heat stable alkaline phosphatase
C1148296|Alkaline phosphatase.heat labile
C1148296|Heat labile alkaline phosphatase
C1148296|Heat labile alkaline phosphatase (substance)
C4040565|Macro alkaline phosphatase
C4040565|Macro alkaline phosphatase (substance)
C4041728|alkaline phosphatase, liver-bone-kidney, mouse
C4041728|ALPL protein, mouse
C0625821|progesterone 11-glucuronide-alkaline phosphatase conjugate
C0625821|progesterone-G-AP
C0061237|germ-cell AP isoenzyme
C0061237|Nagao isoenzyme
C0061237|placental-like alkaline phosphatase
C0061237|PLAP-like AP
C1447085|ALPI protein, human
C1447085|alkaline phosphatase, intestinal, human
C1447085|intestinal alkaline phosphatase, human
C1447085|p75-150 antigen, human
C0529894|miniPLAP
C0529894|miniplacental alkaline phosphatase
C0671822|MC14 alkaline phosphatase I
C0671822|MC14 APase I
C0961931|alkaline phosphatase, intestinal, rat
C0961931|intestinal alkaline phosphatase-I, rat
C0961931|Alpi protein, rat
C0961931|r-IAP-I
C0961932|intestinal alkaline phosphatase-II, rat
C0961932|alkaline phosphatase 3, intestine, not Mn requiring protein, rat
C0961932|Akp3 protein, rat
C0961932|alpi2 protein, rat
C0961932|r-IAP-II
C1100624|MUSEAP protein, mouse
C1120950|PafA enzyme
C1120950|periplasmic alkaline phosphatase, Chryseobacterium meningosepticum
C1120950|PafA protein, Chryseobacterium meningosepticum
C1721792|PHO8 protein, S cerevisiae
C1722357|Akp-2 protein, mouse
C1722357|Akp2 protein, mouse
C1722357|alkaline phosphatase 2, mouse
C1722357|tissue-specific alkaline phosphatase, mouse
C1739750|b0383 protein, E coli
C1739750|ECK0378 protein, E coli
C1739750|phoA protein, E coli
C1958108|alkaline phosphatase 3, mouse
C1958108|alkaline phosphatase 3, intestine, not Mn requiring protein, mouse
C1958108|Akp3 protein, mouse
C0201850|Alkaline phosphatase measurement
C0201850|Phosphatase, alkaline
C0201850|ALP
C0201850|Test;alkaline phosphatase
C0201850|Measurement of alkaline phosphatase
C0201850|ASSAY OF PHOSPHATASE ALKALINE
C0201850|Alkaline Phosphatase
C0201850|ALK phosph
C0201850|Alk phos
C0201850|Alkaline phosphatase measurement (procedure)
C0201850|ASSAY ALKALINE PHOSPHATASE
C0201850|alkaline phosphatase test
C0036776|serum alkaline phosphatase
C0036776|SAP
C0036776|Serum Alkaline Phosphatase Measurement
C0036776|serum alkaline phosphatase measurement (lab test)
C0036776|Serum alkaline phosphatase (& level)
C0036776|Serum alkaline phosphatase (& level) (procedure)
C0036776|Alk. phosphatase -serum
C0036776|Alkaline phosphatase (& level (& serum))
C0036776|Phosph.- alk. - serum
C0036776|Serum alkaline phosphatase NOS
C0036776|Alkaline phosphatase (& level (& serum)) (procedure)
C0036776|Serum alkaline phosphatase NOS (procedure)
C0036776|Serum Alkaline Phosphatase Test
C0036776|Serum alkaline phosphatase level
C0036776|Serum alkaline phosphatase measurement (procedure)
C1293930|Measurement of ratio of analyte to alkaline phosphatase (procedure)
C1293930|Measurement of ratio of analyte to alkaline phosphatase
C0201851|Phosphatase, alkaline; isoenzymes
C0201851|Measurement of alkaline phosphatase isoenzymes
C0201851|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|Alkaline phosphatase isoenzymes measurement
C0201851|Alkaline phosphatase isoenzymes measurement (procedure)
C0201851|ASSAY ALKALINE PHOSPHATASES
C0201855|Alkaline phosphatase, heat stable measurement
C0201855|Phosphatase, alkaline; heat stable (total not included)
C0201855|Measurement of heat stable alkaline phosphatase
C0201855|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|Thermostable alkaline phosphatase measurement
C0201855|Alkaline phosphatase, heat stable measurement (procedure)
C0201855|ASSAY ALKALINE PHOSPHATASE
C2984961|Bone Specific Alkaline Phosphatase Measurement
C2984961|Bone Alkaline Phosphatase Measurement
C2984961|Bone Specific Alkaline Phosphatase
C2984961|ALPBS
C2984961|Bone ALP Measurement
C3898585|Liver Specific Alkaline Phosphatase Measurement
C3898585|ALPLS
C3898585|Liver Specific Alkaline Phosphatase
C3898710|Intestinal Specific Alkaline Phosphatase
C3898710|ALPIS
C3898710|Intestinal Specific Alkaline Phosphatase Measurement
C0200697|Leukocyte alkaline phosphatase level
C0200697|Leucocyte alkaline phosphatase level
C0200697|Leucocyte alkaline phosphatase level (procedure)
C0200697|Leukocyte alkaline phosphatase score
C0200697|Leucocyte alkaline phosphatase score
C0200697|Leukocyte alkaline phosphatase score (procedure)
C0200697|Leukocyte alkaline phosphatase score (observable entity)
C0200697|Neutrophil alkaline phosphatase score
C0200697|LAP score
C0200697|LAP - Neutrophil alkaline phosphatase score
C0200697|LAP - Neutrophil alkaline phosphatase score measurement
C0201852|Placental alkaline phosphatase measurement
C0201852|PLAP measurement
C0201852|Placental alkaline phosphatase measurement (procedure)
C0201853|Intestinal alkaline phosphatase measurement
C0201853|IAP measurement
C0201853|Intestinal alkaline phosphatase measurement (procedure)
C0201854|Germ cell alkaline phosphatase measurement
C0201854|GCAP measurement
C0201854|Germ cell alkaline phosphatase measurement (procedure)
C0428333|Fluid sample alkaline phosphatase level
C0428333|Fluid sample alkaline phosphatase measurement (procedure)
C0428333|Fluid sample alkaline phosphatase measurement
C1272113|Plasma alkaline phosphatase level (procedure)
C1272113|Plasma alkaline phosphatase level
