C0519825|COMPREHENSIVE METABOLIC PANEL
C0519825|Comprehensive metabolic panel This panel must include the following: Albumin (82040) Bilirubin, total (82247) Calcium, total (82310) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Phosphatase, alkaline (84075) Potassium (84132) Protein, total (84155) Sodium (84295) Transferase, alanine amino (ALT) (SGPT) (84460) Transferase, aspartate amino (AST) (SGOT) (84450) Urea nitrogen (BUN) (84520)
C0519825|comprehensive metabolic chemical panel
C0519825|Blood test, comprehensive group of blood chemicals
C0519825|comprehensive metabolic panel (lab test)
C0519825|comprehensive metabolic chem panel
C0519825|COMPREHEN METABOLIC PANEL
C2041458|blood chemistry test panels (lab test)
C2041458|blood chemistry test panels
C0438930|Chem. metabolic function tests
C0438930|Chem. metabolic function tests (procedure)
C0201838|Albumin measurement
C0201838|Test;albumin
C0201838|Measurement of albumin
C0201838|Albumin
C0201838|ALB
C0201838|Microalbumin
C0201838|Albumin measurement (procedure)
C0201838|albumin test
C0201925|Calcium; total
C0201925|Calcium Measurement
C0201925|Ca
C0201925|CALCIUM TOTAL
C0201925|Measurement of calcium
C0201925|Calcium level
C0201925|lab-based chem measurements calcium
C0201925|measurement of calcium (lab test)
C0201925|Calcium
C0201925|Ca++
C0201925|Calcium measurement (procedure)
C0201925|Calcium measurement, NOS
C0201925|ASSAY OF CALCIUM
C0201925|Calcium total each test
C0201925|Ca tot ea.tst
C0337438|Glucose
C0337438|Glucose measurement
C0337438|Test;glucose
C0337438|Measurement of glucose
C0337438|GLUC
C0337438|Glucose measurement (procedure)
C0337438|Glucose measurement, NOS
C0337438|glucose test
C0201850|Alkaline phosphatase measurement
C0201850|Phosphatase, alkaline
C0201850|ALP
C0201850|Test;alkaline phosphatase
C0201850|Measurement of alkaline phosphatase
C0201850|ASSAY OF PHOSPHATASE ALKALINE
C0201850|Alkaline Phosphatase
C0201850|ALK phosph
C0201850|Alk phos
C0201850|Alkaline phosphatase measurement (procedure)
C0201850|ASSAY ALKALINE PHOSPHATASE
C0201850|alkaline phosphatase test
C0201952|Chloride Measurement
C0201952|Measurement of chloride
C0201952|Chloride
C0201952|CL
C0201952|Cl-
C0201952|Chloride measurement (procedure)
C0201952|Chloride measurement, NOS
C0201952|Chloride each test
C0201952|chloride ea.tst
C0201975|Creatinine measurement
C0201975|Creatinine; blood
C0201975|Blood creatinine
C0201975|Creatinine
C0201975|Test;creatinine
C0201975|CREATININE BLOOD
C0201975|Blood creatinine level
C0201975|Measurement of creatinine
C0201975|Cr
C0201975|lab-based chem measurements creatinine
C0201975|measurement of creatinine (lab test)
C0201975|CREAT
C0201975|blood creatinine level (lab test)
C0201975|Creatinine measurement (procedure)
C0201975|Creatinine measurement, NOS
C0201975|ASSAY OF CREATININE
C0201975|creatinine test
C0201930|Carbon dioxide content measurement
C0201930|Carbon dioxide
C0201930|CO2 content measurement
C0201930|PCO2, blood
C0201930|CO<sub>2</sub> content measurement
C0201930|PCO<sub>2</sub>, blood
C0201930|Carbon Dioxide Measurement
C0201930|Carbon dioxide (bicarbonate)
C0201930|ASSAY BLOOD CARBON DIOXIDE
C0201930|CARBON DIOXIDE BICARBONATE
C0201930|Measurement of carbon dioxide
C0201930|CO2
C0201930|PCO>2<, blood
C0201930|CO>2< content measurement
C0201930|Carbon dioxide content measurement (procedure)
C0201930|Carbon dioxide measurement (procedure)
C0005845|Blood Urea Nitrogen
C0005845|BUN
C0005845|Nitrogen, Blood Urea
C0005845|Urea Nitrogen, Blood
C0005845|Blood urea nitrogen measurement
C0005845|Urea nitrogen; quantitative
C0005845|Blood urea
C0005845|BUN level
C0005845|Measurement of blood urea nitrogen (BUN)
C0005845|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|Measurement of urea nitrogen (BUN)
C0005845|Urea - blood
C0005845|Blood urea (procedure)
C0005845|blood urea nitrogen measurement (lab test)
C0005845|BUN measurement
C0005845|Blood urea measurement (procedure)
C0005845|Blood urea measurement
C0005845|Blood urea nitrogen measurement (procedure)
C0005845|ASSAY OF UREA NITROGEN
C0200379|GENERAL HEALTH PANEL
C0200379|General health panel (procedure)
C0200379|General health panel This panel must include the following: Comprehensive metabolic panel (80053) Blood count, complete (CBC), automated and automated differential WBC count (85025 or 85027 and 85004) OR Blood count, complete (CBC), automated (85027) and appropriate manual differential WBC count (85007 or 85009) Thyroid stimulating hormone (TSH) (84443)
C0200379|General health panel, NOS
C0201836|Alanine aminotransferase measurement
C0201836|Alanine aminotransferase
C0201836|ALT
C0201836|Transferase; alanine amino (ALT) (SGPT)
C0201836|Test;alanine aminotransferase
C0201836|TRANSFERASE ALANINE AMINO ALT SGPT
C0201836|Measurement of alanine amino transferase (ALT) (SGPT)
C0201836|Measurement of alanine amino transferase
C0201836|Liver enzyme (SGPT), level
C0201836|Alanine amino (alt) (sgpt)
C0201836|SGPT
C0201836|Glutamic-pyruvate transaminase
C0201836|GPT
C0201836|GPT measurement
C0201836|Glutamic pyruvate transaminase measurement
C0201836|SGPT measurement
C0201836|ALT measurement
C0201836|Alanine aminotransferase measurement (procedure)
C0201836|alanine aminotransferase test
C0201913|Bilirubin; total
C0201913|Total Bilirubin Measurement
C0201913|BILIRUBIN TOTAL
C0201913|Measurement of total bilirubin
C0201913|Total bilirubin
C0201913|Total bilirubin (& level) (procedure)
C0201913|Bilirubin, total measurement
C0201913|Bilirubin, total measurement (procedure)
C0201913|Total bilirubin (& level)
C0201913|Bilirubin
C0201913|BILI
C0201913|Total bilirubin level
C0201913|Bilirubin, total measurement (procedure) [Ambiguous]
C0523465|Serum albumin
C0523465|Serum Albumin Measurement
C0523465|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|Albumin; serum, plasma or whole blood
C0523465|serum albumin measurement (lab test)
C0523465|Measurement of albumin in serum
C0523465|Serum albumin (& level) (procedure)
C0523465|Albumin - serum
C0523465|Serum albumin (& level)
C0523465|Serum Albumin Test
C0523465|Albumin measurement, serum
C0523465|Serum albumin level
C0523465|SA - Serum albumin
C0523465|Albumin measurement, serum (procedure)
C0523465|ASSAY OF SERUM ALBUMIN
C0523658|ASSAY GLUCOSE BLOOD QUANT
C0523658|Glucose; quantitative, blood (except reagent strip)
C0523658|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP
C0523658|Glucose measurement, quantitative
C0523658|Glucose measurement, quantitative (procedure)
C0201899|serum SGOT
C0201899|serum AST
C0201899|Aspartate aminotransferase
C0201899|GOT
C0201899|AST
C0201899|Aspartate Aminotransferase Measurement
C0201899|Transferase; aspartate amino (AST) (SGOT)
C0201899|TRANSFERASE ASPARTATE AMINO AST SGOT
C0201899|Liver enzyme (SGOT), level
C0201899|Measurement of aspartate amino transferase
C0201899|Measurement of aspartate amino transferase (AST) (SGOT)
C0201899|AST - aspartate transam SGOT (& level) (procedure)
C0201899|AST - aspartate transam SGOT (& level)
C0201899|Transferase (ast) (sgot)
C0201899|SGOT
C0201899|ASPT
C0201899|Aspartate transferase
C0201899|Asp transferase
C0201899|Serum glutamic-oxaloacetic transferase
C0201899|Glutamic-oxaloacetic transferase
C0201899|Serum Aspartate Transaminase Test
C0201899|AST measurement
C0201899|Glutamic oxaloacetic transaminase measurement
C0201899|GOT measurement
C0201899|SGOT measurement
C0201899|Aspartate aminotransferase measurement (procedure)
C0391938|Chloride; blood
C0391938|Blood chloride
C0391938|Blood chloride level
C0391938|Measurement of chloride in blood
C0391938|Blood chloride level (procedure)
C0391938|blood chloride level (lab test)
C0391938|Chloride measurement, blood
C0391938|Chloride measurement, blood (procedure)
C0391938|ASSAY OF BLOOD CHLORIDE
C0391938|Blood chloride level measurement
C0391938|CHLORIDE BLD
C0523891|serum sodium
C0523891|serum Na+
C0523891|Serum Sodium Measurement
C0523891|serum sodium measurement (lab test)
C0523891|Sodium; serum, plasma or whole blood
C0523891|SODIUM SERUM PLASMA OR WHOLE BLOOD
C0523891|Measurement of sodium in serum
C0523891|Serum sodium (& level) (procedure)
C0523891|Serum sodium (& level)
C0523891|Sodium - serum
C0523891|Serum Sodium Ion Test
C0523891|Sodium measurement, serum
C0523891|Serum sodium level
C0523891|Sodium measurement, serum (procedure)
C0523891|ASSAY OF SERUM SODIUM
C0523891|Serum sodium each test
C0523891|serum sodium ea.tst
C0302353|serum K+
C0302353|Serum Potassium
C0302353|Serum Potassium Measurement
C0302353|serum potassium measurement (lab test)
C0302353|potassium level
C0302353|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|Potassium; serum, plasma or whole blood
C0302353|Measurement of potassium in serum
C0302353|Potassium - serum
C0302353|Serum potassium (& level) (procedure)
C0302353|Serum potassium (& level)
C0302353|Serum potassium level
C0302353|Serum potassium measurement (procedure)
C0302353|ASSAY OF SERUM POTASSIUM
C0373708|Protein, total, except by refractometry; serum, plasma or whole blood
C0373708|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C0373708|ASSAY OF PROTEIN SERUM
C4048459|OBSTETRIC PANEL
C4048459|Obstetric panel This panel must include the following: Blood count, complete (CBC), automated and automated differential WBC count (85025 or 85027 and 85004) OR Blood count, complete (CBC), automated (85027) and appropriate manual differential WBC count (85007 or 85009) Hepatitis B surface antigen (HBsAg) (87340) Antibody, rubella (86762) Syphilis test, non-treponemal antibody; qualitative (eg, VDRL, RPR, ART) (86592) Antibody screen, RBC, each serum technique (86850) Blood typing, ABO (86900) AND Blood typing, Rh (D) (86901)
C0812553|ACUTE HEPATITIS PANEL
C0812553|Acute hepatitis panel This panel must include the following: Hepatitis A antibody (HAAb), IgM antibody (86709) Hepatitis B core antibody (HBcAb), IgM antibody (86705) Hepatitis B surface antigen (HBsAg) (87340) Hepatitis C antibody (86803)
C0519824|ELECTROLYTE PANEL
C0519824|Electrolytes panel
C0519824|Electrolyte panel This panel must include the following: Carbon dioxide (bicarbonate) (82374) Chloride (82435) Potassium (84132) Sodium (84295)
C0519824|blood electrolyte panel
C0519824|blood electrolyte panel (lab test)
C1964052|BASIC METABOLIC PANEL CALCIUM IONIZED
C1964052|METABOLIC PANEL IONIZED CA
C1964052|BMP with ionized calcium
C1964052|basic metabolic panel with ionized calcium (lab test)
C1964052|basic metabolic panel with ionized calcium
C1964052|Basic metabolic panel (Calcium, ionized) This panel must include the following: Calcium, ionized (82330) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Potassium (84132) Sodium (84295) Urea Nitrogen (BUN) (84520)
C0200382|LIPID PANEL
C0200382|lipids test panel
C0200382|lipid panel (lab test)
C0200382|Lipid panel This panel must include the following: Cholesterol, serum, total (82465) Lipoprotein, direct measurement, high density cholesterol (HDL cholesterol) (83718) Triglycerides (84478)
C0200382|Blood test, lipids (cholesterol and triglycerides)
C0200382|Lipid panel (procedure)
C0519823|METABOLIC PANEL TOTAL CA
C0519823|BASIC METABOLIC PANEL CALCIUM TOTAL
C0519823|Basic metabolic panel (Calcium, total) This panel must include the following: Calcium, total (82310) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Potassium (84132) Sodium (84295) Urea nitrogen (BUN) (84520)
C0374833|Organ or Disease Oriented Panels
C0812554|HEPATIC FUNCTION PANEL
C0812554|Hepatic function panel This panel must include the following: Albumin (82040) Bilirubin, total (82247) Bilirubin, direct (82248) Phosphatase, alkaline (84075) Protein, total (84155) Transferase, alanine amino (ALT) (SGPT) (84460) Transferase, aspartate amino (AST) (SGOT) (84450)
C0812554|Hepatic function panel This panel must include the following: Albumin (82040) Bilirubin, total (82247) Bilirubin, direct (82248) Phosphatase, alkaline (84075) Protein, total (84155) Transferase, alanine amino (ALT) (SGPT) (84460) Transferase, aspartate amino (AST) (SGOT)
C0812554|Liver function blood test panel
C0812552|renal function panel (lab test)
C0812552|renal function panel
C0812552|Renal function panel This panel must include the following: Albumin (82040) Calcium, total (82310) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Phosphorus inorganic (phosphate) (84100) Potassium (84132) Sodium (84295) Urea nitrogen (BUN) (84520)
C0812552|Kidney function blood test panel
C0430174|Metabolic function tested
C0430174|Metabolic function test NOS (procedure)
C0430174|Metabolic function test NOS
C0430174|Metabolic function tested (finding)
C0430174|Metabolic function test
C0430174|Metabolic function test (procedure)
C0430174|Metabolic function tested (procedure)
C4050228|OBSTETRIC PANEL
C4050228|Obstetric panel (includes HIV testing) This panel must include the following: Blood count, complete (CBC), and automated differential WBC count (85025 or 85027 and 85004) OR Blood count, complete (CBC), automated (85027) and appropriate manual differential WBC count (85007 or 85009) Hepatitis B surface antigen (HBsAg) (87340) HIV-1 antigen(s), with HIV-1 and HIV-2 antibodies, single result (87389) Antibody, rubella (86762) Syphilis test, non-treponemal antibody; qualitative (eg, VDRL, RPR, ART) (86592) Antibody screen, RBC, each serum technique (86850) Blood typing, ABO (86900) AND Blood typing, Rh (D) (86901)
C0519825|COMPREHENSIVE METABOLIC PANEL
C0519825|Comprehensive metabolic panel This panel must include the following: Albumin (82040) Bilirubin, total (82247) Calcium, total (82310) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Phosphatase, alkaline (84075) Potassium (84132) Protein, total (84155) Sodium (84295) Transferase, alanine amino (ALT) (SGPT) (84460) Transferase, aspartate amino (AST) (SGOT) (84450) Urea nitrogen (BUN) (84520)
C0519825|comprehensive metabolic chemical panel
C0519825|Blood test, comprehensive group of blood chemicals
C0519825|comprehensive metabolic panel (lab test)
C0519825|comprehensive metabolic chem panel
C0519825|COMPREHEN METABOLIC PANEL
C0519824|ELECTROLYTE PANEL
C0519824|Electrolytes panel
C0519824|Electrolyte panel This panel must include the following: Carbon dioxide (bicarbonate) (82374) Chloride (82435) Potassium (84132) Sodium (84295)
C0519824|blood electrolyte panel
C0519824|blood electrolyte panel (lab test)
C0812552|renal function panel (lab test)
C0812552|renal function panel
C0812552|Renal function panel This panel must include the following: Albumin (82040) Calcium, total (82310) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Phosphorus inorganic (phosphate) (84100) Potassium (84132) Sodium (84295) Urea nitrogen (BUN) (84520)
C0812552|Kidney function blood test panel
C2010717|general health test panel (lab test)
C2010717|general health test panel
C0023901|Function Test, Liver
C0023901|Function Tests, Liver
C0023901|Liver Function Test
C0023901|Liver Function Tests
C0023901|Test, Liver Function
C0023901|Tests, Liver Function
C0023901|hepatic function panel
C0023901|hepatic function panel (lab test)
C0023901|Liver function analyses
C0023901|LFTs
C0023901|LFT
C0023901|Liver Study
C0023901|Test;liver function
C0023901|Liver function tests NOS
C0023901|Liver function tests (& [general])
C0023901|Liver funct. test -gen.
C0023901|Liver function tests (& general)
C0023901|Liver function tests (& [general]) (procedure)
C0023901|Liver function tests (procedure)
C0023901|Liver function tests (& general) (procedure)
C0023901|Liver function tests NOS (procedure)
C0023901|Liver function tests - general
C0023901|LFT - Liver function test
C0023901|Hepatic function panel (procedure)
C0023901|Liver function tests - general (procedure)
C0023901|LFT's
C2030682|hepatitis screen panel (lab test)
C2030682|hepatitis screen panel
C0200382|LIPID PANEL
C0200382|lipids test panel
C0200382|lipid panel (lab test)
C0200382|Lipid panel This panel must include the following: Cholesterol, serum, total (82465) Lipoprotein, direct measurement, high density cholesterol (HDL cholesterol) (83718) Triglycerides (84478)
C0200382|Blood test, lipids (cholesterol and triglycerides)
C0200382|Lipid panel (procedure)
C2041460|arthritis test panel
C2041460|arthritis test panel (lab test)
C2041461|torch antibody panel (lab test)
C2041461|torch antibody panel
C0027617|Neonatal Screening
C0027617|Neonatal Screenings
C0027617|Newborn Infant Screenings
C0027617|Screening, Neonatal
C0027617|Screening, Newborn Infant
C0027617|Screenings, Neonatal
C0027617|Screenings, Newborn Infant
C0027617|newborn screen (lab test)
C0027617|newborn screen
C0027617|Newborn Assessment
C0027617|Newborn Screening
C0027617|Screening, Newborn
C0027617|Infant, Newborn, Screening
C0027617|Newborn Infant Screening
C0027617|Neonatal screening (procedure)
C0027617|Neonatal screening, NOS
C0027617|Neonatal screening test
C2210821|basic thyroid panel
C2210821|basic thyroid panel (lab test)
C2106943|comprehensive thyroid panel (lab test)
C2106943|comprehensive thyroid panel
C2237045|Chem 7
C2237045|SMAC 7
C2237045|basic metabolic panel
C2237045|basic metabolic panel (lab test)
C2237045|BMP (basic metabolic panel)
C2237045|Blood test, basic group of blood chemicals
C1315055|Cardiac studies order set
C1315055|cardiac panel (lab test)
C1315055|cardiac panel
C1315055|PANEL.CARDIAC
C3836618|obstetric 1996 panel in serum and blood (lab test)
C3836618|obstetric 1996 panel in serum and blood
C4064645|maternal serum or plasma screening
C4064645|maternal serum or plasma screening (lab test)
C2122148|basic metabolic chem panel
C2122148|basic metabolic chemistry panel
C2122148|basic metabolic chem panel (lab test)
C0438930|Chem. metabolic function tests
C0438930|Chem. metabolic function tests (procedure)
C0523464|Albumin renal clearance measurement
C0523464|Albumin renal clearance measurement (procedure)
C0201837|Albumin/Globulin ratio
C0201837|Albumin globulin ratio
C0201837|A/G ratio
C0201837|Albumin/Globulin ratio (procedure)
C0523465|Serum albumin
C0523465|Serum Albumin Measurement
C0523465|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|Albumin; serum, plasma or whole blood
C0523465|serum albumin measurement (lab test)
C0523465|Measurement of albumin in serum
C0523465|Serum albumin (& level) (procedure)
C0523465|Albumin - serum
C0523465|Serum albumin (& level)
C0523465|Serum Albumin Test
C0523465|Albumin measurement, serum
C0523465|Serum albumin level
C0523465|SA - Serum albumin
C0523465|Albumin measurement, serum (procedure)
C0523465|ASSAY OF SERUM ALBUMIN
C0201838|Albumin measurement
C0201838|Test;albumin
C0201838|Measurement of albumin
C0201838|Albumin
C0201838|ALB
C0201838|Microalbumin
C0201838|Albumin measurement (procedure)
C0201838|albumin test
C1278236|24 hour urine albumin output
C1278236|24 hour urine albumin output (procedure)
C1278236|24 hour urine albumin output measurement (procedure)
C1278236|24 hour urine albumin output measurement
C0523466|Albumin; urine or other source, quantitative, each specimen
C0523466|ALBUMIN URINE/OTHER SOURCE QUAN EACH SPECIMEN
C0523466|Albumin measurement, urine, quantitative
C0523466|Albumin measurement, urine, quantitative (procedure)
C0523466|ASSAY OF URINE ALBUMIN
C0373533|Albumin; urine, microalbumin, semiquantitative (eg, reagent strip assay)
C0373533|MICROALBUMIN SEMIQUANT
C0373533|ALBUMIN URINE MICROALBUMIN SEMIQUANTITATIVE
C0373533|Semiquantitative analysis of microalbumin in urine
C1504155|serum albumin ischemia modified (lab test)
C1504155|serum albumin ischemia modified
C1504155|ischemia-modified serum albumin
C1504155|ALBUMIN ISCHEMIA MODIFIED
C1504155|serum albumin ischemia modified lab procedure
C1504155|Albumin; ischemia modified
C0373532|Albumin; urine, microalbumin, quantitative
C0373532|MICROALBUMIN QUANTITATIVE
C0373532|ALBUMIN URINE MICROALBUMIN QUANTIATIVE
C0523674|ALBGLYCA
C0523674|Glycated Albumin
C0523674|Glycated Albumin Measurement
C0523674|Glycated albumin measurement (procedure)
C1278275|Cerebrospinal fluid albumin level
C1278275|Cerebrospinal fluid albumin level (procedure)
C1278275|Cerebrospinal fluid albumin measurement (procedure)
C1278275|Cerebrospinal fluid albumin measurement
C0428520|Fluid sample albumin level
C0428520|Fluid sample albumin measurement (procedure)
C0428520|Fluid sample albumin measurement
C0428623|Albumin/immunoglobulin G ratio
C0428623|IgG - Albumin/immunoglobulin G ratio
C0428623|Albumin/immunoglobulin G ratio measurement (procedure)
C0428623|Albumin/immunoglobulin G ratio measurement
C1272106|Plasma albumin level (procedure)
C1272106|Plasma albumin level
C1273508|Serum prealbumin level
C1273508|Serum prealbumin level (procedure)
C1318429|Measurement of albumin in urine
C1318429|Urine albumin (& level) (procedure)
C1318429|Urine albumin (& level)
C1318429|Urine albumin level
C1318429|Urine albumin measurement (procedure)
C1318429|Urine albumin measurement
C0523463|CSF albumin/plasma albumin ratio measurement (procedure)
C0523463|Cerebrospinal fluid albumin/plasma albumin ratio measurement (procedure)
C0523463|Cerebrospinal fluid albumin/plasma albumin ratio measurement
C0523463|CSF albumin/plasma albumin ratio measurement
C0025634|Methemalbumin
C0025634|Methemalbumin Assay
C0025634|Methemalbumin (protein) level
C0025634|Measurement of methemalbumin
C0025634|Methemalbumin measurement
C0025634|Methaemalbumin measurement
C0025634|Methemalbumin measurement (procedure)
C0025634|ASSAY OF METHEMALBUMIN
C1293929|Measurement of ratio of analyte to albumin (procedure)
C1293929|Measurement of ratio of analyte to albumin
C0201925|Calcium; total
C0201925|Calcium Measurement
C0201925|Ca
C0201925|CALCIUM TOTAL
C0201925|Measurement of calcium
C0201925|Calcium level
C0201925|lab-based chem measurements calcium
C0201925|measurement of calcium (lab test)
C0201925|Calcium
C0201925|Ca++
C0201925|Calcium measurement (procedure)
C0201925|Calcium measurement, NOS
C0201925|ASSAY OF CALCIUM
C0201925|Calcium total each test
C0201925|Ca tot ea.tst
C0728876|serum calcium
C0728876|serum Ca++
C0728876|Serum Calcium Measurement
C0728876|Serum calcium (& level) (procedure)
C0728876|Serum calcium (& level)
C0728876|Calcium - serum
C0728876|Serum Calcium Test
C0728876|Serum calcium level
C0728876|Serum calcium measurement (procedure)
C0428303|Urine calcium
C0428303|Urine Calcium Measurement
C0428303|urine calcium measurement (lab test)
C0428303|Urine calcium level
C0428303|Calcium - urine
C0428303|Urine calcium (& level) (procedure)
C0428303|Urine calcium (& level)
C0428303|Urine Calcium Test
C0428303|Calcium measurement, urine
C0428303|Calcium measurement, urine (procedure)
C0430040|Calcium profile
C0430040|Calcium profile (procedure)
C1278284|Calculus calcium content
C1278284|Calculus calcium content (finding)
C1278284|Calculus calcium content measurement (procedure)
C1278284|Calculus calcium content measurement
C1271835|Fluid sample calcium level (procedure)
C1271835|Fluid sample calcium level
C2711247|Calculation of ionized calcium concentration
C2711247|Calculation of ionised calcium concentration
C2711247|Calculation of ionized calcium concentration (procedure)
C2732404|Corrected measurement of calcium
C2732404|Corrected measurement of calcium (procedure)
C2732404|Calcium Corrected
C2732404|CACR
C2732404|Calcium Corrected Measurement
C3272884|Calcium Clearance Measurement
C3272884|Calcium Clearance
C3272884|CACLR
C0201927|Measurement of serum ionized calcium
C0201927|Measurement of serum ionised calcium
C0201927|Serum ionized calcium measurement
C0201927|Serum ionised calcium measurement (procedure)
C0201927|Measurement of serum ionized calcium (procedure)
C0201927|serum ionized calcium measurement (lab test)
C0201927|ionized calcium level
C0201927|Ionized Calcium Measurement
C0201927|Measurement of ionized calcium
C0201927|Serum ionised calcium level (procedure)
C0201927|Serum ionised calcium level
C0201927|Calcium, serum, ionized measurement
C0201927|Calcium, serum, ionized measurement (procedure)
C0201927|Calcium, serum, ionised measurement
C0201927|CAION
C0201927|Calcium, Ionized
C0201927|Serum ionized calcium level
C0201927|Serum ionised calcium measurement
C0373563|Calcium; urine quantitative, timed specimen
C0373563|CALCIUM URINE QUANTITATIVE TIMED SPECIMEN
C0373563|ASSAY OF CALCIUM IN URINE
C0523539|Calcium; after calcium infusion test
C0523539|Calcium challenge tests (procedure)
C0523539|CALCIUM AFTER CALCIUM INFUSION TEST
C0523539|Measurement of calcium after calcium infusion test
C0523539|Calcium challenge tests
C0523539|Calcium measurement after calcium infusion
C0523539|Calcium infusion test
C0489943|Calcium; ionized
C0489943|Ionized Calcium Assay
C0489943|Calcium ionized
C0489943|Ionized calcium
C0489943|Calcium ionised
C0489943|ASSAY OF CALCIUM
C0489943|Calcium ionized each test
C0489943|Ca ionized ea.tst
C3830083|FECA
C3830083|Fractional Excretion of Calcium
C3830083|Fractional Excretion of Ca
C3830083|Fractional Calcium Excretion
C0201928|Calcium excretion, 2-hour collection, fasting, urine
C0201928|Calcium excretion, 2-hour collection, fasting, urine (procedure)
C0278369|Calcium measurement in 24 hour excretion in feces
C0278369|Calcium measurement in 24 hour excretion in faeces
C0278369|Calcium measurement in 24 hour excretion in feces (procedure)
C0278369|Calcium measurement, 24H stool
C0278369|Calcium total measurement, 24 hour excretion in stool
C0729820|Blood calcium
C0729820|Blood calcium level
C0729820|Blood calcium level (procedure)
C0729820|blood calcium measurement (lab test)
C0729820|calcium blood
C0729820|blood calcium measurement
C0729820|Blood calcium measurement (procedure)
C0428613|Calcium to Creatinine Ratio Measurement
C0428613|Calcium/creatinine ratio
C0428613|Calcium/creatinine ratio (procedure)
C0428613|CACREAT
C0428613|Calcium/Creatinine
C0428613|Calcium/creatinine ratio measurement (procedure)
C0428613|Calcium/creatinine ratio measurement
C0523660|Glucose measurement, post glucose dose
C0523660|Glucose measurement, post glucose dose (procedure)
C0337438|Glucose
C0337438|Glucose measurement
C0337438|Test;glucose
C0337438|Measurement of glucose
C0337438|GLUC
C0337438|Glucose measurement (procedure)
C0337438|Glucose measurement, NOS
C0337438|glucose test
C0392201|Blood glucose
C0392201|blood glucose tests (lab test)
C0392201|blood glucose tests
C0392201|Blood glucose measurement
C0392201|blood glucose level
C0392201|blood glucose measurement (lab test)
C0392201|Blood glucose (sugar) level
C0392201|Measurement of glucose in blood
C0392201|Blood Sugar
C0392201|Glucose Measurement, Blood
C0392201|Blood sugar level
C0392201|BS - Blood glucose level
C0392201|Glucose measurement, blood (procedure)
C0202048|Glucose measurement by monitoring device
C0202048|Glucose measurement by monitoring device (procedure)
C0202048|Glucose measurement by monitoring device (procedure) [Ambiguous]
C2732668|Urea, electrolytes and glucose measurement
C2732668|Measurement of urea, sodium, potassium, chloride, bicarbonate and glucose (procedure)
C2732668|Measurement of urea, sodium, potassium, chloride, bicarbonate and glucose
C2732640|Calculation of estimated average glucose based on hemoglobin A1c (procedure)
C2732640|Calculation of estimated average glucose based on hemoglobin A1c
C2732640|Estimated average glucose measurement
C2732640|Calculation of estimated average glucose based on haemoglobin A1c
C0204885|Ward glucometer test
C0204885|Ward glucometer test (procedure)
C0202040|cerebrospinal fluid glucose (lab test)
C0202040|cerebrospinal fluid glucose
C0202040|CSF glucose
C0202040|Glucose CSF
C0202040|Glucose measurement, cerebrospinal fluid
C0202040|Glucose measurement, cerebrospinal fluid (procedure)
C0202040|Glucose measurement, CSF (procedure)
C0202040|CSF Glucose Test
C0202040|Glucose measurement, CSF
C1271625|Urine clinitest
C1271625|Urine clinitest (procedure)
C0202041|serum glucose
C0202041|Serum Glucose Measurement
C0202041|Serum Glucose Test
C0202041|Glucose measurement, serum
C0202041|Glucose measurement, serum (procedure)
C0202042|Plasma Glucose Measurement
C0202042|plasma glucose measurement (lab test)
C0202042|plasma glucose
C0202042|Plasma glucose level
C0202042|Plasma glucose level (procedure)
C0202042|Glucose measurement, plasma
C0202042|Glucose measurement, plasma (procedure)
C0523655|Glucose cerebrospinal fluid/glucose plasma ratio measurement (procedure)
C0523655|Glucose cerebrospinal fluid/glucose plasma ratio measurement
C0523655|Glucose CSF/glucose plasma ratio measurement (procedure)
C0523655|Glucose CSF/glucose plasma ratio measurement
C0004076|urine glucose
C0004076|Glucose measurement, urine
C0004076|urine glucose measurement (lab test)
C0004076|urine glucose measurement
C0004076|Glucose urine
C0004076|Urine screen for sugar (& [glucose]) (procedure)
C0004076|Sugar - urine test (& glucose)
C0004076|Urine glucose test NOS
C0004076|Urine glucose test NOS (procedure)
C0004076|Sugar - urine test (& glucose) (procedure)
C0004076|Urine test for glucose (procedure)
C0004076|Urine screen for sugar (& [glucose])
C0004076|Urine test for glucose
C0004076|Glucose - urine test
C0004076|Sugar - urine test
C0004076|Urine Glucose Test
C0004076|Glucose measurement, urine (procedure)
C0373621|Glucose test; post glucose dose (includes glucose)
C0373621|Glucose; post glucose dose (includes glucose)
C0373621|GLUCOSE POST GLUCOSE DOSE
C0373621|Blood glucose (sugar) level after receiving dose of glucose
C0373621|Measurement of glucose after glucose dose
C0373621|GLUCOSE TEST
C0523658|ASSAY GLUCOSE BLOOD QUANT
C0523658|Glucose; quantitative, blood (except reagent strip)
C0523658|GLUCOSE QUANTITATIVE BLOOD XCPT REAGENT STRIP
C0523658|Glucose measurement, quantitative
C0523658|Glucose measurement, quantitative (procedure)
C0373622|Glucose; tolerance test (GTT), 3 specimens (includes glucose)
C0373622|GLUCOSE TOLERANCE TEST GTT 3 SPECIMENS
C0373622|Glucose tolerance test (gtt)
C0373623|GLUCOSE TOLERANCE EA ADDL BEYOND 3 SPECIMENS
C0373623|Glucose; tolerance test, each additional beyond 3 specimens (List separately in addition to code for primary procedure)
C0373623|Gtt-added samples
C0373620|Glucose; blood, reagent strip
C0373620|blood glucose determination by reagent strip (lab test)
C0373620|blood glucose determination by reagent strip
C0373620|blood glucose level by reagent strip
C0373620|GLUCOSE BLOOD REAGENT STRIP
C0373620|Blood glucose (sugar) measurement using reagent strip
C0373620|Measurement of glucose in blood using reagent strip
C0373620|REAGENT STRIP/BLOOD GLUCOSE
C4064987|glucose in serum or plasma (lab test)
C4064987|glucose in serum or plasma
C0202045|Glucose measurement, fasting
C0202045|Glucose measurement, fasting (procedure)
C0202045|fasting glucose test
C0202045|Test;glucose;fasting
C0202046|Glucose measurement, random
C0202046|Glucose measurement, random (procedure)
C0202046|random glucose test
C0202046|Test;glucose;random
C0017741|Glucose Tolerance Test
C0017741|Glucose Tolerance Tests
C0017741|Test;glucose tolerance
C0017741|Glucose tolerance test (GTT)
C0017741|Blood glucose (sugar) tolerance test
C0017741|Glucose tolerance test NOS
C0017741|Glucose tolerance test NOS (procedure)
C0017741|GTT
C0017741|GTT - Glucose tolerance test
C0017741|OGTT - Oral glucose tolerance test
C0017741|Glucose challenge test
C0017741|Glucose tolerance test (procedure)
C0017741|Glucose tolerance test, NOS
C0523657|Glucose measurement, tolbutamide tolerance test
C0523657|Glucose measurement, tolbutamide tolerance test (procedure)
C1272314|Fecal clinitest (procedure)
C1272314|Faecal clinitest (procedure)
C1272314|Faecal clinitest
C1272314|Fecal clinitest
C0427743|Glucose concentration
C0427743|Glucose concentration, test strip measurement (procedure)
C0427743|Glucose concentration, test strip measurement
C1295145|Glucose measurement estimated from glycated haemoglobin
C1295145|Glucose measurement estimated from glycated hemoglobin (procedure)
C1295145|Glucose measurement estimated from glycated hemoglobin
C0428549|Fluid sample glucose measurement
C0428549|body fluid glucose measurement (lab test)
C0428549|body fluid glucose
C0428549|body fluid glucose measurement
C0428549|Measurement of glucose in body fluid
C0428549|Body Fluid Glucose Test
C0428549|Fluid sample glucose level
C0428549|Fluid sample glucose measurement (procedure)
C0428549|Glucose measurement, body fluid
C1319276|Faecal glucose level
C1319276|Faecal glucose measurement
C1319276|Fecal glucose level (procedure)
C1319276|Fecal glucose level
C1319276|Fecal glucose measurement
C0201850|Alkaline phosphatase measurement
C0201850|Phosphatase, alkaline
C0201850|ALP
C0201850|Test;alkaline phosphatase
C0201850|Measurement of alkaline phosphatase
C0201850|ASSAY OF PHOSPHATASE ALKALINE
C0201850|Alkaline Phosphatase
C0201850|ALK phosph
C0201850|Alk phos
C0201850|Alkaline phosphatase measurement (procedure)
C0201850|ASSAY ALKALINE PHOSPHATASE
C0201850|alkaline phosphatase test
C0036776|serum alkaline phosphatase
C0036776|SAP
C0036776|Serum Alkaline Phosphatase Measurement
C0036776|serum alkaline phosphatase measurement (lab test)
C0036776|Serum alkaline phosphatase (& level)
C0036776|Serum alkaline phosphatase (& level) (procedure)
C0036776|Alk. phosphatase -serum
C0036776|Alkaline phosphatase (& level (& serum))
C0036776|Phosph.- alk. - serum
C0036776|Serum alkaline phosphatase NOS
C0036776|Alkaline phosphatase (& level (& serum)) (procedure)
C0036776|Serum alkaline phosphatase NOS (procedure)
C0036776|Serum Alkaline Phosphatase Test
C0036776|Serum alkaline phosphatase level
C0036776|Serum alkaline phosphatase measurement (procedure)
C1293930|Measurement of ratio of analyte to alkaline phosphatase (procedure)
C1293930|Measurement of ratio of analyte to alkaline phosphatase
C0201851|Phosphatase, alkaline; isoenzymes
C0201851|Measurement of alkaline phosphatase isoenzymes
C0201851|ASSAY OF PHOSPHATASE ALKALINE ISOENZYMES
C0201851|Alkaline phosphatase isoenzymes measurement
C0201851|Alkaline phosphatase isoenzymes measurement (procedure)
C0201851|ASSAY ALKALINE PHOSPHATASES
C0201855|Alkaline phosphatase, heat stable measurement
C0201855|Phosphatase, alkaline; heat stable (total not included)
C0201855|Measurement of heat stable alkaline phosphatase
C0201855|ASSAY OF PHOSPHATASE ALKALINE HEAT STABLE
C0201855|Thermostable alkaline phosphatase measurement
C0201855|Alkaline phosphatase, heat stable measurement (procedure)
C0201855|ASSAY ALKALINE PHOSPHATASE
C2984961|Bone Specific Alkaline Phosphatase Measurement
C2984961|Bone Alkaline Phosphatase Measurement
C2984961|Bone Specific Alkaline Phosphatase
C2984961|ALPBS
C2984961|Bone ALP Measurement
C3898585|Liver Specific Alkaline Phosphatase Measurement
C3898585|ALPLS
C3898585|Liver Specific Alkaline Phosphatase
C3898710|Intestinal Specific Alkaline Phosphatase
C3898710|ALPIS
C3898710|Intestinal Specific Alkaline Phosphatase Measurement
C0200697|Leukocyte alkaline phosphatase level
C0200697|Leucocyte alkaline phosphatase level
C0200697|Leucocyte alkaline phosphatase level (procedure)
C0200697|Leukocyte alkaline phosphatase score
C0200697|Leucocyte alkaline phosphatase score
C0200697|Leukocyte alkaline phosphatase score (procedure)
C0200697|Leukocyte alkaline phosphatase score (observable entity)
C0200697|Neutrophil alkaline phosphatase score
C0200697|LAP score
C0200697|LAP - Neutrophil alkaline phosphatase score
C0200697|LAP - Neutrophil alkaline phosphatase score measurement
C0201852|Placental alkaline phosphatase measurement
C0201852|PLAP measurement
C0201852|Placental alkaline phosphatase measurement (procedure)
C0201853|Intestinal alkaline phosphatase measurement
C0201853|IAP measurement
C0201853|Intestinal alkaline phosphatase measurement (procedure)
C0201854|Germ cell alkaline phosphatase measurement
C0201854|GCAP measurement
C0201854|Germ cell alkaline phosphatase measurement (procedure)
C0428333|Fluid sample alkaline phosphatase level
C0428333|Fluid sample alkaline phosphatase measurement (procedure)
C0428333|Fluid sample alkaline phosphatase measurement
C1272113|Plasma alkaline phosphatase level (procedure)
C1272113|Plasma alkaline phosphatase level
C0391938|Chloride; blood
C0391938|Blood chloride
C0391938|Blood chloride level
C0391938|Measurement of chloride in blood
C0391938|Blood chloride level (procedure)
C0391938|blood chloride level (lab test)
C0391938|Chloride measurement, blood
C0391938|Chloride measurement, blood (procedure)
C0391938|ASSAY OF BLOOD CHLORIDE
C0391938|Blood chloride level measurement
C0391938|CHLORIDE BLD
C1317978|Serum Chloride Measurement
C1317978|serum chloride measurement (lab test)
C1317978|chloride level
C1317978|Serum chloride (& level)
C1317978|Serum chloride (& level) (procedure)
C1317978|Serum chloride level
C1317978|Serum chloride measurement (procedure)
C2711521|Measurement of chloride in stool specimen (procedure)
C2711521|Measurement of chloride in stool specimen
C2732591|Urea, electrolytes and creatinine measurement
C2732591|Measurement of urea, sodium, potassium, chloride, bicarbonate and creatinine
C2732591|Measurement of urea, sodium, potassium, chloride, bicarbonate and creatinine (procedure)
C2732591|lab-based chem measure urea, na, potassium chloride, bicarbonate, creatinine
C2732591|measurement of urea, sodium, potassium chloride, bicarbonate, and creatinine
C2732591|measurement of urea, sodium, potassium chloride, bicarbonate, and creatinine (lab test)
C0729818|Blood chloride level result
C0428295|sweat test for chloride (lab test)
C0428295|sweat test for chloride
C0428295|Sweat chloride (& level) (procedure)
C0428295|Sweat chloride (& level)
C0428295|Sweat chloride
C0428295|Sweat chloride test
C0428295|Chloride Sweat Test
C0428295|Cystic fibrosis sweat test
C0428295|Chloride measurement, sweat
C0428295|Sweat chloride level
C0428295|Cystic fibrosis sweat test (procedure)
C0201953|Chloride; urine
C0201953|urine chloride measurement (lab test)
C0201953|urine chloride measurement
C0201953|urine chloride
C0201953|Urine chloride level
C0201953|Measurement of chloride in urine
C0201953|Urine chloride level (procedure)
C0201953|Urine Chloride Test
C0201953|Chloride measurement, urine
C0201953|Chloride measurement, urine (procedure)
C0201953|ASSAY OF URINE CHLORIDE
C0201953|CHLORIDE URINE
C0373575|Chloride; other source
C0373575|ASSAY OTHER FLUID CHLORIDES
C0373575|CHLORIDE OTHER SOURCE
C3830082|Fractional Excretion of Chloride
C3830082|Fractional Chloride Excretion
C3830082|FECl
C3830082|Fractional Excretion of Cl
C0201952|Chloride Measurement
C0201952|Measurement of chloride
C0201952|Chloride
C0201952|CL
C0201952|Cl-
C0201952|Chloride measurement (procedure)
C0201952|Chloride measurement, NOS
C0201952|Chloride each test
C0201952|chloride ea.tst
C0428297|CSF chloride measurement (procedure)
C0428297|CSF: chloride level NOS (procedure)
C0428297|Cerebrospinal fluid chloride measurement (procedure)
C0428297|Cerebrospinal fluid chloride measurement
C0428297|CSF Cl
C0428297|CSF chloride
C0428297|CSF chloride level
C0428297|cerebrospinal fluid chloride measurement (lab test)
C0428297|Cerebrospinal fluid: chloride level NOS (procedure)
C0428297|Cerebrospinal fluid: chloride level NOS
C0428297|CSF: chloride level NOS
C0428297|CSF Chloride Test
C0428297|CSF: chloride level
C0428297|CSF chloride measurement
C0428296|Body Fluid Chloride Test
C0428296|Fluid sample chloride
C0428296|Fluid sample chloride level
C0428296|Chloride measurement, body fluid (procedure)
C0428296|Chloride measurement, body fluid
C0428296|Body fluid chloride measurement
C0428296|Chloride measurement, body fluid, NOS
C1276037|Plasma chloride level
C1276037|Plasma chloride measurement (procedure)
C1276037|Plasma chloride measurement
C0430179|Sweat test
C0430179|Sweat test NOS
C0430179|Sweat test (procedure)
C0430179|Sweat test NOS (procedure)
C0430179|sweat tests
C0430179|sweat tests (lab test)
C0430179|Sweat screening test
C0201975|Creatinine measurement
C0201975|Creatinine; blood
C0201975|Blood creatinine
C0201975|Creatinine
C0201975|Test;creatinine
C0201975|CREATININE BLOOD
C0201975|Blood creatinine level
C0201975|Measurement of creatinine
C0201975|Cr
C0201975|lab-based chem measurements creatinine
C0201975|measurement of creatinine (lab test)
C0201975|CREAT
C0201975|blood creatinine level (lab test)
C0201975|Creatinine measurement (procedure)
C0201975|Creatinine measurement, NOS
C0201975|ASSAY OF CREATININE
C0201975|creatinine test
C2981749|Urinary Creatinine Assay
C2981751|Serum Creatinine Assay
C0201976|serum creatinine
C0201976|Serum Creatinine Measurement
C0201976|Creatinine measurement, serum (procedure)
C0201976|serum creatinine level
C0201976|serum creatinine measurement (lab test)
C0201976|Creatinine.serum
C0201976|Serum creatinine (& level) (procedure)
C0201976|Creatinine - serum
C0201976|Serum creatinine NOS (procedure)
C0201976|Serum creatinine NOS
C0201976|Serum creatinine (& level)
C0201976|Serum Creatinine Test
C0201976|Creatinine measurement, serum
C1278055|plasma creatinine measurement
C1278055|Plasma creatinine level
C1278055|Plasma creatinine level (procedure)
C1278055|plasma creatinine
C1278055|Plasma creatinine measurement (lab test)
C1278055|Plasma creatinine measurement (procedure)
C1318439|Urine Creatinine Measurement
C1318439|urine creatinine measurement (lab test)
C1318439|urine creatinine
C1318439|creatinine level
C1318439|Creatinine urine
C1318439|Urine creatinine (& level) (procedure)
C1318439|Urine creatinine (& level)
C1318439|Creatinine - urine
C1318439|Creatinine measurement, urine
C1318439|Urine creatinine measurement (procedure)
C1318439|Urine creatinine level
C0201977|urine creatinine 12-hour
C0201977|12-hour urine creatinine measurement
C0201977|12-hour urine creatinine measurement (lab test)
C0201977|12-hour creatinine level
C0201977|Creatinine measurement, 12 hour urine
C0201977|Creatinine measurement, 12 hour urine (procedure)
C3694999|creatinine concentration (serum or plasma)
C3694999|serum or plasma creatinine concentration (lab test)
C3694999|serum or plasma creatinine concentration
C3694393|lab-based chem measurements creatinine clearance - glomerular filtration (lab test)
C3694393|lab-based chem measurements creatinine clearance - glomerular filtration
C0373594|Creatinine; other source
C0373594|CREATININE OTHER SOURCE
C0373594|ASSAY OF URINE CREATININE
C0373595|Creatinine; clearance
C0373595|Creatinine renal clearance
C0373595|Measurement of renal clearance of creatinine
C0373595|Creatinine clearance test
C0373595|Creatinine clearance test (procedure)
C0373595|Measurement of renal clearance of creatinine (procedure)
C0373595|Creatinine clearance measurement
C0373595|Creatinine renal clearance measurement (procedure)
C0373595|Creatinine clearance-glom filt
C0373595|Creatinine clearance study (procedure)
C0373595|Creatinine renal clearance measurement
C0373595|Creatinine clearance
C0373595|Creatinine clearance study
C0373595|CREATCLR
C0373595|renal function creatinine clearance
C0373595|creatinine renal clearance (procedure)
C0428279|Finding of creatinine level
C0428279|lab-based chem measurements creatinine level finding
C0428279|creatinine level finding (lab test)
C0428279|creatinine level finding
C0428279|Creatinine level
C0428279|Creatinine level - finding
C0428279|Finding of creatinine level (finding)
C0523586|Creatinine challenge tests
C0523586|Creatinine challenge tests (procedure)
C1278053|Corrected plasma creatinine level
C1278053|Corrected plasma creatinine level (procedure)
C1278053|Corrected plasma creatinine measurement (procedure)
C1278053|Corrected plasma creatinine measurement
C1261396|Fluid sample creatinine measurement
C1261396|Body Fluid Creatinine Test
C1261396|Creatinine measurement, body fluid
C1261396|Fluid sample creatinine measurement (procedure)
C1261396|Fluid sample creatinine level
C1293927|Measurement of ratio of analyte to creatinine (procedure)
C1293927|Measurement of ratio of analyte to creatinine
C1446045|5-Hydroxyindoleacetic acid/creatinine ratio measurement (procedure)
C1446045|5-Hydroxyindoleacetic acid/creatinine ratio measurement
C1446045|5HIAA/creatinine ratio
C1446063|Aminolaevulinic acid / creatinine ratio measurement
C1446063|Aminolaevulinic acid/creatinine ratio measurement
C1446063|Aminolevulinic acid / creatinine ratio measurement
C1446063|Aminolevulinic acid/creatinine ratio measurement (procedure)
C1446063|Aminolevulinic acid/creatinine ratio measurement
C1446063|ALA/creatinine ratio
C1446080|Magnesium to Creatinine Ratio Measurement
C1446080|Magnesium/Creatinine
C1446080|MGCREAT
C1446080|Magnesium / creatinine ratio measurement (procedure)
C1446080|Magnesium / creatinine ratio measurement
C1446080|Magnesium/creatinine ratio
C1446178|Retinol binding protein / creatinine ratio measurement (procedure)
C1446178|Retinol binding protein / creatinine ratio measurement
C1531635|Citrate:creatinine ratio (procedure)
C1531635|Citrate:creatinine ratio
C1531635|Measurement of ratio of citrate to creatinine (procedure)
C1531635|Measurement of ratio of citrate to creatinine
C1531635|Meausrement of ratio of citrate to creatinine
C1531635|Meausrement of ratio of citrate to creatinine (procedure)
C1531635|Citrate/Creatinine
C1531635|Citrate to Creatinine Ratio Measurement
C1531635|Citric Acid/Creatinine
C1531635|CITCREAT
C0596252|carbon dioxide fixation
C0596253|carbon dioxide tension
C0596254|carbon dioxide transport
C0201930|Carbon dioxide content measurement
C0201930|Carbon dioxide
C0201930|CO2 content measurement
C0201930|PCO2, blood
C0201930|CO<sub>2</sub> content measurement
C0201930|PCO<sub>2</sub>, blood
C0201930|Carbon Dioxide Measurement
C0201930|Carbon dioxide (bicarbonate)
C0201930|ASSAY BLOOD CARBON DIOXIDE
C0201930|CARBON DIOXIDE BICARBONATE
C0201930|Measurement of carbon dioxide
C0201930|CO2
C0201930|PCO>2<, blood
C0201930|CO>2< content measurement
C0201930|Carbon dioxide content measurement (procedure)
C0201930|Carbon dioxide measurement (procedure)
C2144939|Serum Total CO2
C2144939|Serum Total CO2 (lab test)
C2144939|total CO2 content
C0201931|Partial Pressure of Carbon Dioxide Measurement
C0201931|Carbon dioxide measurement, partial pressure
C0201931|PCO2
C0201931|Partial Pressure Carbon Dioxide
C0201931|PaCO2 measurement
C0201931|Carbon dioxide measurement, partial pressure (procedure)
C0005845|Blood Urea Nitrogen
C0005845|BUN
C0005845|Nitrogen, Blood Urea
C0005845|Urea Nitrogen, Blood
C0005845|Blood urea nitrogen measurement
C0005845|Urea nitrogen; quantitative
C0005845|Blood urea
C0005845|BUN level
C0005845|Measurement of blood urea nitrogen (BUN)
C0005845|ASSAY OF UREA NITROGEN QUANTITATIVE
C0005845|Measurement of urea nitrogen (BUN)
C0005845|Urea - blood
C0005845|Blood urea (procedure)
C0005845|blood urea nitrogen measurement (lab test)
C0005845|BUN measurement
C0005845|Blood urea measurement (procedure)
C0005845|Blood urea measurement
C0005845|Blood urea nitrogen measurement (procedure)
C0005845|ASSAY OF UREA NITROGEN
C0455273|Serum urea level
C0455273|Serum urea level (procedure)
C0455273|Serum urea measurement (procedure)
C0455273|Serum urea measurement
C0729828|Plasma urea level
C0729828|Plasma urea level (procedure)
C0729828|Plasma urea measurement (procedure)
C0729828|Plasma urea measurement
C0201922|BUN/Creatinine ratio (procedure)
C0201922|Blood urea nitrogen (BUN)/Creatinine ratio
C0201922|Blood urea nitrogen/creatinine ratio (procedure)
C0201922|Blood urea nitrogen/creatinine ratio
C0201922|Blood urea nitrogen (BUN)/Creatinine ratio (procedure)
C0201922|BUN/Creatinine ratio
C0201922|bun/creatinine ratio (lab test)
C0201922|Urea nitrogen/creatinine ratio, serum
C2208743|serum BUN/creatinine ratio
C2208743|serum BUN/creatinine ratio (lab test)
C2097174|BUN using reagent strip (lab test)
C2097174|BUN using reagent strip
C2097174|BUN by reagent strip
C2097689|BUN was obtained pre-procedure
C2097689|BUN was obtained pre-procedure (lab test)
C2097689|a BUN level was obtained pre-procedure
C0729816|Blood potassium level
C0729816|Blood potassium level (procedure)
C0729816|Blood potassium measurement (procedure)
C0729816|Blood potassium measurement
C4027477|urea nitrogen level in serum or plasma (lab test)
C4027477|urea nitrogen level in serum or plasma
C0200379|GENERAL HEALTH PANEL
C0200379|General health panel (procedure)
C0200379|General health panel This panel must include the following: Comprehensive metabolic panel (80053) Blood count, complete (CBC), automated and automated differential WBC count (85025 or 85027 and 85004) OR Blood count, complete (CBC), automated (85027) and appropriate manual differential WBC count (85007 or 85009) Thyroid stimulating hormone (TSH) (84443)
C0200379|General health panel, NOS
C0201836|Alanine aminotransferase measurement
C0201836|Alanine aminotransferase
C0201836|ALT
C0201836|Transferase; alanine amino (ALT) (SGPT)
C0201836|Test;alanine aminotransferase
C0201836|TRANSFERASE ALANINE AMINO ALT SGPT
C0201836|Measurement of alanine amino transferase (ALT) (SGPT)
C0201836|Measurement of alanine amino transferase
C0201836|Liver enzyme (SGPT), level
C0201836|Alanine amino (alt) (sgpt)
C0201836|SGPT
C0201836|Glutamic-pyruvate transaminase
C0201836|GPT
C0201836|GPT measurement
C0201836|Glutamic pyruvate transaminase measurement
C0201836|SGPT measurement
C0201836|ALT measurement
C0201836|Alanine aminotransferase measurement (procedure)
C0201836|alanine aminotransferase test
C1883008|Serum Alanine Aminotransferase Measurement
C1883008|Serum SGPT Measurement
C1883008|Serum Alanine Transaminase Measurement
C1883008|serum alanine aminotransferase measurement (lab test)
C1883008|ALT (SGPT) level
C0428324|Alanine transaminase level
C0428324|Alanine transaminase level (procedure)
C0428325|ALT/SGPT serum level
C0428325|ALT/SGPT serum level (procedure)
C0523461|ALT measurement, method with pyridoxal-5'-phosphate (procedure)
C0523461|Alanine aminotransferase (ALT) measurement, method with pyridoxal-5'-phosphate
C0523461|Alanine aminotransferase measurement, method with pyridoxal-5'-phosphate (procedure)
C0523461|Alanine aminotransferase (ALT) measurement, method with pyridoxal-5'-phosphate (procedure)
C0523461|Alanine aminotransferase measurement, method with pyridoxal-5'-phosphate
C0523461|ALT measurement, method with pyridoxal-5'-phosphate
C0523462|ALT measurement, method without pyridoxal-5'-phosphate (procedure)
C0523462|Alanine aminotransferase (ALT) measurement, method without pyridoxal-5'-phosphate
C0523462|Alanine aminotransferase measurement, method without pyridoxal-5'-phosphate (procedure)
C0523462|Alanine aminotransferase measurement, method without pyridoxal-5'-phosphate
C0523462|Alanine aminotransferase (ALT) measurement, method without pyridoxal-5'-phosphate (procedure)
C0523462|ALT measurement, method without pyridoxal-5'-phosphate
C0428326|Serum glutamic oxaloacetic transaminase (SGPT) - blood measurement (procedure)
C0428326|Serum glutamic oxaloacetic transaminase (SGPT) - blood measurement
C0428326|SGPT - blood measurement (procedure)
C0428326|SGPT - blood level
C0428326|SGPT - blood measurement
C0428327|ALT - blood measurement (procedure)
C0428327|Alanine aminotransferase (ALT) - blood measurement
C0428327|Liver enzymes (& blood level [ALT] or [SGPT])
C0428327|Liver enzymes (& blood level [ALT] or [SGPT]) (procedure)
C0428327|SGPT - blood level
C0428327|ALT - blood level
C0428327|Alanine aminotransferase - blood measurement
C0428327|Alanine aminotransferase (ALT) - blood measurement (procedure)
C0428327|Alanine aminotransferase - blood measurement (procedure)
C0428327|ALT - blood measurement
C0428327|ALT blood measurement
C0042040|Urine bilirubin tests
C0042040|Bilirubin urine
C0042040|Urine Bilirubin Test
C0042040|Bilirubin measurement, urine
C0042040|Urine bilirubin
C0042040|Urine bilirubin level
C0042040|Bilirubin measurement, urine (procedure)
C0702270|Amniotic Fluid Bilirubin Test
C0702270|Bilirubin measurement, amniotic fluid
C0702270|Bilirubin measurement, amniotic fluid (procedure)
C1278039|serum total bilirubin
C1278039|Serum Total Bilirubin Measurement
C1278039|total serum bilirubin level
C1278039|serum total bilirubin measurement (lab test)
C1278039|Serum total bilirubin level
C1278039|Serum total bilirubin level (procedure)
C1278039|Serum bilirubin total
C1278039|Serum total bilirubin measurement (procedure)
C2711150|Measurement of total bilirubin in cord blood specimen (procedure)
C2711150|Measurement of total bilirubin in cord blood specimen
C0201913|Bilirubin; total
C0201913|Total Bilirubin Measurement
C0201913|BILIRUBIN TOTAL
C0201913|Measurement of total bilirubin
C0201913|Total bilirubin
C0201913|Total bilirubin (& level) (procedure)
C0201913|Bilirubin, total measurement
C0201913|Bilirubin, total measurement (procedure)
C0201913|Total bilirubin (& level)
C0201913|Bilirubin
C0201913|BILI
C0201913|Total bilirubin level
C0201913|Bilirubin, total measurement (procedure) [Ambiguous]
C0373554|Bilirubin; feces, qualitative
C0373554|BILIRUBIN FECES QUALITATIVE
C0373554|FECAL BILIRUBIN TEST
C0697273|Bilirubin; direct
C0697273|Bilirubin conjugated
C0697273|BILIRUBIN DIRECT
C0697273|Conjugated Bilirubin test
C1278036|Plasma total bilirubin level (procedure)
C1278036|Plasma total bilirubin level
C1278036|Plasma bilirubin total
C1278036|Plasma Total Bilirubin Test
C1278036|Plasma total bilirubin measurement (procedure)
C1278036|Plasma total bilirubin measurement
C0201917|Baby bilirubin measurement
C0201917|Bilirubin, neonatal measurement
C0201917|Bilirubin, neonatal measurement (procedure)
C0201917|Total bilirubin, neonatal measurement
C0201917|Microbilirubin measurement
C0201917|Total bilirubin, neonatal measurement (procedure)
C0428441|bilirubin
C0428441|serum bilirubin measurement (lab test)
C0428441|Serum bilirubin (& level) (procedure)
C0428441|Bilirubin - serum
C0428441|Serum bilirubin NOS (procedure)
C0428441|Serum bilirubin NOS
C0428441|Serum bilirubin level
C0428441|Serum bilirubin (& level)
C0428441|Serum bilirubin
C0428441|SB - Serum bilirubin
C0428441|Serum bilirubin measurement (procedure)
C0428441|Serum bilirubin measurement
C1278064|Serum methaemalbumin level (procedure)
C1278064|Serum methaemalbumin level
C1278064|Serum methemalbumin level
C1278064|Serum methaemalbumin measurement
C1278064|Serum methemalbumin measurement (procedure)
C1278064|Serum methemalbumin measurement
C2711642|Measurement of albumin gradient between serum specimen and ascitic fluid specimen (procedure)
C2711642|Measurement of albumin gradient between serum specimen and ascitic fluid specimen
C2711642|Serum ascites albumin gradient
C2097241|serum albumin/globulin ratio (lab test)
C2097241|serum albumin/globulin ratio
C2097241|albumin/globulin ratio
C2097242|serum albumin-globulin capacity (lab test)
C2097242|serum albumin-globulin capacity
C2097242|albumin-globulin capacity
C2732844|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 120 minutes after 75 gram oral glucose challenge (procedure)
C2732844|Quantitative measurement of glucose in serum or plasma specimen 120 minutes after 75 gram oral glucose challenge
C2732844|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 120 minutes after 75 gram oral glucose challenge
C2733143|Quantitative measurement of substance rate of glucose excretion in urine specimen
C2733143|Quantitative measurement of substance rate of glucose excretion in urine
C2733143|Quantitative measurement of substance rate of glucose excretion in urine specimen (procedure)
C2732700|Quantitative measurement of mass concentration of glucose in pericardial fluid specimen (procedure)
C2732700|Quantitative measurement of mass concentration of glucose in pericardial fluid specimen
C2732700|Quantitative measurement of glucose in pericardial fluid specimen
C2732794|Quantitative measurement of mass concentration of glucose in 1 hour postprandial urine specimen (procedure)
C2732794|Quantitative measurement of mass concentration of glucose in 1 hour postprandial urine specimen
C2732794|Quantitative measurement of glucose in 1 hour postprandial urine specimen
C2732897|Quantitative measurement of glucose in peritoneal dialysis fluid specimen
C2732897|Quantitative measurement of mass concentration of glucose in peritoneal dialysis fluid specimen
C2732897|Quantitative measurement of mass concentration of glucose in peritoneal dialysis fluid specimen (procedure)
C2732804|Quantitative measurement of mass concentration of glucose in synovial fluid specimen
C2732804|Quantitative measurement of glucose in synovial fluid specimen
C2732804|Quantitative measurement of mass concentration of glucose in synovial fluid specimen (procedure)
C2733070|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 6 hours after glucose challenge
C2733070|Quantitative measurement of mass concentration of glucose in serum or plasma specimen 6 hours after glucose challenge (procedure)
C2733070|Quantitative measurement of glucose in serum or plasma specimen 6 hours after glucose challenge
C2732796|Quantitative measurement of mass rate of excretion of glucose in 24 hour urine specimen
C2732796|Quantitative measurement of mass rate of excretion of glucose in 24 hour urine specimen (procedure)
C2732796|Quantitative measurement of glucose in 24 hour urine specimen
C2732716|Quantitative measurement of mass concentration of glucose in postcalorie fasting serum or plasma specimen
C2732716|Quantitative measurement of mass concentration of glucose in postcalorie fasting serum or plasma
C2732716|Quantitative measurement of mass concentration of glucose in postcalorie fasting serum or plasma specimen (procedure)
C2732249|Quantitative measurement of mass concentration of glucose in pleural fluid specimen (procedure)
C2732249|Quantitative measurement of mass concentration of glucose in pleural fluid specimen
C2732249|Quantitative measurement of glucose in pleural fluid specimen
C0201899|serum SGOT
C0201899|serum AST
C0201899|Aspartate aminotransferase
C0201899|GOT
C0201899|AST
C0201899|Aspartate Aminotransferase Measurement
C0201899|Transferase; aspartate amino (AST) (SGOT)
C0201899|TRANSFERASE ASPARTATE AMINO AST SGOT
C0201899|Liver enzyme (SGOT), level
C0201899|Measurement of aspartate amino transferase
C0201899|Measurement of aspartate amino transferase (AST) (SGOT)
C0201899|AST - aspartate transam SGOT (& level) (procedure)
C0201899|AST - aspartate transam SGOT (& level)
C0201899|Transferase (ast) (sgot)
C0201899|SGOT
C0201899|ASPT
C0201899|Aspartate transferase
C0201899|Asp transferase
C0201899|Serum glutamic-oxaloacetic transferase
C0201899|Glutamic-oxaloacetic transferase
C0201899|Serum Aspartate Transaminase Test
C0201899|AST measurement
C0201899|Glutamic oxaloacetic transaminase measurement
C0201899|GOT measurement
C0201899|SGOT measurement
C0201899|Aspartate aminotransferase measurement (procedure)
C1261155|AST serum measurement (procedure)
C1261155|Serum Aspartate Transaminase Measurement
C1261155|Serum Aspartate Aminotransferase Measurement
C1261155|Serum SGOT Measurement
C1261155|AST serum level
C1261155|AST serum level (procedure)
C1261155|Aspartate aminotransferase (AST) serum measurement (procedure)
C1261155|Aspartate aminotransferase serum measurement (procedure)
C1261155|Aspartate aminotransferase (AST) serum measurement
C1261155|Aspartate aminotransferase serum measurement
C1261155|AST serum measurement
C0523517|Aspartate amino transferase/alanine amino transferase ratio measurement
C0523517|Aspartate amino transferase/alanine amino transferase ratio measurement (procedure)
C1278050|Plasma aspartate transaminase level (procedure)
C1278050|Plasma aspartate transaminase level
C1278050|Plasma aspartate transaminase measurement (procedure)
C1278050|Plasma aspartate transaminase measurement
C0523891|serum sodium
C0523891|serum Na+
C0523891|Serum Sodium Measurement
C0523891|serum sodium measurement (lab test)
C0523891|Sodium; serum, plasma or whole blood
C0523891|SODIUM SERUM PLASMA OR WHOLE BLOOD
C0523891|Measurement of sodium in serum
C0523891|Serum sodium (& level) (procedure)
C0523891|Serum sodium (& level)
C0523891|Sodium - serum
C0523891|Serum Sodium Ion Test
C0523891|Sodium measurement, serum
C0523891|Serum sodium level
C0523891|Sodium measurement, serum (procedure)
C0523891|ASSAY OF SERUM SODIUM
C0523891|Serum sodium each test
C0523891|serum sodium ea.tst
C2016757|sodium measurement from other source (lab test)
C2016757|sodium measurement from other source
C2016757|sodium level from source other than urine
C2702997|whole blood sodium measurement (lab test)
C2702997|whole blood sodium measurement
C2702997|Measurement of sodium in whole blood
C3161784|serum sodium after fludrocortisone
C3161784|serum sodium after fludrocortisone (lab test)
C3161785|serum sodium after demeclocyline
C3161785|serum sodium after demeclocyline (lab test)
C0302353|serum K+
C0302353|Serum Potassium
C0302353|Serum Potassium Measurement
C0302353|serum potassium measurement (lab test)
C0302353|potassium level
C0302353|POTASSIUM SERUM PLASMA/WHOLE BLOOD
C0302353|Potassium; serum, plasma or whole blood
C0302353|Measurement of potassium in serum
C0302353|Potassium - serum
C0302353|Serum potassium (& level) (procedure)
C0302353|Serum potassium (& level)
C0302353|Serum potassium level
C0302353|Serum potassium measurement (procedure)
C0302353|ASSAY OF SERUM POTASSIUM
C0553704|Potassium, increased level
C0553704|Serum potasium increased
C0553704|Serum potassium increased
C0553704|Potassium serum increased
C2229880|serum total body potassium measurement
C2229880|serum total body potassium measurement (lab test)
C2229880|total body potassium level
C0373708|Protein, total, except by refractometry; serum, plasma or whole blood
C0373708|PROTEIN XCPT REFRACTOMETRY SERUM PLASMA/WHL BLD
C0373708|ASSAY OF PROTEIN SERUM
C4048459|OBSTETRIC PANEL
C4048459|Obstetric panel This panel must include the following: Blood count, complete (CBC), automated and automated differential WBC count (85025 or 85027 and 85004) OR Blood count, complete (CBC), automated (85027) and appropriate manual differential WBC count (85007 or 85009) Hepatitis B surface antigen (HBsAg) (87340) Antibody, rubella (86762) Syphilis test, non-treponemal antibody; qualitative (eg, VDRL, RPR, ART) (86592) Antibody screen, RBC, each serum technique (86850) Blood typing, ABO (86900) AND Blood typing, Rh (D) (86901)
C0812553|ACUTE HEPATITIS PANEL
C0812553|Acute hepatitis panel This panel must include the following: Hepatitis A antibody (HAAb), IgM antibody (86709) Hepatitis B core antibody (HBcAb), IgM antibody (86705) Hepatitis B surface antigen (HBsAg) (87340) Hepatitis C antibody (86803)
C1964052|BASIC METABOLIC PANEL CALCIUM IONIZED
C1964052|METABOLIC PANEL IONIZED CA
C1964052|BMP with ionized calcium
C1964052|basic metabolic panel with ionized calcium (lab test)
C1964052|basic metabolic panel with ionized calcium
C1964052|Basic metabolic panel (Calcium, ionized) This panel must include the following: Calcium, ionized (82330) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Potassium (84132) Sodium (84295) Urea Nitrogen (BUN) (84520)
C3836932|lipids test panel serum or plasma
C3836932|lipids test panel serum or plasma (lab test)
C0430044|fasting lipid panel (lab test)
C0430044|fasting lipid panel
C0430044|lipids test panel fasting
C0430044|Fasting lipid profile
C0430044|FLP - Fasting lipid profile
C0430044|Fasting lipid profile (procedure)
C0523942|Triglyceride and ester in HDL measurement (procedure)
C0523942|Triglyceride and ester in high density lipoprotein measurement (procedure)
C0523942|Triglyceride and ester in high density lipoprotein measurement
C0523942|Triglyceride and ester in HDL measurement
C0523943|Triglyceride and ester in intermediate density lipoprotein measurement (procedure)
C0523943|Triglyceride and ester in IDL measurement (procedure)
C0523943|Triglyceride and ester in intermediate density lipoprotein measurement
C0523943|Triglyceride and ester in IDL measurement
C0523944|Triglyceride and ester in low density lipoprotein measurement
C0523944|Triglyceride and ester in LDL measurement (procedure)
C0523944|Triglyceride and ester in low density lipoprotein measurement (procedure)
C0523944|Triglyceride and ester in LDL measurement
C0523945|Triglyceride and ester in VLDL measurement (procedure)
C0523945|Triglyceride and ester in very low density lipoprotein measurement
C0523945|Triglyceride and ester in very low density lipoprotein measurement (procedure)
C0523945|Triglyceride and ester in VLDL measurement
C0519823|METABOLIC PANEL TOTAL CA
C0519823|BASIC METABOLIC PANEL CALCIUM TOTAL
C0519823|Basic metabolic panel (Calcium, total) This panel must include the following: Calcium, total (82310) Carbon dioxide (bicarbonate) (82374) Chloride (82435) Creatinine (82565) Glucose (82947) Potassium (84132) Sodium (84295) Urea nitrogen (BUN) (84520)
C0812554|HEPATIC FUNCTION PANEL
C0812554|Hepatic function panel This panel must include the following: Albumin (82040) Bilirubin, total (82247) Bilirubin, direct (82248) Phosphatase, alkaline (84075) Protein, total (84155) Transferase, alanine amino (ALT) (SGPT) (84460) Transferase, aspartate amino (AST) (SGOT) (84450)
C0812554|Hepatic function panel This panel must include the following: Albumin (82040) Bilirubin, total (82247) Bilirubin, direct (82248) Phosphatase, alkaline (84075) Protein, total (84155) Transferase, alanine amino (ALT) (SGPT) (84460) Transferase, aspartate amino (AST) (SGOT)
C0812554|Liver function blood test panel
C4050228|OBSTETRIC PANEL
C4050228|Obstetric panel (includes HIV testing) This panel must include the following: Blood count, complete (CBC), and automated differential WBC count (85025 or 85027 and 85004) OR Blood count, complete (CBC), automated (85027) and appropriate manual differential WBC count (85007 or 85009) Hepatitis B surface antigen (HBsAg) (87340) HIV-1 antigen(s), with HIV-1 and HIV-2 antibodies, single result (87389) Antibody, rubella (86762) Syphilis test, non-treponemal antibody; qualitative (eg, VDRL, RPR, ART) (86592) Antibody screen, RBC, each serum technique (86850) Blood typing, ABO (86900) AND Blood typing, Rh (D) (86901)
C0430174|Metabolic function tested
C0430174|Metabolic function test NOS (procedure)
C0430174|Metabolic function test NOS
C0430174|Metabolic function tested (finding)
C0430174|Metabolic function test
C0430174|Metabolic function test (procedure)
C0430174|Metabolic function tested (procedure)
C2368348|basic metabolic panel and renal function tests (lab test)
C2368348|basic metabolic panel and renal function tests
C0430175|Chem. metab. function test NOS
C0430175|Chem. metab. function test NOS (procedure)
C0006779|Calorimetry
C0006779|Calorimetry (procedure)
C0204047|Ischaemic forearm exercise test
C0204047|Ischaemic forearm exercise test (procedure)
C0204047|Ischemic forearm exercise test
C0204047|Ischaemic forearm exercise test [Ambiguous]
C0204047|Ischemic forearm exercise test (procedure)
C0204047|Ischemic forearm exercise test (regime/therapy)
C0204048|Ischemic limb exercise with electromyography and lactic acid determination (procedure)
C0204048|Ischemic limb exercise with electromyography and lactic acid determination
C0204048|Ischemic limb exercise with EMG and lactic acid determination
C0204048|Ischaemic limb exercise with EMG and lactic acid determination
C0204048|Ischemic limb exercise with EMG and lactic acid determination (procedure)
C0204048|Ischemic limb exercise with EMG and lactic acid determination (regime/therapy)
C1283822|Ischaemic lactate test
C1283822|Ischemic lactate test
C1283822|Ischemic lactate test (procedure)
C0430180|Body water test
C0430180|Body water test (procedure)
C0430177|Flush provocation test
C0430177|Flush provocation test (procedure)
C0430603|Metabolic function not tested (situation)
C0430603|Metabolic function not tested (procedure)
C0430603|Metabolic function not tested
C0430178|Nicotinic acid loading test
C0430178|Nicotinic acid loading test (procedure)
C0430176|Nitrogen balance test
C0430176|Nitrogen balance test (procedure)
C1273413|Endocrine studies
C1273413|Endocrine studies (procedure)
