C0011849|Diabetes Mellitus
C0011880|Acidoses, Diabetic
C0011880|Diabetic Acidoses
C0011880|Diabetic Ketoacidoses
C0011880|Diabetic Ketoacidosis
C0011880|Ketoacidoses, Diabetic
C0011880|Ketosis, Diabetic
C0011880|diabetic acidosis
C0011880|Diabetes mellitus with ketoacidosis
C0011880|Ketoacidosis in diabetes mellitus (disorder)
C0011880|Ketoacidosis in diabetes mellitus
C0011880|diabetes with ketoacidosis
C0011880|diabetes mellitus with ketoacidosis (diagnosis)
C0011880|Acidosis, Diabetic
C0011880|Diabetic Ketosis
C0011880|Ketoacidosis, Diabetic
C0011880|Diabetic Ketoacidosis [Disease/Finding]
C0011880|Diabetes mellitus NOS with ketoacidosis (disorder)
C0011880|Ketoacidosis - diabetic
C0011880|Diabetes mellitus NOS with ketoacidosis
C0011880|Diabetes mellitus (& [ketoacidosis]) (disorder)
C0011880|Diabetes mellitus (& [ketoacidosis])
C0011880|Diabetes with ketoacidosis (disorder)
C0011880|DKA - Diabetic ketoacidosis
C0011880|DKA
C0011880|Ketoacidosis (diabetic)
C0011880|Acidosis diabetic
C0011880|Diabetic acidosis without coma
C0011880|Diabetic ketosis without coma
C0011880|Diabetic acidosis, NOS
C0011880|Diabetic Ketoses
C0011880|Ketoses, Diabetic
C0011875|Angiopathies, Diabetic
C0011875|Diabetic Angiopathies
C0011875|Angiopathy, Diabetic
C0011875|Diabetic Angiopathy
C0011875|Diabetic Angiopathies [Disease/Finding]
C0011875|Diabetic Vascular Diseases
C0011875|Diabetic Vascular Complications
C0011875|Diabetic vascular disorder
C0011875|Diabetic vascular disorder NOS
C0011875|diabetes; angiopathy (manifestation)
C0011875|angiopathy; diabetes (manifestation)
C0011875|Diabetic Vascular Complication
C0011875|Diabetic Vascular Disease
C0011875|Vascular Complication, Diabetic
C0011875|Vascular Complications, Diabetic
C0011875|Vascular Disease, Diabetic
C0011875|Vascular Diseases, Diabetic
C0011881|Diabetic Nephropathies
C0011881|Nephropathies, Diabetic
C0011881|Diabetes with renal manifestations
C0011881|Nephropathy, Diabetic
C0011881|diabetic nephropathy
C0011881|Renal disorder associated with diabetes mellitus
C0011881|diabetic nephropathy (diagnosis)
C0011881|Diabetic Kidney Disease
C0011881|Diabetic Nephropathies [Disease/Finding]
C0011881|Nephropathy;diabetic
C0011881|diabetes with renal manifestations (diagnosis)
C0011881|Diabetic Kidney Problems
C0011881|Diabetes + nephropathy
C0011881|Diabetes with renal manifestations (disorder)
C0011881|Nephropathy - diabetic
C0011881|-- Diabetic Kidney Disease
C0011881|Diabetic nephropathy NOS
C0011881|Diabetic renal disease
C0011881|Diabetic renal disease (disorder)
C0011881|diabetes; nephropathy (manifestation)
C0011881|nephropathy; diabetes (manifestation)
C0011881|Diabetic Kidney Diseases
C0011881|Kidney Disease, Diabetic
C0011881|Kidney Diseases, Diabetic
C0011882|Diabetic Neuropathies
C0011882|Neuropathies, Diabetic
C0011882|Diabetes with neurological manifestations
C0011882|Diabetic Neuropathy
C0011882|Neuropathy, Diabetic
C0011882|Diabetic Neuropathies [Disease/Finding]
C0011882|Neuropathy;diabetic
C0011882|Neuropathy - diabetic
C0011882|Diabetes + neuropathy
C0011882|Diabetic neuropathy (disorder)
C0011882|Diabetes mellitus with neuropathy
C0011882|Diabetes mellitus with neurological manifestation
C0011882|Diabetes mellitus NOS with neurological manifestation (disorder)
C0011882|Diabetes mellitus NOS with neurological manifestation
C0011882|neuropathy; diabetes (manifestation)
C0011882|Diabetic neuropathy (disorder) [Ambiguous]
C0085207|Diabetes, Gestational
C0085207|Diabetes, Pregnancy Induced
C0085207|Gestational Diabetes Mellitus
C0085207|Pregnancy-Induced Diabetes
C0085207|GDM
C0085207|Diabetes mellitus arising in pregnancy
C0085207|Gestational diabetes
C0085207|Diabetes in Pregnancy
C0085207|DIABETES PREGN IND
C0085207|gestational diabetes mellitus (diagnosis)
C0085207|Gestational diabetes mellitus NOS
C0085207|Diabetes, Pregnancy-Induced
C0085207|Diabetes, Gestational [Disease/Finding]
C0085207|Diabetes Mellitus, Gestational
C0085207|Diabetes;during pregnancy
C0085207|Diabetes and Pregnancy
C0085207|Gestational diabetes mellitus (disorder)
C0085207|Maternal gestational diabetes mellitus
C0085207|Maternal gestational diabetes mellitus (disorder)
C0085207|-- Gestational Diabetes
C0085207|Maternal diabetes
C0085207|Diabetes mellitus gestational
C0085207|GDM - Gestational diabetes mellitus
C0085207|Gestational diabetes mellitus, NOS
C0011854|Brittle Diabetes Mellitus
C0011854|Diabetes Mellitus, Insulin-Dependent
C0011854|Diabetes Mellitus, Juvenile Onset
C0011854|Diabetes Mellitus, Ketosis Prone
C0011854|IDDM
C0011854|Insulin-Dependent Diabetes Mellitus
C0011854|Juvenile-Onset Diabetes Mellitus
C0011854|Ketosis-Prone Diabetes Mellitus
C0011854|Diabetes Mellitus, Insulin Dependent
C0011854|insulin dependent diabetes mellitus
C0011854|Diabetes Mellitus, Sudden Onset
C0011854|Mellitus, Sudden-Onset Diabetes
C0011854|Sudden-Onset Diabetes Mellitus
C0011854|JOD
C0011854|IDDM1
C0011854|INSULIN-DEPENDENT DIABETES MELLITUS 1
C0011854|Insulin-dependent diabetes mellitus (type I)
C0011854|DIABETES MELLITUS, INSULIN-DEPENDENT, 1
C0011854|DIABETES MELLITUS TYPE 01
C0011854|insulin dependent diabetes
C0011854|type I diabetes mellitus
C0011854|juvenile diabetes mellitus
C0011854|ketosis prone diabetes
C0011854|IDD
C0011854|Type 1 diabetes mellitus
C0011854|Type 1 Diabetes
C0011854|Type I Diabetes
C0011854|Juvenile Diabetes
C0011854|DIABETES MELLITUS, KETOSIS-PRONE
C0011854|KPD
C0011854|brittle diabetes (mellitus)
C0011854|juvenile onset diabetes (mellitus)
C0011854|ketosis-prone diabetes (mellitus)
C0011854|Diabetes Mellitus, Type 1 [Disease/Finding]
C0011854|Diabetes Mellitus, Brittle
C0011854|Diabetes Mellitus, Type 1
C0011854|Diabetes Mellitus, Juvenile-Onset
C0011854|Diabetes Mellitus, Sudden-Onset
C0011854|Diabetes Mellitus, Type I
C0011854|Diabetes;Type 1
C0011854|Diabetes;insulin dependent
C0011854|Diabetes;juvenile onset
C0011854|Insulin Dependent Diabetes Mellitus 1
C0011854|Juvenile Onset Diabetes
C0011854|Diabetes, Juvenile-Onset
C0011854|Juvenile-Onset Diabetes
C0011854|Diabetes Type 1
C0011854|Insulin-dependent diabetes
C0011854|Diabetes mellitus: [juvenile] or [insulin dependent]
C0011854|Diabetes mellitus - juvenile
C0011854|Diabetes mellitus: [juvenile] or [insulin dependent] (disorder)
C0011854|Diabetes mellitus type 1
C0011854|Juvenile onset diabetes mellitus
C0011854|Type I diabetes mellitus (disorder)
C0011854|IDDM - Insulin-dependent diabetes mellitus
C0011854|Insulin dependent diabetes mel
C0011854|-- Diabetes Type 1
C0011854|Diabetes mellitus Type I
C0011854|Type 1 diabetes mellitus (diagnosis)
C0011854|Diabetes mellitus juvenile onset
C0011854|Diabetes mellitus insulin-dependent
C0011854|Insulin dependent diabetic
C0011854|Diabetes mellitus type 1 (disorder)
C0011854|diabetes; insulin-dependent
C0011854|diabetes; juvenile-onset
C0011854|diabetes; ketosis-prone
C0011854|diabetes; type I
C0011854|insulin-dependent; diabetes
C0011854|juvenile-onset; diabetes
C0011854|ketosis, prone; diabetes
C0011854|type I; diabetes
C0011854|juvenile onset of diabetes
C0011860|Adult-Onset Diabetes Mellitus
C0011860|Diabetes Mellitus, Adult Onset
C0011860|Diabetes Mellitus, Ketosis Resistant
C0011860|Diabetes Mellitus, Non-Insulin-Dependent
C0011860|Ketosis-Resistant Diabetes Mellitus
C0011860|NIDDM
C0011860|Non-Insulin-Dependent Diabetes Mellitus
C0011860|Stable Diabetes Mellitus
C0011860|Diabetes Mellitus, Maturity Onset
C0011860|Maturity Onset Diabetes Mellitus
C0011860|noninsulin dependent diabetes mellitus
C0011860|Diabetes Mellitus, Slow Onset
C0011860|Slow-Onset Diabetes Mellitus
C0011860|Noninsulin-dependent diabetes mellitus
C0011860|Diabetes mellitus, noninsulin-dependent
C0011860|DIABETES MELLITUS TYPE 02
C0011860|adult onset diabetes mellitus
C0011860|type II diabetes mellitus
C0011860|ketosis resistant diabetes
C0011860|Diabetes mellitus non insulin-dep
C0011860|Type 2 diabetes mellitus
C0011860|AODM
C0011860|type 2 diabetes
C0011860|non-insulin dependent diabetes mellitus
C0011860|Adult-Onset Diabetes
C0011860|Type 2 Diabetes Mellitus Non-Insulin Dependent
C0011860|Type II Diabetes
C0011860|T2D
C0011860|T2DM - Type 2 Diabetes mellitus
C0011860|Diabetes, Type 2
C0011860|Diabetes Mellitus, Stable
C0011860|MODY
C0011860|Diabetes Mellitus, Type 2
C0011860|Diabetes Mellitus, Ketosis-Resistant
C0011860|Diabetes Mellitus, Non Insulin Dependent
C0011860|Diabetes Mellitus, Slow-Onset
C0011860|Diabetes Mellitus, Noninsulin Dependent
C0011860|Diabetes Mellitus, Type 2 [Disease/Finding]
C0011860|Maturity-Onset Diabetes Mellitus
C0011860|Diabetes Mellitus, Maturity-Onset
C0011860|Diabetes Mellitus, Adult-Onset
C0011860|Diabetes Mellitus, Type II
C0011860|Diabetes;Type 2
C0011860|Diabetes;adult onset
C0011860|Diabetes;non insulin depend
C0011860|Diabetes mellitus (NIDDM)
C0011860|Maturity-Onset Diabetes
C0011860|Diabetes Type 2
C0011860|Diabetes mellitus type 2
C0011860|Diabetes mellitus - adult onset
C0011860|Diabetes mellitus: [adult onset] or [noninsulin dependent]
C0011860|Diabetes mellitus: [adult onset] or [noninsulin dependent] (disorder)
C0011860|Diabetes mellitus -adult onset
C0011860|NIDDM - Non-insulin dependent diabetes mellitus
C0011860|Type II diabetes mellitus (disorder)
C0011860|Maturity onset diabetes
C0011860|Noninsulin dependent diab.mell
C0011860|Non-insulin-dependent diabetes
C0011860|-- Diabetes Type 2
C0011860|Noninsulin Dependent Diabetes
C0011860|Type I I Diabetes
C0011860|Adult Onset Diabetes
C0011860|Noninsulin dependent diabetes mellitus (NIDDM)
C0011860|Noninsulin-dependent diabetes
C0011860|Diabetes mellitus Type II
C0011860|NIDDM diabetes mellitus
C0011860|Type 2 diabetes mellitus (diagnosis)
C0011860|Diabetes mellitus maturity onset
C0011860|Diabetes mellitus non-insulin-dependent
C0011860|Diabetes mellitus type 2 (disorder)
C0011860|diabetes
C0011860|NIDDM; diabetes
C0011860|diabetes; NIDDM
C0011860|diabetes; adult-onset
C0011860|diabetes; maturity-onset
C0011860|diabetes; non-insulin-dependent
C0011860|diabetes; nonketotic
C0011860|diabetes; type II
C0011860|maturity-onset; diabetes
C0011860|non-insulin-dependent; diabetes
C0011860|nonketotic; diabetes
C0011860|adult-onset; diabetes
C0011860|type II; diabetes
C0011860|NCDMM
C0011860|Non-Insulin Dependent Diabetes
C0011860|non insulin dependent diabetes
C0362046|Prediabetic State
C0362046|Prediabetic States
C0362046|State, Prediabetic
C0362046|States, Prediabetic
C0362046|Prediabetes
C0362046|Prediabetic State [Disease/Finding]
C0362046|Pre diabetes
C0362046|Prediabetes (disorder)
C0362046|Pre-diabetic
C0362046|Borderline diabetes
C0362046|Pre-diabetes
C0362046|Prediabetes (finding)
C0362046|Prediabetes syndrome
C0362046|Pre-diabetes NOS
C0271646|drug related diabetes mellitus
C0271646|Drug-induced diabetes mellitus (disorder)
C0271646|Drug-induced diabetes mellitus
C0597655|virus related diabetes mellitus
C0920358|diabetic ophthalmopathy
C0853897|Diabetic cardiomyopathy
C0853897|Diabetic Cardiomyopathies
C0853897|Cardiomyopathy, Diabetic
C0853897|Cardiomyopathies, Diabetic
C0853897|Diabetic Cardiomyopathies [Disease/Finding]
C0348447|Other specified diabetes mellitus
C0348447|[X]Other specified diabetes mellitus
C0348447|[X]Other specified diabetes mellitus (disorder)
C0271641|Malnutrition-related diabetes mellitus
C0271641|Diabetes mellitus malnutrition-related
C0271641|Malnutrition-related diabetes mellitus (disorder)
C0271641|malnutrition-related diabetes mellitus (diagnosis)
C0271641|diabetes mellitus secondary malnutrition-related
C0271641|MRDM
C0271641|Malnutrition related diabetes mellitus
C0271641|Malnutrition related diabetes mellitus (disorder)
C0271641|diabetes; malnutrition-related
C0271641|malnutrition; diabetes
C0011849|Diabetes Mellitus
C0011849|Unspecified diabetes mellitus
C0011849|diabetes mellitus (diagnosis)
C0011849|DM
C0011849|diabetes NOS
C0011849|Diabetes Mellitus [Disease/Finding]
C0011849|Diabetes mellitus (E08-E13)
C0011849|Diabetes
C0011849|Diabetes mellitus (disorder)
C0011849|Diabetes mellitus NOS
C0011849|Diabetes Melllitus
C0011849|Med: Diabetes mellitus
C0011849|DM - Diabetes mellitus
C0011849|Diabetes mellitus, NOS
C0348939|Unspecified diabetes mellitus with multiple complications
C0348939|Unspecified diabetes mellitus with multiple complications (disorder)
C0348450|Unspecified diabetes mellitus with renal complications
C0348450|[X]Unspecified diabetes mellitus with renal complications (disorder)
C0348450|[X]Unspecified diabetes mellitus with renal complications
C0494295|Unspecified diabetes mellitus with coma
C0494296|Unspecified diabetes mellitus with ketoacidosis
C2362567|Unspecified diabetes mellitus with neurological complications
C1744704|Unspecified diabetes mellitus with ophthalmic complications
C0494300|Unspecified diabetes mellitus with other specified complications
C0011871|Unspecified diabetes mellitus with peripheral circulatory complications
C0011871|Diabetic peripheral angiopathy
C0011871|diabetes mellitus with peripheral circulatory disorder
C0011871|diabetes mellitus with peripheral circulatory disorder (diagnosis)
C0011871|diabetes with peripheral circulatory disorder
C0011871|Diabetes with peripheral circulatory disorders
C0011871|Diabetes mellitus with peripheral circulatory disorder (disorder)
C0011871|Diabetes with peripheral circulatory disorders (disorder)
C0011871|Diabetes mellitus NOS with peripheral circulatory disorder (disorder)
C0011871|Diabetes mellitus NOS with peripheral circulatory disorder
C0011871|Diabetes + periph.circulat.dis
C0011871|Diabetic peripheral vascular disease
C0011871|Diabetic peripheral angiopathy (disorder)
C0011871|Diabetic peripheral vascular disorder
C0342257|Disorder associated with diabetes mellitus
C0342257|Unspecified diabetes mellitus with unspecified complications
C0342257|DIABETES COMPL
C0342257|COMPL DIABETES MELLITUS
C0342257|DIABETES RELAT COMPL
C0342257|DIABETIC COML
C0342257|diabetes mellitus with complication (diagnosis)
C0342257|diabetes mellitus with complication
C0342257|Diabetes with unspecified complications
C0342257|Diabetic complications
C0342257|Diabetes mellitus with complications
C0342257|Diabetes Complication
C0342257|Diabetes Complications
C0342257|Diabetes-Related Complications
C0342257|Diabetes Complications [Disease/Finding]
C0342257|Complications of Diabetes Mellitus
C0342257|Diabetes;complicated
C0342257|Diabetes mellitus NOS with unspecified complication
C0342257|Diabetes mellitus with unspecified complication
C0342257|Diabetes with diabetic complications
C0342257|Diabetes mellitus with unspecified complication (disorder)
C0342257|Diabetes mellitus with complication (disorder)
C0342257|Diabetes mellitus NOS with unspecified complication (disorder)
C0342257|Diabetes--Complications
C0342257|Diabetes with unspecified complication
C0342257|Diabetic complication
C0342257|Diabetic complication NOS
C0342257|Diabetic complication (disorder)
C0342257|Diabetic complication, NOS
C0342257|Diabetes Mellitus Complications
C0342257|Diabetes Mellitus Complication
C0342257|Diabetes Related Complications
C0342257|Diabetes-Related Complication
C0342257|complicated diabetes
C0271635|Diabetes mellitus without complication
C0271635|Unspecified diabetes mellitus without complications
C0271635|diabetes mellitus without complication (diagnosis)
C0271635|Diabetes mellitus NOS with no mention of complication
C0271635|Diabetes mellitus with no mention of complication (disorder)
C0271635|Diabetes mellitus with no mention of complication
C0271635|Diabetes mellitus NOS with no mention of complication (disorder)
C0271635|Diabetes mellitus without mention of complication
C0271635|Diabetes mellitus without complication (disorder)
C0011853|Diabetes Mellitus, Experimental
C0011853|EXPER DIABETES MELLITUS
C0011853|DIABETES MELLITUS EXPER
C0011853|Experimental Diabetes Mellitus
C0011853|Diabetes Mellitus, Experimental [Disease/Finding]
C2711205|Multiple complications due to diabetes mellitus (disorder)
C2711205|Multiple complications due to diabetes mellitus
C0265344|DONOHUE SYNDROME
C0265344|Leprechaunisms
C0265344|Syndrome, Donohue
C0265344|Donohue Syndrome [Disease/Finding]
C0265344|Leprechaunism
C0265344|Leprechaunism syndrome
C0265344|Donohue's syndrome
C0265344|Leprechaunism syndrome (disorder)
C0265344|Donohue
C2827448|Childhood Diabetes Mellitus
C2873880|Diabetes mellitus due to underlying condition
C2873948|Drug or chemical induced diabetes mellitus
C2919615|Posttransplant diabetes mellitus (disorder)
C2919615|Posttransplant diabetes mellitus
C0554876|poorly controlled diabetes mellitus (diagnosis)
C0554876|diabetes mellitus poorly controlled
C0554876|poorly controlled diabetes mellitus
C1720078|Diabetic neurologic disease
C1720078|Neurologic complication of diabetes mellitus
C1720078|Neurologic disorder associated with diabetes mellitus (disorder)
C1720078|Neurologic disorder associated with diabetes mellitus
C1720078|diabetes mellitus with neurological complications (diagnosis)
C1720078|diabetes with neurological complications
C1720078|diabetes mellitus with neurological complications
C0342245|Diabetes with ophthalmic manifestations
C0342245|diabetes mellitus with ophthalmic manifestations (diagnosis)
C0342245|diabetes mellitus with ophthalmic manifestations
C0342245|Diabetic Eye Disease
C0342245|Diabetic Eye Problems
C0342245|Diabetes mellitus NOS with ophthalmic manifestation
C0342245|Diabetes mellitus with ophthalmic manifestation (disorder)
C0342245|Diabetes mellitus with ophthalmic manifestation
C0342245|Diabetes + eye manifestation
C0342245|Diabetes mellitus NOS with ophthalmic manifestation (disorder)
C0342245|Diabetic eye disease NOS
C0342245|Ophthalmic manifestations of diabetes
C0342245|Diabetic oculopathy (disorder)
C0342245|Diabetic oculopathy
C0342245|Diabetic oculopathy, NOS
C0342245|Diabetic eye disease, NOS
C2062378|diabetes mellitus under control
C2062378|diabetes mellitus under control (diagnosis)
C0553772|diabetes mellitus with hyperosmolar nonketotic state (diagnosis)
C0553772|diabetes mellitus with hyperosmolar nonketotic state
C0553772|hyperglycemic hyperosmolar nonketotic state
C0553772|Diabetic hyperosmolar non-ketotic state
C0553772|HONKS - Diabetic hyperosmolar non-ketotic state
C0553772|Diabetic hyperosmolar non-ketotic state (disorder)
C0860163|diabetic gastropathy
C0860163|diabetes mellitus with gastropathy (diagnosis)
C0860163|diabetes mellitus with gastropathy
C0271640|Secondary diabetes mellitus
C0271640|Secondary diabetes mellitus NOS
C0271640|secondary diabetes mellitus (diagnosis)
C0271640|Secondary diabetes mellitus (disorder)
C0271640|Secondary diabetes mellitus, NOS
C0158981|Neonatal diabetes mellitus
C0158981|neonatal diabetes mellitus (diagnosis)
C0158981|Neonatal diabetes
C0158981|Neonat diabetes mellitus
C0158981|Diabetes mellitus syndrome in newborn infant
C0158981|Congenital Diabetes Mellitus
C0158981|Neonatal diabetes mellitus (disorder)
C0158981|diabetes; neonatal
C0158981|neonatal; diabetes
C0865166|Diabetic hypoglycemia NOS
C0865166|diabetes mellitus with hypoglycemia
C0865166|diabetic hypoglycemia
C0865166|diabetic hypoglycemia (diagnosis)
C2930860|Premature aging, Okamoto type
C2931057|Lipoatrophy with diabetes, hepatic steatosis, cardiomyopathy, and leukomelanodermic papules
C2931125|Feigenbaum Bergeron Richardson syndrome
C0342287|TRMA
C0342287|THIAMINE-RESPONSIVE MEGALOBLASTIC ANEMIA SYNDROME
C0342287|Thiamine responsive myelodysplasia
C0342287|Thiamine responsive megaloblastic anemia syndrome
C0342287|Abboud syndrome
C0342287|Rogers syndrome
C0342287|THMD1
C0342287|Megaloblastic Anemia, Thiamine-Responsive, With Diabetes Mellitus And Sensorineural Deafness
C0342287|Thiamine-Responsive Myelodysplasia
C0342287|Thiamine-Responsive Anemia Syndrome
C0342287|THIAMINE METABOLISM DYSFUNCTION SYNDROME 1 (MEGALOBLASTIC ANEMIA, DIABETES MELLITUS, AND DEAFNESS TYPE)
C0342287|Megaloblastic anaemia, thiamine-responsive, with diabetes mellitus and sensorineural deafness
C0342287|Megaloblastic anemia, thiamine-responsive, with diabetes mellitus and sensorineural deafness (disorder)
C2931296|Pancreatic hypoplasia diabetes heart disease
C2931296|Yorifuji Okuno syndrome
C0342286|Hypogonadism, diabetes mellitus, alopecia ,mental retardation and electrocardiographic abnormalities
C0342286|Woodhouse Sakati syndrome
C0342286|Extrapyramidal Disorder, Progressive, With Primary Hypogonadism, Mental Retardation, and Alopecia
C0342286|Hypogonadism, Alopecia, Diabetes Mellitus, Mental Retardation, and Extrapyramidal Syndrome
C0342286|Woodhouse-Sakati Syndrome
C0342286|HYPOGONADISM, ALOPECIA, DIABETES MELLITUS, MENTAL RETARDATION, DEAFNESS, AND EXTRAPYRAMIDAL SYNDROME
C0342286|Hypogonadism, diabetes mellitus, alopecia, mental retardation and electrocardiographic abnormalities (disorder)
C0342286|Hypogonadism, diabetes mellitus, alopecia, mental retardation and electrocardiographic abnormalities
C0342286|Hypogonadism, diabetes mellitus, alopecia ,mental retardation and electrocardiographic abnormalities (disorder)
C1838655|PANCREATIC BETA CELL AGENESIS WITH NEONATAL DIABETES MELLITUS
C1838655|Congenital absence of insulin-producing beta cells with diabetes mellitus
C1809475|PHOTOMYOCLONUS, DIABETES MELLITUS, DEAFNESS, NEPHROPATHY, AND CEREBRAL DYSFUNCTION
C1809475|Herrmann syndrome
C1809475|Photomyoclonus, diabetes mellitus, deafness, nephropathy and cerebral dysfunction
C1809475|Photomyoclonus, diabetes mellitus, deafness, nephropathy and cerebral dysfunction (disorder)
C2931765|Furukawa Takagi Nakao syndrome
C0431693|RENAL CYSTS AND DIABETES SYNDROME
C0431693|MODY5
C0431693|Hyperuricemic nephropathy, familial juvenile, atypical
C0431693|Glomerulocystic kidney disease, hypoplastic type
C0431693|Glomerulocystic kidney, familial hypoplastic
C0431693|Maturity-onset diabetes of the young, type 5
C0431693|Renal cysts and diabetes syndrome (disorder)
C0431693|Maturity-onset diabetes of the young, type 5 (disorder)
C0431693|Familial hypoplastic, glomerulocystic kidney
C0431693|familial hypoplastic, glomerulocystic kidney (diagnosis)
C0431693|RCAD
C0431693|maturity-onset diabetes of the young - type 5 (diagnosis)
C0431693|maturity-onset diabetes of the young - type 5
C0431693|FJHN, ATYPICAL
C0431693|CONGENITAL ANOMALIES OF THE KIDNEY AND URINARY TRACT WITH DIABETES
C0431693|CAKUT WITH DIABETES
C0431693|RCAD Syndrome
C0431693|Familial hypoplastic, glomerulocystic kidney (disorder)
C0406682|Diabetic dermopathy
C0406682|diabetes mellitus with dermatological manifestations
C0406682|diabetes mellitus with dermatological manifestations (diagnosis)
C0406682|diabetes mellitus with diabetic dermatitis
C0406682|diabetes mellitus with diabetic dermatitis (diagnosis)
C0406682|diabetic dermatitis
C0406682|Diabetic dermopathy (disorder)
C3250577|diabetes mellitus with oral cavity manifestations (diagnosis)
C3250577|diabetes mellitus with oral cavity manifestations
C0375121|diabetes mellitus with hyperosmolarity
C0375121|diabetes mellitus with hyperosmolarity (diagnosis)
C3534592|Diabetes in Children and Teens
C0011878|Diabetic Diets
C0011878|Diets, Diabetic
C0011878|diabetic diet
C0011878|diabetic diet (treatment)
C0011878|Diabetic diet (finding)
C0011878|Diabetes--Diet therapy
C0011878|Diet, Diabetic
C0011878|DD - Diabetic diet
C0011878|diabetes mellitus diet
C0524620|Syndrome X, Reaven
C0524620|dysmetabolic syndrome X
C0524620|dysmetabolic syndrome X (diagnosis)
C0524620|Insulin resistance syndrome
C0524620|Metabolic syndrome
C0524620|Metabolic Syndrome X
C0524620|Insulin Resistance Syndrome X
C0524620|Metabolic X Syndrome
C0524620|Syndrome X, Insulin Resistance
C0524620|Metabolic Syndrome X [Disease/Finding]
C0524620|Metabolic Cardiovascular Syndrome
C0524620|Reaven Syndrome X
C0524620|Syndrome X, Metabolic
C0524620|Cardiovascular Syndrome, Metabolic
C0524620|Cardiovascular Syndromes, Metabolic
C0524620|Syndrome, Metabolic Cardiovascular
C0524620|Syndrome X (Metabolic)
C0524620|Metabolic syndrome X (disorder)
C0524620|Equine metabolic syndrome
C0524620|Syndrome X, Dysmetabolic
C0524620|Syndrome, Metabolic X
C0524620|X Syndrome, Metabolic
C0524620|Reaven's syndrome
C0206172|Diabetic Foot
C0206172|Feet, Diabetic
C0206172|Foot, Diabetic
C0206172|Diabetic Feet
C0206172|Diabetic Foot [Disease/Finding]
C0206172|Diabetic foot (disorder)
C3534591|Diabetic Heart Disease
C0020616|Agents, Hypoglycemic
C0020616|Hypoglycemic Agents
C0020616|hypoglycemic agent
C0020616|Drugs, Hypoglycemic
C0020616|antihyperglycemic
C0020616|Hypoglycaemic drug
C0020616|Hypoglycemic drug
C0020616|Anti-hyperglycemics
C0020616|Agents, Antihyperglycemic
C0020616|Hypoglycemic Medicines
C0020616|Diabetes Medicines
C0020616|Drugs for hypoglycemia
C0020616|Drugs for hypoglycaemia
C0020616|Hypoglycemic product (product)
C0020616|Hypoglycaemic product
C0020616|Hypoglycemic product
C0020616|Drugs for hypoglycemia (product)
C0020616|Hypoglycemic
C0020616|Hypoglycemic agent (substance)
C0020616|Hypoglycaemic
C0020616|Antihyperglycemics
C0020616|Hypoglycemics
C0020616|Antihyperglycemic Agents
C0020616|Hypoglycemic Drugs
C0020616|Hypoglycaemic agent
C0020616|Hypoglycemic agent (product)
C0020616|Hypoglycemic drug, NOS
C0020616|Hypoglycaemic drug, NOS
C0020616|Drugs for hypoglycemia (substance)
C0020616|Hypoglycemic drug (substance)
C1456657|Diabetic Nerve Problems
C0559093|Diabetes with other complications (disorder)
C0559093|Diabetes with other complications
C0011870|Diabetes with other coma
C0011870|Diabetes with non-ketotic non-hyperosmolar coma (disorder)
C0011870|Diabetes with non-ketotic non-hyperosmolar coma
C1275078|Carpenter syndrome
C1275078|Type II Acrocephalopolysyndactyly
C1275078|Acrocephalopolysyndactyly Type II
C1275078|ACPS II
C1275078|CARPENTER SYNDROME 1
C1275078|CRPT1
C1275078|Carpenter syndrome (disorder)
C1275078|Carpenter 's Syndrome
C1275078|Carpenter's syndrome
C1275078|Carpenter's syndrome (disorder)
C1275078|Acrocephalopolysyndactyly type II (disorder)
C1275078|Acrocephalopolysyndactyly type 2
C1275078|Carpenter
C0342254|Diabetes mellitis with nephropathy NOS (disorder)
C0342254|Diabetes mellitus with renal manifestation
C0342254|Diabetes mellitus with renal manifestation (disorder)
C0342254|Diabetes mellitis with nephropathy NOS
C0342290|Abnormal metabolic state in diabetes mellitus
C0342290|Abnormal metabolic state in diabetes mellitus (disorder)
C0342264|Diabetes mellitus, juvenile type, with no mention of complication
C0342264|Diabetes mellitus, juvenile type, with no mention of complication (disorder)
C1282941|Diabetes mellitus with neurological manifestation (disorder)
C1282941|Diabetes mellitus with neurological manifestation
C1282941|diabetic neuropathy with neurological complication (diagnosis)
C1282941|diabetic neuropathy with neurological complication
C1282941|Diabetes with neurological manifestations
C1282941|Diabetic neuropathy with neurologic complication
C1282941|Diabetic neuropathy with neurologic complication (disorder)
C0342265|Diabetes mellitus, adult onset, with no mention of complication (disorder)
C0342265|Diabetes mellitus, adult onset, with no mention of complication
C0554436|Diabetic gangrene
C0554436|Gangrene associated with diabetes mellitus (disorder)
C0554436|Gangrene associated with diabetes mellitus
C0554436|Gangrene - diabetic
C0554436|Diabetes mellitus with gangrene
C0554436|Diabetes mellitus with gangrene (disorder)
C0554436|Diabetes with gangrene
C0554436|diabetic gangrene (diagnosis)
C0554436|gangrene associated with diabetes mellitus (diagnosis)
C0554436|Diabetic gangrene (disorder)
C0341893|Diabetes mellitus complicating pregnancy, childbirth, or the puerperium
C0341893|Diabetes mellitus of mother, comp pregnancy,childbirth, or the puerp, unspec as to eoc
C0341893|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as t
C0341893|Diabetes in preg-unspec
C0341893|Diabetes mellitus in pregnancy, childbirth, and the puerperium
C0341893|Unspecified diabetes mellitus in pregnancy, childbirth and the puerperium
C0341893|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care
C0341893|Diabetes mellitus of mother, complicating pregnancy, childbirth, or the puerperium, unspecified as to episode of care or not applicable
C0341893|diabetes mellitus in pregnancy, childbirth, and puerperium (diagnosis)
C0341893|diabetes mellitus in pregnancy, childbirth, and puerperium
C0341893|Diabetes mellitus during pregnancy, childbirth and the puerperium (disorder)
C0341893|Diabetes mellitus during pregnancy, childbirth and the puerperium
C0341893|Diabetes mellitus during pregnancy, childbirth or the puerperium NOS (disorder)
C0341893|Diabetes mellitus during pregnancy, childbirth or the puerperium NOS
C0341893|diabetes mellitus in mother complicating pregnancy, childbirth, and puerperium
C0341893|diabetes mellitus in mother complicating pregnancy, childbirth, and puerperium (diagnosis)
C0341893|Diabetes mellitus in mother complicating pregnancy, childbirth AND/OR puerperium (disorder)
C0341893|Diabetes mellitus in mother complicating pregnancy, childbirth AND/OR puerperium
C0341893|Diabetes mellitus in mother complicating pregnancy, childbirth or puerperium
C0341893|Gestational diabetes complicating pregnancy, childbirth, or the puerperium
C0348933|Other specified diabetes mellitus with coma
C0348933|Other specified diabetes mellitus with coma (disorder)
C0342260|Diabetes mellitus NOS with other specified manifestation (disorder)
C0342260|Diabetes mellitus with other specified manifestation (disorder)
C0342260|Diabetes mellitus NOS with other specified manifestation
C0342260|Diabetes mellitus with other specified manifestation
C0348931|Other specified diabetes mellitus with other specified complications
C0348931|Other specified diabetes mellitus with other specified complication
C0348931|Oth diabetes mellitus with other specified complication
C0348931|Other specified diabetes mellitus with other specified complications (disorder)
C0342261|Type I diabetes mellitus with other specified manifestations
C0342261|Insulin-dependent diabetes mellitus with other specified complications
C0342261|Type 1 diabetes mellitus with other specified complications
C0342261|Type 1 diabetes mellitus with other specified complication
C0342261|Diabetes mellitus, juvenile type, with other specified manifestation
C0342261|Diabetes mellitus, juvenile type, with other specified manifestation (disorder)
C0348938|Other specified diabetes mellitus with multiple complications
C0348938|Other specified diabetes mellitus with multiple complications (disorder)
C0342262|Type II diabetes mellitus with other specified manifestations
C0342262|Non-insulin-dependent diabetes mellitus with other specified complications
C0342262|Type 2 diabetes mellitus with other specified complications
C0342262|Type 2 diabetes mellitus with other specified complication
C0342262|Diabetes mellitus, adult onset, with other specified manifestation (disorder)
C0342262|Diabetes mellitus, adult onset, with other specified manifestation
C3646651|pregnancy complications: chronic diabetes mellitus
C3646651|pregnancy complicated by chronic diabetes mellitus (diagnosis)
C3646651|pregnancy complications: diabetes mellitus chronic
C3646651|pregnancy complicated by chronic diabetes mellitus
C2874125|diabetes mellitus due to genetic defects of beta-cell function
C2874125|Diabetes mellitus due to genetic defect in beta cell function
C2874125|Diabetes mellitus due to genetic defect in beta cell function (disorder)
C2874124|diabetes mellitus due to genetic defects in insulin action
C2874124|Diabetes mellitus due to genetic defect in insulin action (disorder)
C2874124|Diabetes mellitus due to genetic defect in insulin action
C0392201|Blood glucose
C0392201|blood glucose tests (lab test)
C0392201|blood glucose tests
C0392201|Blood glucose measurement
C0392201|blood glucose level
C0392201|blood glucose measurement (lab test)
C0392201|Blood glucose (sugar) level
C0392201|Measurement of glucose in blood
C0392201|Blood Sugar
C0392201|Glucose Measurement, Blood
C0392201|Blood sugar level
C0392201|BS - Blood glucose level
C0392201|Glucose measurement, blood (procedure)
C0020456|Hyperglycemia
C0020456|Hyperglycemias
C0020456|Hyperglycaemia, unspecified
C0020456|Hyperglycemia, unspecified
C0020456|Hyperglycemia NOS
C0020456|[D]Hyperglycemia (context-dependent category)
C0020456|hyperglycemia (diagnosis)
C0020456|Hyperglycaemia
C0020456|Hyperglycemia [Disease/Finding]
C0020456|[X]Hyperglycaemia, unspecified
C0020456|[D]Hyperglycaemia
C0020456|[D]Hyperglycemia
C0020456|[D]Hyperglycaemia (situation)
C0020456|Hyperglycaemia (disorder)
C0020456|[D]Hyperglycemia (situation)
C0020456|[X]Hyperglycemia, unspecified (finding)
C0020456|[X]Hyperglycemia, unspecified
C0020456|Hyperglycemic disorder
C0020456|High blood sugar
C0020456|High Blood Glucose
C0020456|Blood Glucose, High
C0020456|Glucose, High Blood
C0020456|Hyperglycaemia NOS
C0020456|Elevated Blood Glucose
C0020456|Hyperglycaemic disorder
C0020456|Hyperglycemia (disorder)
C0020456|Hyperglycemic disorder (disorder)
C0020456|blood sugar; high
C0020456|blood; sugar, high
C0020456|high; blood sugar
C0020456|sugar; blood, high
C0020456|Hyperglycemia, NOS
C0020456|Hyperglycaemia, NOS
C0020456|[X]Hyperglycemia, unspecified (context-dependent category)
C0271687|diabetes mellitus due to structurally abnormal insulin (diagnosis)
C0271687|Diabetes mellitus due to structurally abnormal insulin
C0271687|Diabetes mellitus due to structurally abnormal insulin (disorder)
C0271687|Insulinopathy
C0271687|Diabetes mellitus due to abnormal insulin
C0271687|Insulinopathy, NOS
C0342274|diabetes mellitus associated with genetic syndrome (diagnosis)
C0342274|Diabetes mellitus associated with genetic syndrome
C0342274|Genetic syndromes of diabetes mellitus
C0342274|Diabetes mellitus associated with genetic syndrome (disorder)
C0342283|Hyperproinsulinemia
C0342283|Hyperproinsulinemia (diagnosis)
C0342283|diabetes mellitus hyperproinsulinemia
C0342283|Hyperproinsulinaemia
C0342283|Hyperproinsulinemia (disorder)
C1263962|Houssay syndrome
C1263962|Houssay's syndrome
C1263962|Houssay's syndrome (diagnosis)
C1263962|Houssay's syndrome (disorder)
C1960272|Latent autoimmune diabetes mellitus in adult (disorder)
C1960272|Latent autoimmune diabetes mellitus in adult
C1960272|Latent autoimmune diabetes mellitus in adult (LADA)
C1960272|diabetes mellitus latent autoimmune in adult
C1960272|Latent autoimmune diabetes mellitus in adult (diagnosis)
C1960626|Diabetes mellitus associated with cystic fibrosis
C1960626|Diabetes mellitus associated with cystic fibrosis (disorder)
C1960626|diabetes mellitus associated with cystic fibrosis (diagnosis)
C0342302|Brittle diabetes
C0342302|Brittle diabetes mellitus (disorder)
C0342302|Unstable diabetes mellitus
C0342302|Brittle diabetes mellitus (finding)
C0342302|Brittle diabetes mellitus
C0342302|Unstable diabetes
C0342302|Unstable diabetes mellitus (disorder)
C0342302|brittle diabetes mellitus (diagnosis)
C0342302|Diabetes brittle
C0342302|Labile diabetes
C0342302|brittle; diabetes
C0342302|diabetes; brittle
C0342302|diabetes; unstable
C0342302|unstable; diabetes
C0342302|Brittle diabetes (disorder)
C0342302|Unstable diabetes (disorder)
C0271701|DM due to insulin receptor ab
C0271701|Diabetes mellitus due to insulin receptor antibodies (disorder)
C0271701|Diabetes mellitus due to insulin receptor antibodies
C0271701|diabetes mellitus due to insulin receptor antibodies (diagnosis)
C0271701|Diabetes mellitus caused by insulin receptor antibodies
C0271701|DM caused by insulin receptor ab
C0271701|Diabetes mellitus caused by insulin receptor antibodies (disorder)
C1720029|Coma associated with diabetes mellitus (disorder)
C1720029|Coma associated with diabetes mellitus
C1720029|coma associated with diabetes mellitus (diagnosis)
C1857775|DIABETES MELLITUS, NEONATAL, WITH CONGENITAL HYPOTHYROIDISM
C1857775|NDH SYNDROME
C1835887|DIABETES MELLITUS, TRANSIENT NEONATAL, 2
C1835887|DIABETES MELLITUS, TRANSIENT NEONATAL, 2 (disorder)
C1835887|Diabetes mellitus, transient neonatal 2 (disorder)
C1835887|Diabetes mellitus, transient neonatal 2
C1835887|TNDM2
C1853564|DEND
C1853564|DEVELOPMENTAL DELAY, EPILEPSY, AND NEONATAL DIABETES
C1839028|MITOCHONDRIAL MYOPATHY WITH DIABETES
C1839028|Mitochondrial Myopathy, Lipid Type
C1864623|DIABETES MELLITUS, TRANSIENT NEONATAL, 3
C1864623|DIABETES MELLITUS, TRANSIENT NEONATAL, 3 (disorder)
C1864623|Diabetes mellitus, transient neonatal 3
C1864623|TNDM3
C1864623|Diabetes mellitus, transient neonatal 3 (disorder)
C0342278|DIABETES MELLITUS, INSULIN-RESISTANT, WITH ACANTHOSIS NIGRICANS
C0342278|Insulin Receptor Defect with Insulin-Resistant Diabetes Mellitus and Acanthosis Nigricans
C0342278|IRAN, Type A
C0342278|Diabetes Mellitus, Insulin-Resistant, with Acanthosis Nigricans, Type A
C0342278|INSULIN RECEPTOR, DEFECT IN, WITH INSULIN-RESISTANT DIABETES MELLITUS AND ACANTHOSIS NIGRICANS
C0342278|Hereditary benign acanthosis nigricans with insulin resistance
C0342278|Insulin-resistant acanthosis nigricans type A
C0342278|Hereditary benign acanthosis nigricans with insulin resistance (disorder)
C1864839|MODY7
C1864839|MATURITY-ONSET DIABETES OF THE YOUNG, TYPE 7
C1864839|MATURITY-ONSET DIABETES OF THE YOUNG, TYPE 7 (disorder)
C1864839|maturity-onset diabetes of the young - type 7
C1864839|maturity-onset diabetes of the young - type 7 (diagnosis)
C2748662|Mitchell-Riley Syndrome
C2748662|MTCHRS
C2748662|DIABETES, NEONATAL, WITH PANCREATIC HYPOPLASIA, INTESTINAL ATRESIA, AND GALLBLADDER APLASIA OR HYPOPLASIA
C0342281|MUSCULAR ATROPHY, ATAXIA, RETINITIS PIGMENTOSA, AND DIABETES MELLITUS
C0342281|Muscular atrophy, ataxia, retinitis pigmentosa, and diabetes mellitus (disorder)
C3711391|Tndm Type 1
C3711391|6q24-Related Transient Neonatal Diabetes Mellitus
C3711391|6q24-Tndm
C1857958|DIABETES MELLITUS, CONGENITAL AUTOIMMUNE
C1836780|PANCREATIC AND CEREBELLAR AGENESIS
C1836780|PACA
C1836780|Diabetes Mellitus, Permanent Neonatal, with Cerebellar Agenesis
C1859965|ALANINURIA WITH MICROCEPHALY, DWARFISM, ENAMEL HYPOPLASIA, AND DIABETES MELLITUS
C1859965|Stimmler Syndrome
C1859596|ATHEROSCLEROSIS, PREMATURE, WITH DEAFNESS, NEPHROPATHY, DIABETES MELLITUS, PHOTOMYOCLONUS, AND DEGENERATIVE NEUROLOGIC DISEASE
C1838782|WOLFRAM SYNDROME, MITOCHONDRIAL FORM
C1838782|DIDMOAD Syndrome, Mitochondrial Form
C1838782|Diabetes Insipidus And Mellitus With Optic Atrophy And Deafness, Mitochondrial Form
C1832386|DIABETES MELLITUS, TRANSIENT NEONATAL, 1
C1832386|TNDM1
C1832386|Diabetes mellitus, transient neonatal 1
C1832386|Diabetes mellitus, transient neonatal 1 (disorder)
C1832386|TNDM
C1832386|DMTN
C1838780|Pancreatic Hypoplasia, Congenital, with Diabetes Mellitus and Congenital Heart Disease
C2675066|LYMPHEDEMA-DISTICHIASIS SYNDROME WITH RENAL DISEASE AND DIABETES MELLITUS
C1833102|DIABETES MELLITUS, PERMANENT NEONATAL, WITH NEUROLOGIC FEATURES
C1833104|DIABETES MELLITUS, PERMANENT NEONATAL
C1833104|PNDM
C1833104|PDMI
C1833104|Diabetes Mellitus, Permanent, of Infancy
C1833104|Permanent diabetes mellitus of infancy
C1833104|Permanent neonatal diabetes mellitus (disorder)
C1833104|Permanent neonatal diabetes mellitus
C1832443|Martinez Frias syndrome
C1832443|Diabetes, Neonatal, with Pancreatic Hypoplasia, Intestinal Atresia, and Gallbladder Aplasia or Hypoplasia
C1832443|Martinez-Frias Syndrome
C1832443|Pancreatic Hypoplasia, Intestinal Atresia, and Gallbladder Aplasia or Hypoplasia, with or without Tracheoesophageal Fistula
C3828492|Pre-Gestational Diabetes
C3828492|Pregestational Diabetes
C3837964|diabetes mellitus with microvascular complications - MVCD3
C3837964|diabetes mellitus with microvascular complications - MVCD3 (diagnosis)
C3837962|diabetes mellitus with microvascular complications - MVCD5
C3837962|diabetes mellitus with microvascular complications - MVCD5 (diagnosis)
C3837966|diabetes mellitus with microvascular complications - MVCD1
C3837966|diabetes mellitus with microvascular complications - MVCD1 (diagnosis)
C3837963|diabetes mellitus with microvascular complications - MVCD4
C3837963|diabetes mellitus with microvascular complications - MVCD4 (diagnosis)
C3837965|diabetes mellitus with microvascular complications - MVCD2 (diagnosis)
C3837965|diabetes mellitus with microvascular complications - MVCD2
C3837960|diabetes mellitus with microvascular complications - MVCD7
C3837960|diabetes mellitus with microvascular complications - MVCD7 (diagnosis)
C3837961|diabetes mellitus with microvascular complications - MVCD6
C3837961|diabetes mellitus with microvascular complications - MVCD6 (diagnosis)
C3837959|diabetes mellitus with microvascular complications
C3837959|diabetes mellitus with microvascular complications (diagnosis)
C0021655|Insulin Resistance
C0021655|Resistance, Insulin
C0021655|Insulin Resistance [Disease/Finding]
C0021655|insulin resistance (diagnosis)
C0021655|Drug resistance to insulin
C0021655|Drug resistance to insulin (disorder)
C3839440|Diabetes mellitus in remission (disorder)
C3839440|Diabetes mellitus in remission
C3875503|Diabetes mellitus due to pancreatic injury
C3875503|Diabetes mellitus due to pancreatic injury (disorder)
C3896643|NODAT
C3896643|New Onset Diabetes After Transplant
C0342276|Maturity onset diabetes mellitus in young
C0342276|MODY
C0342276|MATURITY-ONSET DIABETES OF THE YOUNG
C0342276|Mason-Type Diabetes
C0342276|Diabetes, maturity-onset, of the young (MODY)
C0342276|Maturity onset diabetes in youth type 1
C0342276|Maturity-onset diabetes of the young (disorder)
C0342276|Maturity onset diabetes mellitus in young (disorder)
C0342276|MODY - Maturity onset diabetes in youth type 1
C0342276|Diabetes mellitus autosomal dominant (disorder)
C0342276|Diabetes mellitus autosomal dominant
C0342276|Autosomal dominant diabetes mellitus
C0342276|MODY - Maturity onset diabetes in youth type I
C0342276|Maturity onset diabetes in youth
C0342276|NIDDY
C0342276|maturity-onset diabetes of the young (diagnosis)
C0342276|Maturity Onset Diabetes of the Young
C0854110|Insulin-resistant diabetes mellitus
C0854110|Insulin resistant diabetes
C0854110|Insulin-resistant diabetes
C0854110|Insulin resistant diabetes mellitus
C0854110|insulin resistant diabetes (mellitus)
C0854110|Diabetes mellitus, insulin-resistant
C4039625|Gingivitis co-occurrent with diabetes mellitus
C4039625|Gingivitis co-occurrent with diabetes mellitus (disorder)
C0477821|Pre-existing diabetes mellitus, unspecified
C0477821|[X]Pre-existing diabetes mellitus, unspecified (disorder)
C0477821|[X]Pre-existing diabetes mellitus, unspecified
C0043207|Syndrome, Wolfram
C0043207|Wolfram Syndrome
C0043207|DIDMOAD
C0043207|WOLFRAM SYNDROME 1
C0043207|WFS1
C0043207|Diabetes mellitus and insipidus with optic atrophy and deafness
C0043207|Wolfram Syndrome [Disease/Finding]
C0043207|DIDMOAD Syndrome
C0043207|Diabetes Insipidus and Mellitus with Optic Atrophy and Deafness
C0043207|diabetes mellitus and insipidus with optic atrophy and deafness (diagnosis)
C0043207|Diabetes Insipidus, Diabetes Mellitus, Optic Atrophy, and Deafness
C0043207|DIDMOADUD
C0043207|Diabetes insipidus,diabetes mellitus, optic atrophy and deafness
C0043207|Diabetes insipidus, diabetes mellitus, optic atrophy and deafness
C0043207|DIDMOAD - Diabetes insipidus, diabetes mellitus, optic atrophy and deafness
C0043207|DIDMOAD - Diabetes insipidus,diabetes mellitus, optic atrophy and deafness
C0043207|WFS
C0043207|Marquardt-Loriaux syndrome
C0043207|Diabetes mellitus AND insipidus with optic atrophy AND deafness (disorder)
C0043207|Diabetes insipidus,diabetes mellitus, optic atrophy and deafness (disorder)
C1283034|Maternal diabetes mellitus
C1283034|Maternal diabetes mellitus (disorder)
C0271695|PINEAL HYPERPLASIA, INSULIN-RESISTANT DIABETES MELLITUS, AND SOMATIC ABNORMALITIES
C0271695|Pineal hyperplasia and diabetes mellitus syndrome
C0271695|Rabson-Mendenhall Syndrome
C0271695|Rabson Mendenhall Syndrome
C0271695|Syndrome, Mendenhall
C0271695|Syndrome, Rabson-Mendenhall
C0271695|Pineal hyperplasia AND diabetes mellitus syndrome (diagnosis)
C0271695|diabetes mellitus associated with genetic syndrome pineal hyperplasia
C0271695|MENDENHALL SYNDROME
C0271695|Pineal hyperplasia, insulin-resistant diabetes mellitus and somatic abnormalities
C0271695|Pineal hyperplasia AND diabetes mellitus syndrome (disorder)
C0271695|Pineal hyperplasia, insulin-resistant diabetes mellitus and somatic abnormalities (disorder)
C0271670|Pregestational diabetes mellitus AND/OR impaired glucose tolerance, modified White class R (disorder)
C0271670|Pregestational diabetes mellitus AND/OR impaired glucose tolerance, modified White class R
C0271670|Pregestational diabetes mellitus or impaired glucose tolerance, modified White class R
C0854359|Insulin autoimmune syndrome
C0854359|autoimmune endocrine disease insulin syndrome
C0854359|autoimmune insulin syndrome
C0854359|autoimmune insulin syndrome (diagnosis)
C0854359|Insulin autoimmune syndrome (disorder)
C0011859|Diabetes Mellitus, Lipoatrophic
C0011859|Lipoatrophic Diabetes Mellitus
C0011859|Lipoatrophic Diabetes
C0011859|Diabetes Mellitus, Lipoatrophic [Disease/Finding]
C0011859|Diabetes, Lipoatrophic
C0011859|Lipoatrophic Diabete
C0011859|Diabete, Lipoatrophic
C0011859|Lipoatrophic diabetes (disorder)
C0011859|Lipodystrophic diabetes
C0011859|Lipoatrophic diabetes, NOS
C0011859|Lipodystrophic diabetes, NOS
C0154183|Diabetes with other specified manifestations
C0154172|Type I diabetes mellitus with hyperosmolar coma
C0235397|Diabetes mellitus precipitated
C0235398|Diabetes mellitus aggravated
C0235398|Diabetes mellitus exacerbated
C0235399|Diabetes mellitus reactivated
C0241861|diabetes; stable
C0241861|stable; diabetes
C0342297|Diabetes mellitus, adult onset, with hyperosmolar coma (disorder)
C0342297|Type 2 diabetes mellitus with hyperosmolar coma
C0342297|Type 2 diabetes mellitus with hyperosmolar coma (disorder)
C0342297|Diabetes mellitus, adult onset, with hyperosmolar coma
C0342297|Type II diabetes mellitus with hyperosmolar coma
C0494293|Other specified diabetes mellitus without complications
C0342269|Steroid-induced diabetes
C0342269|Steroid-induced diabetes (disorder)
C0342269|Diabetes steroid-induced
C0546950|Type II diabetes mellitus without mention of complication
C0011884|Diabetic Retinopathies
C0011884|Diabetic Retinopathy
C0011884|Retinopathies, Diabetic
C0011884|Retinopathy, Diabetic
C0011884|DR - Diabetic retinopathy
C0011884|DR
C0011884|Diabetic Retinopathy [Disease/Finding]
C0011884|Retinopathy;diabetic
C0011884|Retinopathy - diabetic
C0011884|Retinal abnormality - diabetes-related (disorder)
C0011884|Retinal abnormality - diabetes-related
C0011884|Diabetic retinopathy NOS (disorder)
C0011884|Diabetic retinopathy (disorder)
C0011884|Diabetic retinopathy NOS
C0011884|diabetes with diabetic retinopathy
C0011884|diabetes with diabetic retinopathy (diagnosis)
C0011884|diabetes mellitus with diabetic retinopathy
C0011884|Retinopathy diabetic
C0011884|Diabetic retinopathy, NOS
C0865162|Diabetes mellitus without mention of complication or manifestation
