C1274583|Non-professional tattoo
C1274583|Amateur tattoo
C1274583|tattoo dirty
C1274583|tattoo infected
