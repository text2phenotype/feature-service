C2367818|hepatitis C treatment prescribed
C2367821|peginterferon and ribavirin therapy considered for hepatitis C
C2367822|peginterferon and ribavirin therapy prescribed for hepatitis C
C2750389|HEPATITIS C VIRUS INFECTION, RESPONSE TO THERAPY OF
C2750389|Previous HCV Treatment
C2750389|Previously treated for HCV
C2750389|Previous treatment for HCV
C2750389|Previous HCV treatment
C2367819|antiviral hepatitis C treatment being received (treatment)
C2367819|antiviral hepatitis C treatment being received
C2367820|antiviral hepatitis C treatment not being received (treatment)
C2367820|antiviral hepatitis C treatment not being received
C2367821|peginterferon and ribavirin therapy considered for hepatitis C (treatment)
C2367821|peginterferon and ribavirin therapy considered for hepatitis C
C2367822|peginterferon and ribavirin therapy prescribed for hepatitis C (treatment)
C2367822|peginterferon and ribavirin therapy prescribed for hepatitis C
