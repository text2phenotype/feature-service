C3871344|Current or former injection drug user (even once)
C3871344|Current or former injection drug user
C3871344|Current or former IV drug user
C3871344|Current or former IV user
C3871344|Current IV user
C3871344|Former IV user
C3871344|Former IV drug user
C3871344|History of injection drug use
C3871344|History of IV drug use
C3871344|History of IV use
C3871344|Hx injec drug use
C3871344|Hx IV use
C3871344|History IV use
C3871344|Uses IV needles
C3871344|IV drug user
C3871344|History of injection drug use
C3871344|Hx injec drug use
