C3160090|HCV NS3/4A Protease Inhibitors [MoA]
C1738934|boceprevir 
C1876229|telaprevir
C2605855|simeprevir
C3154649|boceprevir 200 MG Oral Capsule
C3154711|telaprevir 375 MG Oral Tablet
C0697341|Inderal 10 MG Oral Tablet
C0591636|Inderal
C3226084|Inderal Pill
C3226083|Inderal Oral Product
C2710361|Propranolol Hydrochloride 120 MG [Inderal]
C2710374|Propranolol Hydrochloride 160 MG [Inderal]
C2710406|Propranolol Hydrochloride 60 MG [Inderal]
C2710422|Propranolol Hydrochloride 80 MG [Inderal]
C1577533|Propranolol Extended Release Oral Capsule [Inderal]
C0697868|24 HR Propranolol Hydrochloride 160 MG Extended Release Oral Capsule [Inderal]
C0697871|24 HR Propranolol Hydrochloride 80 MG Extended Release Oral Capsule [Inderal]
C0709220|24 HR Propranolol Hydrochloride 60 MG Extended Release Oral Capsule [Inderal]
C0709222|24 HR Propranolol Hydrochloride 120 MG Extended Release Oral Capsule [Inderal]
C0022957|Lactulose
C0994966|Lactulose Oral Solution [Enulose]
C1134051|Lactulose 667 MG/ML
C1178770|Lactulose 670 MG/ML
C1252332|Lactulose Oral Solution
C1589308|Lactulose Oral Solution [Constulose]
C1589310|Lactulose Oral Solution [Generlac]
C3216530|Lactulose Oral Liquid Product
C3216531|Lactulose Oral Product
C4306942|Lactulose 10000 MG [Kristalose]
C4306943|Lactulose 20000 MG [Kristalose]
C4307200|Lactulose 10000 MG
C4307201|Lactulose 20000 MG
C4307247|Lactulose Powder for Oral Solution
C4307286|Lactulose Oral Powder Product
C1589307|Lactulose 667 MG/ML [Constulose]
C1589309|Lactulose 667 MG/ML [Generlac]
C1600254|Lactulose 667 MG/ML [Enulose]
C4307030|Lactulose Powder for Oral Solution [Kristalose]
C0353982|Lactulose 670 MG/ML Oral Solution
C0708296|Lactulose 667 MG/ML Oral Solution [Enulose]
C0978083|Lactulose 10000 MG Powder for Oral Solution
C1298316|Lactulose 667 MG/ML Oral Solution
C1586235|Lactulose 667 MG/ML Oral Solution [Constulose]
C1586236|Lactulose 667 MG/ML Oral Solution [Generlac]
C1613498|Lactulose 20000 MG Powder for Oral Solution [Kristalose] 
C1620382|Lactulose 10000 MG Powder for Oral Solution [Kristalose] 
C1737835|Lactulose 20000 MG Powder for Oral Solution
C0043031|Warfarin
C3154650|Victrelis
C3154650|vicrtelis
C1738934|N-(3-amino-1-(cyclobutylmethyl)-2,3-dioxopropyl)-3-(2-((((1,1-dimethylethyl)amino)carbonyl)amino)-3,3-dimethyl-1-oxobutyl)-6,6-dimethyl-3-azabicyclo(3.1.0)hexan-2-carboxamide
C1738934|boceprevir
C1738934|antivirals boceprevir
C1738934|antivirals boceprevir (medication)
C1738934|Boceprevir (substance)
C1738934|Boceprevir (product)
C1738934|3-Azabicyclo(3.1.0)hexane-2-carboxamide, N-(3-amino-1-(cyclobutylmethyl)-2,3-dioxopropyl)-3-((2S)-2-((((1,1- dimethylethyl)amino)carbonyl)amino)-3,3-dimethyl-1-oxobutyl)-6,6- dimethyl-, (1R,2S,5S)-
C3154649|Boceprevir Cap 200 MG
C3154649|BOCEPREVIR 200MG CAP
C3154649|boceprevir 200 mg oral capsule
C3154649|BOCEPREVIR 200MG CAP [VA Product]
C3154649|Boceprevir 200mg Oral capsule
C3154649|Boceprevir 200mg capsule (product)
C3154649|Boceprevir 200mg capsule
C1741239|Sch-503034
C1741239|Sch 503034
C1741239|Sch503034
C3896865|EBP 520
C3154701|Incivek
C1876229|telaprevir
C1876229|antiviral telaprevir
C1876229|antiviral telaprevir (medication)
C1876229|Telaprevir (substance)
C1876229|Telaprevir (product)
C3281323|VRT-111950
C3281324|MP-424
C3281325|LY-570310
C1956374|VX-950
C1956374|VX 950
C1956374|VX950 cpd
C3154711|telaprevir 375 MG Oral Tablet
C3154711|Telaprevir Tab 375 MG
C3154711|TELAPREVIR 375MG TAB
C3154711|TELAPREVIR 375MG TAB,28 [VA Product]
C3154711|TELAPREVIR 375MG TAB,28
C3154711|TELAPREVIR 375MG TAB [VA Product]
C3154711|Telaprevir 375mg Oral tablet
C3154711|TELAPREVIR 375MG TAB,UD
C3154711|TELAPREVIR 375MG UD TAB
C3154711|TELAPREVIR 375MG TAB,UD [VA Product]
C3154711|Telaprevir 375mg tablet
C3154711|Telaprevir 375mg tablet (product)
C2605856|435350, TMC
C2605856|TMC435350
C2605856|TMC-435350
C2605856|TMC 435350
C2745868|435, TMC
C2745868|TMC435
C2745868|TMC-435
C2745868|TMC 435
C3696409|Olysio
C2605855|simeprevir
C2605855|simeprevir (medication)
C2605855|antiviral simeprevir
C2605855|Simeprevir (substance)
C2605855|N-(17-(2-(4-isopropylthiazole-2-yl)-7-methoxy-8-methylquinolin-4-yloxy)-13-methyl-2,14-dioxo-3,13-diazatricyclo(13.3.0.04,6)octadec-7-ene-4-carbonyl)(cyclopropyl)sulfonamide
C2605855|Simeprevir [Chemical/Ingredient]
C2605855|Simeprevir (product)
C3696072|simeprevir sodium
C3696072|simeprevir (as sodium)
C3696748|simeprevir Oral Product
C3696748|Oral form simeprevir (product)
C3696748|Oral form simeprevir
C4075528|Simeprevir + sofosbuvir (product)
C4075528|Simeprevir + sofosbuvir
C3154653|BOCEPREVIR 200 mg ORAL CAPSULE [VICTRELIS]
C3154653|Victrelis 200 MG Oral Capsule
C3154653|VICTRELIS 200mg Capsule
C3154653|Victrelis, 200 mg oral capsule
C3154713|telaprevir 375 MG Oral Tablet [Incivek]
C3154713|Incivek 375 MG Oral Tablet
C3154713|INCIVEK 375mg Tablet
C3154713|Incivek, 375 mg oral tablet
C3154713|INCIVEK 375 MG Oral Tablet, Twice Daily
C0697341|Inderal 10mg Tablet
C0697341|Inderal, 10 mg oral tablet
C0697341|Inderal 10 MG Oral Tablet
C0697341|Propranolol Hydrochloride 10 MG Oral Tablet [Inderal]
C0282321|Hydrochloride, Propranolol
C0282321|Propranolol Hydrochloride
C0282321|2-Propanol-1-[(1-methylethyl)amino]-3-(1-naphthalenyloxy) Hydrochloride
C0282321|Propranolol hydrochloride product
C0282321|propranolol hydrochloride (medication)
C0282321|Propranolol Hydrochloride [Chemical/Ingredient]
C0282321|Propranolol hydrochloride [2]
C0282321|Propranolol hydrochloride [2] (product)
C0282321|Propranolol hydrochloride (product)
C0282321|Propranolol hydrochloride (substance)
C0282321|Propranolol hydrochloride [2] (substance)
C0282321|Propranolol hydrochloride product (product)
C0282321|Propranolol hydrochloride product (substance)
C0591636|Inderal
C0697332|Inderal 160 MG Oral Tablet
C0697332|Propranolol Hydrochloride 160 MG Oral Tablet [Inderal]
C1271144|Inderal 80 MG Oral Capsule
C1271144|Propranolol Hydrochloride 80 MG Oral Capsule [Inderal]
C1271144|Inderal 80mg capsule
C1271144|Inderal 80mg capsule (product)
C0709222|propranolol hydrochloride 120 MILLIGRAM In 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [Inderal LA]
C0709222|Inderal LA 120mg Extended-Release Capsule
C0709222|Inderal LA, 120 mg oral capsule, extended release
C0709222|Propranolol Hydrochloride 120 MG Oral Capsule, Extended Release [INDERAL LA]
C0709222|PROPRANOLOL HYDROCHLORIDE 120 mg ORAL CAPSULE, EXTENDED RELEASE [INDERAL XL]
C0709222|Inderal XL, 120 mg oral capsule, extended release
C0709222|Inderal XL 120mg Extended-Release Capsule
C0709222|24 HR Propranolol Hydrochloride 120 MG Extended Release Oral Capsule [Inderal]
C0709222|Inderal LA 120 MG 24HR Extended Release Oral Capsule
C0709222|Inderal XL 120 MG 24 HR Extended Release Oral Capsule
C2710362|Inderal 120 MG Extended Release Oral Capsule
C2710362|Propranolol Hydrochloride 120 MG Extended Release Oral Capsule [Inderal]
C0697868|propranolol hydrochloride 160 MILLIGRAM In 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [Inderal LA]
C0697868|Inderal LA 160mg Extended-Release Capsule
C0697868|Inderal LA, 160 mg oral capsule, extended release
C0697868|Propranolol Hydrochloride 160 MG Oral Capsule, Extended Release [INDERAL LA]
C0697868|Inderal LA 160 MG 24 HR Extended Release Oral Capsule
C0697868|Inderal LA 160 MG 24HR Extended Release Oral Capsule
C0697868|24 HR Inderal LA 160 MG Extended Release Oral Capsule
C0697868|24 HR Propranolol Hydrochloride 160 MG Extended Release Oral Capsule [Inderal]
C2710375|Propranolol Hydrochloride 160 MG Extended Release Oral Capsule [Inderal]
C2710375|Inderal 160 MG Extended Release Oral Capsule
C0709233|Inderal 20mg Tablet
C0709233|Inderal, 20 mg oral tablet
C0709233|Propranolol Hydrochloride 20 MG Oral Tablet [Inderal]
C0709233|Inderal 20 MG Oral Tablet
C0697330|Inderal 40mg Tablet
C0697330|Inderal, 40 mg oral tablet
C0697330|Propranolol Hydrochloride 40 MG Oral Tablet [Inderal]
C0697330|Inderal 40 MG Oral Tablet
C0709220|propranolol hydrochloride 60 MILLIGRAM In 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [Inderal LA]
C0709220|Inderal LA 60mg Extended-Release Capsule
C0709220|Inderal LA, 60 mg oral capsule, extended release
C0709220|Propranolol Hydrochloride 60 MG Oral Capsule, Extended Release [INDERAL LA]
C0709220|Inderal LA 60 MG 24 HR Extended Release Oral Capsule
C0709220|24 HR Propranolol Hydrochloride 60 MG Extended Release Oral Capsule [Inderal]
C0709220|24 HR Inderal LA 60 MG Extended Release Oral Capsule
C0709220|Inderal LA 60 MG 24HR Extended Release Oral Capsule
C2710407|Inderal 60 MG Extended Release Oral Capsule
C2710407|Propranolol Hydrochloride 60 MG Extended Release Oral Capsule [Inderal]
C0709234|Inderal 60mg Tablet
C0709234|Inderal, 60 mg oral tablet
C0709234|Inderal 60 MG Oral Tablet
C0709234|Propranolol Hydrochloride 60 MG Oral Tablet [Inderal]
C0697871|propranolol hydrochloride 80 MILLIGRAM In 1 CAPSULE ORAL CAPSULE, EXTENDED RELEASE [Inderal LA]
C0697871|Inderal LA 80mg Extended-Release Capsule
C0697871|Inderal LA, 80 mg oral capsule, extended release
C0697871|Propranolol Hydrochloride 80 MG Oral Capsule, Extended Release [INDERAL LA]
C0697871|PROPRANOLOL HYDROCHLORIDE 80 mg ORAL CAPSULE, EXTENDED RELEASE [INDERAL XL]
C0697871|Inderal XL 80mg Extended-Release Capsule
C0697871|Inderal XL, 80 mg oral capsule, extended release
C0697871|24 HR Propranolol Hydrochloride 80 MG Extended Release Oral Capsule [Inderal]
C0697871|Inderal XL 80 MG 24 HR Extended Release Oral Capsule
C0697871|Inderal LA 80 MG 24HR Extended Release Oral Capsule
C2710423|Inderal 80 MG Extended Release Oral Capsule
C2710423|Propranolol Hydrochloride 80 MG Extended Release Oral Capsule [Inderal]
C0697347|Inderal 80mg Tablet
C0697347|Inderal, 80 mg oral tablet
C0697347|Propranolol Hydrochloride 80 MG Oral Tablet [Inderal]
C0697347|Inderal 80 MG Oral Tablet
C1306227|Propranolol Oral Capsule [Inderal]
C1577533|Propranolol Extended Release Oral Capsule [Inderal]
C0306453|Propranolol Oral Tablet [Inderal]
C0059478|epsilon-N-1-(1-deoxylactulosyl)lysine
C0701236|Normase
C0701237|Amivalex
C0719221|Cephulac
C0719324|Cholac
C0719340|Chronulac
C0719488|Constilac
C0719489|Constulose
C0720231|Enulose
C0720316|Evalose
C0720632|Generlac
C0720849|Heptalac
C0721265|Kristalose
C0116371|epsilon-(deoxylactulose)lysine
C0125215|lactose-lysine
C0125227|lactulose-lysine
C0284752|lactuloselysine
C0022957|Lactulose
C0022957|D-Fructose, 4-O-beta-D-galactopyranosyl-
C0022957|lactulose (medication)
C0022957|laxatives lactulose
C0022957|4-O-beta-D-Galactopyranosyl-D-fructofuranose
C0022957|Lactulose [Chemical/Ingredient]
C0022957|Lactulose product
C0022957|Lactulose (product)
C0022957|Lactulose (substance)
C1737835|Lactulose 20g Powder for Oral sol/PWD [Constipation]
C1737835|LACTULOSE 20GM/PKT PWDR
C1737835|Lactulose Oral Crystal Packet 20 GM
C1737835|LACTULOSE 20GM/PKT PWDR [VA Product]
C1737835|Lactulose 167 MG/ML Oral Solution
C1737835|lactulose 20 GM per 4 OZ. Powder for Oral Solution
C1737835|lactulose 20 g oral powder for reconstitution
C1298316|Lactulose 667 MG/ML Oral Solution
C1298316|Lactulose (Encephalopathy) Solution 10 GM/15ML
C1298316|Lactulose Solution 10 GM/15ML
C1298316|Lactulose 10g/15mL Oral solution [Encephalopathy]
C1298316|Lactulose 10g/15mL Oral solution [Constipation]
C1298316|LACTULOSE 10GM/15ML SYRUP
C1298316|Lactulose 10 GM/15 ML Solution
C1298316|LACTULOSE 10 g in 15 mL ORAL SOLUTION
C1298316|lactulose 10 GM per 15 ML Oral Solution
C1298316|LACTULOSE 10 g in 15 mL ORAL SOLUTION [Lactulose]
C1298316|lactulose 20 GM per 30 ML Oral Solution
C1298316|LACTULOSE 10GM/15ML SYRUP [VA Product]
C1298316|LACTULOSE 20 g in 30 mL ORAL SOLUTION
C1298316|LACTULOSE 10 g in 15 mL RECTAL SOLUTION
C1298316|Lactulose, 10 g/15 mL oral and rectal liquid
C1298316|lactulose 10 g/15 mL oral and rectal liquid
C1298316|LACTULOSE 10GM/15ML ORAL SOLN
C1298316|LACTULOSE 10GM/15ML SOLN,ORAL
C1298316|LACTULOSE 10GM/15ML SOLN,ORAL [VA Product]
C1298316|Lactulose 10g/15 mL solution (product)
C1298316|Lactulose 10g/15 mL solution
C1298316|Acilac 10g/15ml Solution
C1298316|Lactulose 10g/15mL solution (product)
C1298316|Lactulose 10g/15mL solution
C1298316|Lactulose 10g/15mL syrup (product)
C1298316|Lactulose 10g/15mL syrup
C1298316|Lactulose 10 GM/15 ML Oral Solution
C1298316|Lactulose 10 GM/15 ML Oral Syrup
C1298316|Lactulose, 10 g/15 mL oral syrup
C1298316|lactulose 10 g/15 mL oral syrup
C3216531|Lactulose Oral Product
C3216531|Oral form lactulose (product)
C3216531|Oral form lactulose
C0353982|Lactulose 670 MG/ML Oral Solution
C0353982|lactulose 3.35 GM per 5 ML Oral Solution
C0353982|Lactulose 3.35g/5mL oral solution
C0353982|Lactulose 3.35g/5mL oral solution (product)
C0353982|Lactulose 3.35g/5mL oral solution (substance)
C0591418|Duphalac
C1589304|Catulac
C1589311|RO-Lactulose
C0605673|Cholan-24-oic acid, 3,7,12-trioxo-, (5beta)-, mixt. with (3(S)-endo)-8-(2-(1,1'-biphenyl)-4-yl-2-oxoethyl)-3-(3-hydroxy-1-oxo-2-phenylpropoxy)-8-methyl-8-azoniabicyclo(3.2.1)octane bromide, 4-O-beta-D-galactopyranosyl-D-fructose and pancreatin
C0605673|FZ 560
C0605673|FZ-560
C0708296|lactulose 10 GRAM In 15 MILLILITER ORAL LIQUID [Enulose]
C0708296|lactulose 10 GRAM In 15 MILLILITER RECTAL LIQUID [Enulose]
C0708296|Lactulose 667 MG/ML Oral Solution [Enulose]
C0708296|Enulose 667 MG/ML Oral Solution
C0708296|Enulose 10 GM per 15 ML Syrup
C0708296|Lactulose 10 GM/15 ML Oral Solution [ENULOSE]
C0708296|Lactulose 10 GM/15 ML Oral Syrup [ENULOSE]
C0708296|LACTULOSE 10 g in 15 mL RECTAL SOLUTION [Enulose]
C0708296|LACTULOSE 10 g in 15 mL ORAL SOLUTION [Enulose]
C0708296|Enulose, 10 g/15 mL oral and rectal liquid
C0708296|Enulose 10g/15ml Solution
C0994966|Lactulose Oral Solution [Enulose]
C0994966|LACTULOSE 10GM/15ML SYRUP
C0994966|ENULOSE SYRUP
C0994966|ENULOSE SYRUP [VA Product]
C1589305|Lactulose 667 MG/ML [Catulac]
C1589307|Lactulose 667 MG/ML [Constulose]
C1589309|Lactulose 667 MG/ML [Generlac]
C1589312|Lactulose 667 MG/ML [RO-Lactulose]
C1600249|Lactulose 667 MG/ML [Cephulac]
C1600250|Lactulose 667 MG/ML [Cholac]
C1600251|Lactulose 667 MG/ML [Chronulac]
C1600252|Lactulose 667 MG/ML [Constilac]
C1600253|Lactulose 667 MG/ML [Duphalac]
C1600254|Lactulose 667 MG/ML [Enulose]
C1600255|Lactulose 667 MG/ML [Evalose]
C1600256|Lactulose 667 MG/ML [Heptalac]
C0978083|Lactulose 10g Powder for Oral sol/PWD [Constipation]
C0978083|LACTULOSE 10GM/PKT PWDR
C0978083|Lactulose Oral Crystal Packet 10 GM
C0978083|LACTULOSE 10GM/PKT PWDR [VA Product]
C0978083|lactulose 10 GM per 4 OZ. Powder for Oral Solution
C0978083|Lactulose 83.3 MG/ML Oral Solution
C0978083|lactulose 10 g oral powder for reconstitution
C1352027|Lactulose 660 MG/ML Oral Solution
C1238377|Lactulose Oral Solution [Kristalose]
C1589308|Lactulose Oral Solution [Constulose]
C1589310|Lactulose Oral Solution [Generlac]
C1589313|Lactulose Oral Solution [RO-Lactulose]
C1355127|Lactulose 606 MG/ML Oral Solution
C1355126|Lactulose 650 MG/ML Oral Solution
C1355125|Lactulose 666 MG/ML Oral Solution
C1589306|Lactulose Oral Solution [Catulac]
C2240661|Lactulose Oral Solution [Cephulac]
C1239130|Lactulose Oral Solution [Cholac]
C2240662|Lactulose Oral Solution [Chronulac]
C1239069|Lactulose Oral Solution [Constilac]
C2240663|Lactulose Oral Solution [Duphalac]
C1239128|Lactulose Oral Solution [Evalose]
C1239126|Lactulose Oral Solution [Heptalac]
C1586235|Lactulose 667 MG/ML Oral Solution [Constulose]
C1586235|Constulose 667 MG/ML Oral Solution
C1586235|Constulose 10 GM per 15 ML Syrup
C1586235|Lactulose 10 GM/15 ML Oral Solution [CONSTULOSE]
C1586235|Lactulose 10 GM/15 ML Oral Syrup [CONSTULOSE]
C1586235|LACTULOSE 10 g in 15 mL ORAL SOLUTION [Constulose]
C1586235|Constulose 10g/15ml Solution
C1586235|Constulose, 10 g/15 mL oral syrup
C1586236|Generlac 667 MG/ML Oral Solution
C1586236|Lactulose 667 MG/ML Oral Solution [Generlac]
C1586236|Lactulose 10 GM/15 ML Oral Solution [GENERLAC]
C1586236|Lactulose 10 g in 15 mL ORAL SOLUTION [Generlac]
C1586236|Generlac 10 GM per 15 ML Oral Solution
C1586236|Generlac, 10 g/15 mL oral and rectal liquid
C1586236|Generlac 10g/15ml Solution
C3221021|Cephulac Oral Liquid Product
C3221216|Duphalac Oral Liquid Product
C3221248|Enulose Oral Liquid Product
C3222920|Constilac Oral Liquid Product
C3222922|Constulose Oral Liquid Product
C3223259|Heptalac Oral Liquid Product
C3223942|Generlac Oral Liquid Product
C3224342|Cholac Oral Liquid Product
C3224366|Chronulac Oral Liquid Product
C3225241|Evalose Oral Liquid Product
C3228268|Kristalose Oral Liquid Product
C3230348|Catulac Oral Liquid Product
C3231581|RO-Lactulose Oral Liquid Product
C1252332|Lactulose Oral Solution
C0787976|Lactulose 0.4 MG/MG Oral Gel
C1359419|Lactulose 2500 MG Oral Tablet
C1363276|Lactulose 2865 MG Chewable Tablet
C3221022|Cephulac Oral Product
C3221217|Duphalac Oral Product
C3221249|Enulose Oral Product
C3222921|Constilac Oral Product
C3222923|Constulose Oral Product
C3223260|Heptalac Oral Product
C3223943|Generlac Oral Product
C3224343|Cholac Oral Product
C3224367|Chronulac Oral Product
C3225242|Evalose Oral Product
C3228269|Kristalose Oral Product
C3230349|Catulac Oral Product
C3231582|RO-Lactulose Oral Product
C1252272|Lactulose Oral Gel
C1370590|Lactulose Oral Tablet
C1370592|Lactulose Chewable Tablet
C1620382|Lactulose 10 GM/PACKET Oral Powder for Suspension [KRISTALOSE]
C1620382|Kristalose 83.3 MG/ML Oral Solution
C1620382|Kristalose 10 GM per 4 OZ. Powder for Oral Solution
C1620382|Lactulose 83.3 MG/ML Oral Solution [Kristalose]
C1620382|lactulose 10 g in 10 g ORAL POWDER, FOR SOLUTION [Kristalose]
C1620382|Kristalose 10g Powder for Solution
C1620382|Kristalose, 10 g oral powder for reconstitution
C0708295|Lactulose 667 MG/ML Oral Solution [Duphalac]
C0708295|Duphalac 667 MG/ML Oral Solution
C0708295|Duphalac 10 GM per 15 ML Syrup
C0708295|Lactulose 10 GM/15 ML Oral Syrup [DUPHALAC]
C0708295|Duphalac, 10 g/15 mL oral syrup
C1695496|Lactulose 667 MG/ML Oral Solution [RO-Lactulose]
C1695496|RO-Lactulose 667 MG/ML Oral Solution
C1586234|Lactulose 667 MG/ML Oral Solution [Catulac]
C1586234|Catulac 667 MG/ML Oral Solution
C0708290|Cephulac 10g/15ml Solution
C0708290|Cephulac 667 MG/ML Oral Solution
C0708290|Lactulose 667 MG/ML Oral Solution [Cephulac]
C0708290|Cephulac 10 GM per 15 ML Syrup
C0708290|Lactulose 10 GM/15 ML Oral Syrup [CEPHULAC]
C0708290|Cephulac, 10 g/15 mL oral syrup
C0708291|Cholac 667 MG/ML Oral Solution
C0708291|Lactulose 667 MG/ML Oral Solution [Cholac]
C0708291|Cholac 10 GM per 15 ML Syrup
C0708291|Lactulose 10 GM/15 ML Oral Syrup [CHOLAC]
C0708291|Cholac 10g/15ml Solution
C0708291|Cholac, 10 g/15 mL oral syrup
C0708292|Chronulac 10g/15ml Solution
C0708292|Lactulose 667 MG/ML Oral Solution [Chronulac]
C0708292|Chronulac 667 MG/ML Oral Solution
C0708292|Chronulac 10 GM per 15 ML Syrup
C0708292|Lactulose 10 GM/15 ML Oral Syrup [CHRONULAC]
C0708292|Chronulac, 10 g/15 mL oral syrup
C0708293|Lactulose 667 MG/ML Oral Solution [Constilac]
C0708293|Constilac 667 MG/ML Oral Solution
C0708293|Constilac 10 GM per 15 ML Syrup
C0708293|Lactulose 10 GM/15 ML Oral Syrup [CONSTILAC]
C0708293|Constilac 10g/15ml Solution
C0708293|Constilac, 10 g/15 mL oral syrup
C0708297|Evalose 667 MG/ML Oral Solution
C0708297|Lactulose 667 MG/ML Oral Solution [Evalose]
C0708297|Evalose 10 GM per 15 ML Syrup
C0708297|Lactulose 10 GM/15 ML Oral Syrup [EVALOSE]
C0708297|Evalose, 10 g/15 mL oral syrup
C0708299|Lactulose 667 MG/ML Oral Solution [Heptalac]
C0708299|Heptalac 667 MG/ML Oral Solution
C0708299|Lactulose 10 GM/15 ML Oral Solution [HEPTALAC]
C0708299|Lactulose 10 GM/15 ML Oral Syrup [HEPTALAC]
C0708299|Heptalac, 10 g/15 mL oral syrup
C1613498|Lactulose 20 GM/PACKET Oral Powder for Suspension [KRISTALOSE]
C1613498|Lactulose 167 MG/ML Oral Solution [Kristalose]
C1613498|Kristalose 20 GM per 4 OZ. Powder for Oral Solution
C1613498|Kristalose 167 MG/ML Oral Solution
C1613498|lactulose 20 g in 20 g ORAL POWDER, FOR SOLUTION [Kristalose]
C1613498|Kristalose 20g Powder for Solution
C1613498|Kristalose, 20 g oral powder for reconstitution
C0981135|Warfarin Sodium 1mg Oral tablet
C0981135|Warfarin Sodium, 1 mg oral tablet
C0981135|warfarin 1 mg oral tablet
C0981135|WARFARIN (COUMADIN) NA 1MG TAB UD
C0981135|WARFARIN (COUMADIN) NA 1MG TAB
C0981135|Warfarin Sodium Tab 1 MG
C0981135|Warfarin Sodium 1 MG Oral Tablet
C0981135|WARFARIN NA (GOLDEN STATE) 1MG TAB
C0981135|WARFARIN NA 1MG TAB
C0981135|WARFARIN NA (GOLDEN STATE) 1MG TAB [VA Product]
C0981135|WARFARIN NA 1MG TAB,UD
C0981135|WARFARIN NA 1MG TAB,UD [VA Product]
C0981135|WARFARIN NA 1MG TAB [VA Product]
C0981135|WARFARIN SODIUM 1 mg ORAL TABLET [Warfarin Sodium]
C0981135|WARFARIN NA (EXELAN) 1MG TAB
C0981135|WARFARIN NA (EXELAN) 1MG TAB [VA Product]
C0981135|Warfarin sodium 1mg tablet
C0981135|Warfarin sodium 1mg tablet (product)
C0981135|Warfarin sodium 1mg tablet (substance)
C0690746|Warfarin Sodium 4mg Oral tablet
C0690746|WARFARIN NA 4MG TAB,UD
C0690746|Warfarin Sodium, 4 mg oral tablet
C0690746|warfarin 4 mg oral tablet
C0690746|WARFARIN (COUMADIN) NA 4MG TAB UD
C0690746|WARFARIN (COUMADIN) NA 4MG TAB
C0690746|Warfarin Sodium Tab 4 MG
C0690746|Warfarin Sodium 4 MG Oral Tablet
C0690746|WARFARIN NA (GOLDEN STATE) 4MG TAB
C0690746|WARFARIN NA 4MG TAB [VA Product]
C0690746|WARFARIN NA (GOLDEN STATE) 4MG TAB [VA Product]
C0690746|WARFARIN NA 4MG TAB
C0690746|WARFARIN NA 4MG TAB,UD [VA Product]
C0690746|Warfarin Sodium 4 mg ORAL TABLET [Warfarin Sodium]
C0690746|WARFARIN NA (EXELAN) 4MG TAB
C0690746|WARFARIN NA (EXELAN) 4MG TAB [VA Product]
C0690746|Warfarin sodium 4mg tablet (product)
C0690746|Warfarin sodium 4mg tablet
C0981139|Warfarin 2mg/mL powder for injection solution (product)
C0981139|Warfarin 2mg/mL powder for injection solution
C0981139|warfarin 5 mg intravenous powder for injection
C0981139|WARFARIN SODIUM 5MG/VIL INJ
C0981139|Warfarin Sodium For Inj 5 MG
C0981139|Warfarin Sodium 2 MG/ML Injectable Solution
C0981139|WARFARIN NA 5MG/VIL INJ
C0981139|WARFARIN NA 5MG/VIL INJ [VA Product]
C0981139|Warfarin 5mg Lyophilisate for solution for injection
C0981139|Warfarin Sodium 5 MG Intravenous Powder for Solution
C0981141|Warfarin Sodium 7.5mg Oral tablet
C0981141|Warfarin Sodium, 7.5 mg oral tablet
C0981141|warfarin 7.5 mg oral tablet
C0981141|WARFARIN (COUMADIN) NA 7.5MG TAB
C0981141|WARFARIN (COUMADIN) NA 7.5MG TAB UD
C0981141|Warfarin Sodium Tab 7.5 MG
C0981141|Warfarin Sodium 7.5 MG Oral Tablet
C0981141|WARFARIN NA (GOLDEN STATE) 7.5MG TAB
C0981141|WARFARIN NA 7.5MG TAB,UD [VA Product]
C0981141|WARFARIN SODIUM 7.5 mg ORAL TABLET [Warfarin Sodium]
C0981141|WARFARIN NA (GOLDEN STATE) 7.5MG TAB [VA Product]
C0981141|WARFARIN NA 7.5MG TAB,UD
C0981141|WARFARIN NA 7.5MG TAB [VA Product]
C0981141|WARFARIN NA 7.5MG TAB
C0981141|WARFARIN NA (EXELAN) 7.5MG TAB
C0981141|WARFARIN NA (EXELAN) 7.5MG TAB [VA Product]
C0981141|Warfarin sodium 7.5mg tablet (product)
C0981141|Warfarin sodium 7.5mg tablet
C0981794|Warfarin Sodium 3mg Oral tablet
C0981794|Warfarin Sodium, 3 mg oral tablet
C0981794|warfarin 3 mg oral tablet
C0981794|WARFARIN (COUMADIN) NA 3MG TAB
C0981794|WARFARIN (COUMADIN) NA 3MG TAB UD
C0981794|Warfarin Sodium Tab 3 MG
C0981794|Warfarin Sodium 3 MG Oral Tablet
C0981794|WARFARIN NA (GOLDEN STATE) 3MG TAB
C0981794|WARFARIN NA (GOLDEN STATE) 3MG TAB [VA Product]
C0981794|WARFARIN NA 3MG TAB [VA Product]
C0981794|WARFARIN NA 3MG TAB,UD
C0981794|WARFARIN SODIUM 3 mg ORAL TABLET [Warfarin Sodium]
C0981794|WARFARIN NA 3MG TAB
C0981794|WARFARIN NA 3MG TAB,UD [VA Product]
C0981794|WARFARIN NA (EXELAN) 3MG TAB
C0981794|WARFARIN NA (EXELAN) 3MG TAB [VA Product]
C0981794|Warfarin sodium 3mg tablet
C0981794|Warfarin sodium 3mg tablet (product)
C0981794|Warfarin sodium 3mg tablet (substance)
C0981140|Warfarin Sodium 6mg Oral tablet
C0981140|Warfarin Sodium, 6 mg oral tablet
C0981140|warfarin 6 mg oral tablet
C0981140|WARFARIN (COUMADIN) NA 6MG TAB
C0981140|WARFARIN (COUMADIN) NA 6MG TAB UD
C0981140|Warfarin Sodium Tab 6 MG
C0981140|Warfarin Sodium 6 MG Oral Tablet
C0981140|WARFARIN NA (GOLDEN STATE) 6MG TAB
C0981140|WARFARIN NA (GOLDEN STATE) 6MG TAB [VA Product]
C0981140|WARFARIN NA 6MG TAB
C0981140|WARFARIN NA 6MG TAB,UD [VA Product]
C0981140|WARFARIN NA 6MG TAB [VA Product]
C0981140|WARFARIN NA 6MG TAB,UD
C0981140|Warfarin Sodium 6 mg ORAL TABLET [Warfarin Sodium]
C0981140|WARFARIN NA (EXELAN) 6MG TAB
C0981140|WARFARIN NA (EXELAN) 6MG TAB [VA Product]
C0981140|Warfarin sodium 6mg tablet (product)
C0981140|Warfarin sodium 6mg tablet
C0981793|Warfarin Sodium 5mg Oral tablet
C0981793|Warfarin Sodium, 5 mg oral tablet
C0981793|warfarin 5 mg oral tablet
C0981793|WARFARIN (COUMADIN) NA 5MG TAB UD
C0981793|WARFARIN (COUMADIN) NA 5MG TAB
C0981793|Warfarin Sodium Tab 5 MG
C0981793|Warfarin Sodium 5 MG Oral Tablet
C0981793|WARFARIN NA (GOLDEN STATE) 5MG TAB
C0981793|WARFARIN NA 5MG TAB,UD
C0981793|WARFARIN NA 5MG TAB,UD [VA Product]
C0981793|WARFARIN SODIUM 5 mg ORAL TABLET [Warfarin Sodium]
C0981793|WARFARIN NA 5MG TAB
C0981793|WARFARIN NA (GOLDEN STATE) 5MG TAB [VA Product]
C0981793|WARFARIN NA 5MG TAB [VA Product]
C0981793|WARFARIN NA (EXELAN) 5MG TAB
C0981793|WARFARIN NA (EXELAN) 5MG TAB [VA Product]
C0981793|Warfarin sodium 5mg tablet
C0981793|Warfarin sodium 5mg tablet (product)
C0981793|Warfarin sodium 5mg tablet (substance)
C0917972|Athrombin-K
C0981136|Warfarin Sodium 2.5mg Oral tablet
C0981136|Warfarin Sodium, 2.5 mg oral tablet
C0981136|warfarin 2.5 mg oral tablet
C0981136|WARFARIN (COUMADIN) NA 2.5MG TAB
C0981136|WARFARIN (COUMADIN) NA 2.5MG TAB UD
C0981136|Warfarin Sodium Tab 2.5 MG
C0981136|Warfarin Sodium 2.5 MG Oral Tablet
C0981136|WARFARIN NA (GOLDEN STATE) 2.5MG TAB
C0981136|WARFARIN NA 2.5MG TAB,UD
C0981136|WARFARIN NA 2.5MG TAB,UD [VA Product]
C0981136|WARFARIN SODIUM 2.5 mg ORAL TABLET [Warfarin Sodium]
C0981136|WARFARIN NA (GOLDEN STATE) 2.5MG TAB [VA Product]
C0981136|WARFARIN NA 2.5MG TAB [VA Product]
C0981136|WARFARIN NA 2.5MG TAB
C0981136|WARFARIN NA (EXELAN) 2.5MG TAB [VA Product]
C0981136|WARFARIN NA (EXELAN) 2.5MG TAB
C0981136|Warfarin sodium 2.5mg tablet (product)
C0981136|Warfarin sodium 2.5mg tablet
C0043031|Warfarin
C0043031|2H-1-Benzopyran-2-one, 4-hydroxy-3-(3-oxo-1-phenylbutyl)-
C0043031|4-Hydroxy-3-(3-oxo-1-phenylbutyl)-2H-1-benzopyran-2-one
C0043031|3-(Alpha-acetonylbenzyl)-4-hydroxycoumarin
C0043031|3-Alpha-phenyl-beta-acetylethyl-4-hydroxycoumarin
C0043031|1-(4'-Hydroxy-3'-coumarinyl)-1-phenyl-3-butanone
C0043031|Warfarin [Chemical/Ingredient]
C0043031|3-(.alpha.-Acetonylbenzyl)-4-hydroxycoumarin
C0043031|3-(.alpha.-Phenyl-.beta.-acetylethyl)-4-hydroxycoumarin
C0043031|warfarin (medication)
C0043031|anticoagulants warfarin
C0043031|Warfarin (product)
C0043031|Warfarin (substance)
C0043031|WARF
C0981134|Warfarin Sodium 10mg Oral tablet
C0981134|Warfarin Sodium, 10 mg oral tablet
C0981134|warfarin 10 mg oral tablet
C0981134|WARFARIN (COUMADIN) NA 10MG TAB
C0981134|WARFARIN (COUMADIN) NA 10MG TAB UD
C0981134|Warfarin Sodium Tab 10 MG
C0981134|Warfarin Sodium 10 MG Oral Tablet
C0981134|WARFARIN NA (GOLDEN STATE) 10MG TAB
C0981134|WARFARIN NA 10MG TAB,UD
C0981134|WARFARIN NA 10MG TAB
C0981134|WARFARIN NA 10MG TAB,UD [VA Product]
C0981134|WARFARIN SODIUM 10 mg ORAL TABLET [Warfarin Sodium]
C0981134|WARFARIN NA 10MG TAB [VA Product]
C0981134|WARFARIN NA (GOLDEN STATE) 10MG TAB [VA Product]
C0981134|Warfarin Sodium 10 MG Oral Tablet [PANWARFIN]
C0981134|WARFARIN NA (EXELAN) 10MG TAB
C0981134|WARFARIN NA (EXELAN) 10MG TAB [VA Product]
C0981134|Warfarin sodium 10mg tablet (product)
C0981134|Warfarin sodium 10mg tablet
C1584930|Warfarin Sodium 2mg Oral tablet
C1584930|Warfarin Sodium, 2 mg oral tablet
C1584930|warfarin 2 mg oral tablet
C1584930|WARFARIN (COUMADIN) NA 2MG TAB
C1584930|WARFARIN (COUMADIN) NA 2MG TAB UD
C1584930|Warfarin Sodium Tab 2 MG
C1584930|Warfarin Sodium 2 MG Oral Tablet
C1584930|WARFARIN NA (GOLDEN STATE) 2MG TAB
C1584930|WARFARIN NA 2MG TAB [VA Product]
C1584930|WARFARIN NA 2MG TAB
C1584930|WARFARIN SODIUM 2 mg ORAL TABLET [Warfarin Sodium]
C1584930|WARFARIN NA 2MG TAB,UD
C1584930|WARFARIN NA (GOLDEN STATE) 2MG TAB [VA Product]
C1584930|WARFARIN NA 2MG TAB,UD [VA Product]
C1584930|WARFARIN NA (EXELAN) 2MG TAB
C1584930|WARFARIN NA (EXELAN) 2MG TAB [VA Product]
C1584930|Warfarin sodium 2mg tablet (product)
C1584930|Warfarin sodium 2mg tablet
C1584930|Warfaren sodium 2mg tablet usp
C0376218|Sodium, Warfarin
C0376218|Warfarin Sodium
C0376218|warfarin sodium (medication)
C0376218|Warfarin Sodium [Chemical/Ingredient]
C0376218|Warfarin sodium (substance)
C0376218|Prothromadin
C0376218|Sodium warfarin
C0376218|Tintorane
C1572765|WARFARIN SODIUM ISOPROPANOL COMPLEX
C1601608|Warfin
C0163698|2H-1-Benzopyran-2-one, 3-(1-(4-azidophenyl)-3-oxobutyl)-4-hydroxy-
C0163698|azidowarfarin
C0298589|warfarin hexadecyl ether
C0265374|Dysmorphism due to warfarin
C0265374|Foetal warfarin syndrome
C0265374|Congenital warfarin syndrome
C0265374|Warfarin syndrome
C0265374|Fetal anticoagulant syndrome
C0265374|Coumarin syndrome
C0265374|Warfarin embryopathy
C0265374|DiSala syndrome
C0265374|Fetal Warfarin Syndrome
C0265374|Fetal warfarin syndrome (disorder)
C0265374|Fetal Coumadin Syndrome
C0265374|dysmorphism; warfarin
C0265374|warfarin; dysmorphism
C0282378|Potassium, Warfarin
C0282378|Warfarin Potassium
C0282378|warfarin potassium (discontinued) (medication)
C0282378|warfarin potassium (discontinued)
C0282378|Potassium warfarin
C0282378|Potassium warfarin (substance)
C0588999|Warfarin - rodenticide
C0588999|Warfarin - rodenticide (substance)
C1975542|Warfarin &#x7C; urine
C2966895|Warfarin &#x7C; XXX
C0366686|Warfarin:Mass:Pt:Dose:Qn
C0366686|Warfarin [Mass] of Dose
C0366686|Warfarin Dose
C0366686|Warfarin:Mass:Point in time:Dose med or substance:Quantitative
C1975540|Warfarin &#x7C; bld-ser-plas
C1975541|Warfarin &#x7C; gastric fluid
C0647187|3'-hydroxywarfarin
C0648649|N-acetyl-gamma-glutamyl-4'-aminowarfarin
C0648649|AGAW
C0049626|4,6-dihydroxy-3-(3-oxo-1-phenylbutyl)-2H-1- benzopyran-2-one
C0049626|6-hydroxywarfarin
C0639160|6-methyl-6,12-methano-6H,12H,13H-benzopyran(4,3-d)benzodioxocin-13-one
C0639160|MMBBD
C0207897|4'-aminowarfarin
C0207897|3-(1-(4-aminophenyl)-3-oxobutyl)-4-hydroxy-2H-1-benzopyran-2-one
C0529816|8-hydroxywarfarin
C0637401|4-hydroxy-3-(1-(4-hydroxyphenyl)-3-oxobutyl)-2H-1-benzopyran-2-one
C0637401|4'-hydroxywarfarin
C2363289|Coumafuryl
C2363289|Coumafuryl (substance)
C2363289|Coumafuryl (product)
C0627500|MS-warfarin
C0627500|methylsulfinylwarfarin
C0642757|4-hydroxy-3-(2-hydroxy-3-oxo-1-phenylbutyl)-2H-1-benzopyran-2-one
C0642757|10-hydroxywarfarin
C0255975|7-hydroxywarfarin
C0255975|2H-1-Benzopyran-2-one, 4,7-dihydroxy-3-(3-oxo-1-phenylbutyl)-
C1276897|Warfarin Sodium 0.5 MG Oral Tablet
C1276897|Warfarin sodium 0.5mg tablet (product)
C1276897|Warfarin sodium 0.5mg tablet
C1276897|Warfarin sodium 0.5mg tablet (substance)
C1527323|Rodex
C1527323|Rodex brand of warfarin
C1520121|Co-Rax
C1520122|Compound 42
C1520123|WARF Compound 42
C0699129|Coumadin
C0699129|Marevan
C0699129|Bristol-Myers Squibb Brand of Warfarin Sodium
C0699129|Goldshield Brand of Warfarin Sodium
C0699129|Boots Brand of Warfarin Sodium
C1564392|Genpharm Brand of Warfarin Sodium
C1564392|Gen-Warfarin
C1564393|Aldo Brand of Warfarin Sodium
C1564393|Aldocumar
C1564394|Coumadine
C1564394|Bailly Brand of Warfarin Sodium
C1564395|Apo-Warfarin
C1564395|Apotex Brand of Warfarin Sodium
C1564396|Estedi Brand of Warfarin Sodium
C1564396|Tedicumar
C1564397|Warfant
C1564397|Antigen Brand of Warfarin Sodium
C1330361|Jantoven
C1601605|Narfarin
C1601620|Marfarin
C0605881|actosin P
C0605881|pindone, warfarin drug combination
C0605881|pindone - warfarin
C0699130|Panwarfin
C1996947|Parenteral form warfarin
C1996947|Parenteral form warfarin (product)
C1998178|Oral form warfarin
C1998178|Oral form warfarin (product)
