C1122548|NS4A cofactor peptide, Hepatitis C virus
C0015506|Factor VIII
C0086277|Factor VIII Coagulant Antigen
C0015491|factor IX
C1394921|deficiency; clotting factor, VIII, with vascular defect
C0200408|Coagulation factor IX measurement
C4067217|acquired clotting factor inhibitors - factor ix
C1394911|deficiency; clotting factor, IX (congenital) (functional) (hereditary) (with functional defect)
C0199967|Transfusion of coagulation factors
C0852255|Blood and blood product treatment
C0614404|asialo-Factor VIII
C0614404|asialofactor VIII
C0626325|Factor VIII Leiden
C0627512|Kryobulin TIM3
C0633201|(des-797-1562)-factor VIII
C0633201|factor VIII (des-797-1562)
C0644521|factor VIII delta II
C0644521|factor VIII deltaII
C0711027|Koate-HP, human intravenous powder for injection
C0354641|Factor VIII fraction products
C0354641|Human antihaemophilic fraction
C0354641|Human antihemophilic fraction
C0354641|Human coagulation factor VIII
C0354641|Factor VIII fraction products (product)
C0354641|Factor VIII fraction products (substance)
C0724529|Porcine Factor VIII
C0724529|antihemophilic factor, porcine
C0724529|ANTIHEMOPHILIC FACTOR,PORCINE
C0724529|Porcine factor VIII (product)
C0724529|Porcine factor VIII (substance)
C0724529|Porcine antihaemophilic factor agent
C0724529|Porcine antihaemophilic factor
C0724529|Porcine antihemophilic factor agent (substance)
C0724529|Porcine antihemophilic factor agent
C0724529|Porcine antihemophilic factor
C0740130|Hemofil-M
C0740130|Hemofil
C0740130|Hemophil
C0740130|Hemofil M
C0740130|Hemofil HM
C0795577|recombinant antihemophilic factor VIII
C0795577|Factor VIII Recombinant
C0541364|FVIII Ise
C0541364|factor VIII Ise
C0591821|Monoclate-P
C0591821|Monoclate-P (obsolete)
C2342443|Xyntha
C2342443|Factor VIII (Xyntha)
C2342443|Factor VIII (Xyntha) (medication)
C0015514|Activated Factor VIII
C0015514|Factor VIII, Thrombin Activated
C0015514|Factor VIIIa
C0015514|Thrombin-Activated Factor VIII
C0015514|Blood-coagulation factor VIIIa, procoagulant
C0015514|Factor VIIIa, Coagulation
C0015514|VIIIa, Coagulation Factor
C0015514|COAG FACTOR VIIIA
C0015514|BLOOD COAG FACTOR VIII ACTIVATED
C0015514|Factor VIIIa [Chemical/Ingredient]
C0015514|Coagulation Factor VIIIa
C0015514|Factor VIII, Thrombin-Activated
C0015514|Factor VIII, Activated
C0015514|Blood Coagulation Factor VIII, Activated
C0015514|Coagulation factor VIIIa (substance)
C0015506|Factor VIII
C0015506|coagulation factor VIII
C0015506|Blood-coagulation factor VIII, complex
C0015506|antihemophilic factor
C0015506|COAG FACTOR VIII
C0015506|BLOOD COAG FACTOR VIII
C0015506|antihemophilic factor A
C0015506|thromboplastinogen A
C0015506|platelet cofactor I
C0015506|hematological agents antihemophilic factors
C0015506|antihemophilic factors
C0015506|antihemophilic factors (medication)
C0015506|Thromboplastinogen
C0015506|Blood Coagulation Factor VIII
C0015506|Factor VIII [Chemical/Ingredient]
C0015506|Coagulation factor VIII (substance)
C0015506|Factor viii (antihemophilic factor, human) per i.u.
C0015506|AHF
C0015506|AHG
C0015506|Antihemophilic globulin
C0015506|Antihaemophilic factor
C0015506|Factor VIII (substance)
C0015506|Antihaemophilic factor A
C0015506|Antihaemophilic globulin
C0015506|Coagulation factor VIII (substance) [Ambiguous]
C0015506|Factor VIII product (product)
C0015506|Factor VIII product
C0020199|Hyate C
C0020199|Hyatt C
C0020199|Hyate:C
C0020199|Hyate C (obsolete)
C0020199|HyateC
C0020199|HyattC
C0020199|Hyate-C
C0020199|Hyatt-C
C0020199|Speywood Brand of Porcine Factor VIII Preparation
C2825466|Moroctocog alfa (product)
C2825466|Moroctocog alfa
C2825466|Moroctocog alfa (substance)
C2825466|Antihemophilic Factor, Human Recombinant Residues 743-1636 Deleted
C0971600|ReFacto
C0971600|refacto (medication)
C0218184|Kogenate
C0218184|Kogenate Bayer
C0218184|Kogenate (obsolete)
C0218184|Factor VIII (Kogenate)
C0218184|Factor VIII (Kogenate) (medication)
C0218184|recombinant antihemophilic factor VIII
C0700346|antihemophilic factor, human
C0700346|Antihemophilic Factor Human
C0700346|ANTIHEMOPHILIC FACTOR,HUMAN
C2927721|Factor VIII/von Willebrand Factor Complex Human Plasma
C2732002|Recombinant antihemophilic factor agent
C2732002|Recombinant antihaemophilic factor agent
C2732002|antihemophilic factor, recombinant
C2732002|ANTIHEMOPHILIC FACTOR, HUMAN RECOMBINANT
C2732002|FVIII
C2732002|Factor VIII
C2732002|ANTIHEMOPHILIC FACTOR,RECOMBINANT
C2732002|Recombinant human factor VIII - Octocog alpha
C2732002|DNA factor VIII (product)
C2732002|Octocog alpha
C2732002|Recombinant antihaemophilic factor preparation
C2732002|Recombinant antihemophilic factor agent (substance)
C2732002|Recombinant antihemophilic factor preparation
C2732002|DNA factor VIII (substance)
C2732002|Recombinant antihemophilic factor preparation (substance)
C2732002|Recombinant antihemophilic factor agent (product)
C2732002|Recombinant human factor VIII
C2601455|Coagulation factor VIII &#x7C; Platelet poor plasma
C2968287|Factor VIII &#x7C; patient
C1985551|Coagulation factor VIII activity.Xa activator &#x7C; platelet poor plasma
C1976512|Transfuse factor VIII &#x7C; patient
C0086277|FACTOR VIII COAG ANTIGEN
C0086277|Coagulation factor VIII Ag
C0086277|Coagulation factor VIII Antigen
C0086277|Factor VIII Clotting Antigen
C0086277|Factor VIII Ag
C0086277|Factor VIII antigen
C0086277|Factor VIII antigen (substance)
C0086277|Factor VIII Coagulant Antigen
C2968288|Factor VIII units &#x7C; Blood product unit
C1985549|Coagulation factor VIII Ab &#x7C; platelet poor plasma
C1985548|Coagulation factor VIII &#x7C; XXX
C2601456|Coagulation factor VIII activity &#x7C; Platelet poor plasma
C1985550|Coagulation factor VIII activated &#x7C; platelet poor plasma
C2359705|Transfuse factor VIII &#x7C; Blood product unit
C1307126|Antihemophilic Factor
C1307126|factor VIII, human
C1307126|AHF
C1307126|F8 protein, human
C1307126|FVIII protein, human
C1307126|coagulation factor VIII, procoagulant component (hemophilia A) protein, human
C1307126|Factor VIII
C1307126|Coagulation Factor VIII
C1307126|Coagulation Factor VIIIc
C1307126|F8
C1307126|Factor VIII F8B
C1307126|Antihaemophilic Factor
C1307126|Procoagulant Component
C0086428|Humate-P
C0086428|Humate-P (obsolete)
C2726511|Wilate
C0594139|Alphanate
C0594139|Alphanate (obsolete)
C3660038|N8-GP compound
C3529561|N8 rFVIII
C3529561|N8 recombinant factor VIII
C3529561|recombinant factor VIII N8
C1815380|Optivate
C3849397|factor VIII-Fc fusion protein
C3849397|rFVIIIFc protein
C3859470|Obizur
C3859426|antihemophilic factor, porcine B-domain truncated recombinant
C3859426|ANTIHEMOPHILIC FACTOR PORCINE, B-DOMAIN TRUNCATED RECOMBINANT
C4018188|Novoeight
C4031949|antihemophilic factor (recombinant), porcine sequence (medication)
C4031949|antihemophilic factor (recombinant), porcine sequence
C3834170|factor VIII (b-domain deleted recombinant) FC fusion protein
C3834170|antihemophilic factor, recombinant Fc fusion protein
C3834170|antihemophilic factor (recombinant), fc fusion protein (medication)
C3834170|antihemophilic factor (recombinant), fc fusion protein
C3834170|efmoroctocog alfa
C4038482|Factor VIII+von Willebrand factor.ristocetin cofactor
C4045418|BAY 94-9027
C4057564|Koate
C0376176|Monoclate
C1300015|Antihemophilic Factor (Human) For Inj 1000 Unit
C1300015|Antihemophilic Factor (Human) For Inj 220-400 Unit
C1300015|Antihemophilic Factor (Human) For Inj 250 Unit
C1300015|Antihemophilic Factor (Human) For Inj 401-800 Unit
C1300015|Antihemophilic Factor (Human) For Inj 500 Unit
C1300015|Antihemophilic Factor (Human) For Inj Kit 250 Unit
C1300015|Antihemophilic Factor (Human) For Inj Kit 500 Unit
C1300015|antihemophilic factor human intravenous powder for injection
C1300015|antihemophilic factor (obsolete) human intravenous powder for injection
C1300015|Antihemophilic factor agent 500 iu powder for injection solution 5mL vial + diluent (product)
C1300015|Antihemophilic factor agent 1500 iu powder for injection solution 5mL vial + diluent (product)
C1300015|Antihaemophilic factor agent 500 iu powder for injection solution 5mL vial + diluent
C1300015|Antihemophilic factor agent 500 iu powder for injection solution 5mL vial + diluent
C1300015|Antihemophilic factor agent 1000 iu powder for injection solution 5mL vial + diluent
C1300015|Antihaemophilic factor agent 1500 iu powder for injection solution 5mL vial + diluent
C1300015|Antihaemophilic factor agent 1000 iu powder for injection solution 5mL vial + diluent
C1300015|Antihemophilic factor agent 1000 iu powder for injection solution 5mL vial + diluent (product)
C1300015|Antihemophilic factor agent 1500 iu powder for injection solution 5mL vial + diluent
C1300015|Antihemophilic Factor VIII Human 1 IU Intravenous Powder for Solution
C1300015|ANTIHEMOPHILIC FACTOR,HUMAN INJ
C1300015|ANTIHEMOPHILIC FACTOR,HUMAN INJ [VA Product]
C1300015|Antihemophilic Factor VIII Human 1 IU Injection Powder for Solution
C1300015|Antihemophilic Factor VIII Human Intravenous Powder for Solution
C1300015|Antihemophilic Factor VIII Human 1 IU Injection Powder for Solution [FACTOR VIII:C]
C1300015|Antihemophilic Factor (Human) For Inj 801-1500 Unit
C1300015|Antihemophilic Factor (Human) For Inj 1501-2000 Unit
C1300015|Antihemophilic Factor VIII Human/Antihemophilic Factor VIII:C Human 1 IU-1 IU Intravenous Powder for Solution
C1300015|Antihemophilic Factor (Human) For Inj 1700 Unit
C1300015|factor VIII, human 1 UNT Injection
C1300015|antihemophilic factor, human 1 UNT Injection
C1300015|Antihaemophilic factor 500unt/vial powder
C1300015|Antihemophilic factor 500unt/vial powder (product)
C1300015|Antihemophilic factor 500unt/vial powder
C1300015|Antihemophilic Factor VIII:C Human 1 IU Intravenous Powder for Solution
C0543246|antihemophilic factor (obsolete) porcine intravenous powder for injection
C0543246|antihemophilic factor porcine intravenous powder for injection
C0543246|Porcine factor VIII 700iu injection
C0543246|Antihemophilic Factor VIII:C (Porcine) 1 U Injection Powder for Solution
C0543246|Antihemophilic Factor VIII (Porcine) Injection Powder for Solution
C0543246|Antihemophilic Factor VIII (Porcine) 1 IU Injection Powder for Solution
C0543246|Antihemophilic Factor VIII (Porcine) 1 U Intravenous Powder for Solution
C0543246|Porcine factor VIII 700iu powder for injection solution vial (product)
C0543246|Porcine factor VIII 700iu powder for injection solution vial
C0543246|Porcine factor VIII 700iu injection (product)
C0543246|Porcine factor VIII 700iu injection (substance)
C4064080|simoctocog alfa
C4064080|simoctocog alfa (medication)
C4064080|antihemophilic factors simoctocog alfa
C4064080|coagulation factor VIII, B-domain deleted recombinant
C4074414|Nuwiq
C3529563|turoctocog alfa
C3529563|antihemophilic factor, human B-domain truncated recombinant
C0732093|Factor VIII + von Willebrand factor
C0732093|factor VIII, von Willebrand factor drug combination
C0732093|factor VIII - von Willebrand factor
C0732093|Factor VIII / von Willebrand factor
C0732093|Factor VIII+von Willebrand factor
C0732093|Factor VIII+von Willebrand factor (product)
C0732093|Factor VIII+von Willebrand factor (substance)
C0358606|Activated prothrombin complex concentrate
C0358606|Factor VIII by-passing fraction products
C0358606|Factor VIII by-passing fraction products (product)
C0358606|Factor VIII by-passing fraction products (substance)
C0720828|Helixate
C0720828|Helixate (obsolete)
C1815247|Monarc-M
C1815247|Monarc-M (obsolete)
C0218182|Recombinate
C0218182|Recombinate (obsolete)
C1691209|Octocog alfa
C1691209|Octocog alfa (product)
C1691209|DNA factor VIII
C1691209|Deoxyribonucleic acid factor VIII
C1691209|Deoxyribonucleic acid factor VIII (product)
C1691209|Octocog alfa (substance)
C0056540|cryobulin
C0056545|cryoprecipitate coagulum
C0961271|BAY 14-2222
C0961271|BAY-14-2222
C0961271|BAY14-2222
C0966326|malmo protocol
C0966500|r-VIII SQ
C0966500|recombinant factor VIII SQ
C1098523|rFVIII-FS
C1098523|recombinant FVIII, sugar formulated
C1121470|B-domain-deleted factor VIII
C1121470|GC-rAHF
C1121470|rFVIII (B-domain-deleted)
C1175691|8Y factor VIII-von Willebrand factor concentrate
C1175691|factor VIII-von Willebrand factor concentrate 8Y
C1175691|vWF-FVllI 8Y
C0731320|Haemate P
C2002589|Immunate solvent detergent, human
C1815260|Advate
C1985553|Coagulation factor VIII Ag &#x7C; Tissue and Smears
C1985552|Coagulation factor VIII Ag &#x7C; platelet poor plasma
C0015494|Activated Factor IX
C0015494|Factor IXa
C0015494|Factor IXa, Coagulation
C0015494|IXa, Coagulation Factor
C0015494|BLOOD COAG FACTOR IX ACTIVATED
C0015494|COAG FACTOR IXA
C0015494|FACTOR VIIIIA
C0015494|FACTOR VIIII ACTIVATED
C0015494|COAGULATION FACTOR VIIIIA
C0015494|Coagulation factor IXa -RETIRED-
C0015494|Coagulation Factor IXa
C0015494|Factor IX, Activated
C0015494|Blood Coagulation Factor IX, Activated
C0015494|Factor IXa [Chemical/Ingredient]
C0015494|Coagulation factor IXa (substance)
C0015494|Activated Christmas Factor
C0015491|Factor IX
C0015491|Christmas factor
C0015491|coagulation factor IX
C0015491|Blood-coagulation factor IX
C0015491|Complex, Factor IX
C0015491|Fraction, Factor IX
C0015491|IX Complex, Factor
C0015491|IX Fraction, Factor
C0015491|Factor IX, Coagulation
C0015491|IX, Coagulation Factor
C0015491|COAGULATION FACTOR VIIII
C0015491|COAG FACTOR IX
C0015491|FACTOR VIIII
C0015491|BLOOD COAG FACTOR IX
C0015491|antihemophilic factor B
C0015491|autoprothrombin II
C0015491|thromboplastinogen B
C0015491|Factor IX Complex
C0015491|Plasma Thromboplastin Component
C0015491|Factor IX Fraction
C0015491|Blood Coagulation Factor IX
C0015491|Factor IX [Chemical/Ingredient]
C0015491|PTC
C0015491|IX
C0015491|Platelet cofactor II
C0015491|Coagulation factor IX (substance)
C0015491|Antihaemophilic factor B
C1170091|BeneFIX
C1170091|Benefix (obsolete)
C0060018|factor IX Long Beach
C0060018|FIX-LB
C0082540|factor IX-antithrombin III complex
C0082540|factor IX-ATIII complex
C0082536|factor IX Leyden
C0082536|Leyden factor IX
C0060011|BM Lake Elsinore factor IX
C0060011|factor IX BM Lake Elsinore
C0060011|Factor IX BmLE
C0060014|Blood-coagulation factor IX Chapel Hill
C0060014|factor IX Chapel Hill
C0297142|Mononine
C0297142|Mononine (obsolete)
C0297142|Mononine (obsolete1)
C0289773|factor IX (1-47)
C0251224|factor IX Strasbourg 2
C0117201|factor IX Madrid
C0060013|factor IX Cardiff
C0117199|factor IX Cambridge
C0117199|factor IX propeptide
C0718844|Bebulin VH
C0718844|Bebulin VH (obsolete)
C0592047|Replenine
C2826076|Factor IX, recombinant
C2826076|Coagulation Factor IX Recombinant Human
C2826076|FACTOR IX,RECOMBINANT
C2826076|coagulation factor IX (recombinant human)
C3666839|Rixubis
C3644708|Kcentra
C0718417|Alphanine SD
C0718417|Alphanine SD (obsolete)
C0718417|Alphanine SD (obsolete1)
C2972532|Transfuse factor IX &#x7C; patient
C1985535|Coagulation factor IX activated &#x7C; platelet poor plasma
C2601448|Coagulation factor IX &#x7C; Platelet poor plasma
C2972533|Transfuse factor IX units &#x7C; Blood product unit
C1985536|Coagulation factor IX Ag &#x7C; platelet poor plasma
C2601449|Coagulation factor IX activity &#x7C; Platelet poor plasma
C2968286|Factor IX &#x7C; patient
C2749016|THROMBOPHILIA, X-LINKED, DUE TO FACTOR IX DEFECT
C2749016|THPH8
C3657751|IB1001
C3657751|IB1001 trenacog alfa
C4048712|factor IX complex
C4048712|coagulation factor IX
C4048712|Factor IX complex agent
C4048712|factor IX complex, human
C4048712|FACTOR IX COMPLEX,HUMAN
C4048712|Coagulation Factor IX Complex Human
C4048712|Factor IX complex preparation
C4048712|Factor IX preparation
C4048712|Factor IX complex agent (substance)
C4048712|Factor IX agent
C4048712|Factor IX complex preparation (substance)
C3883805|N9-GP compound
C3883805|nonacog beta pegol
C3883952|factor IX Padua
C3883952|factor IX-Padua
C0722828|Profilnine SD
C4041753|rFIXFc protein
C4041753|factor IX Fc fusion protein
C4051373|Ixinity
C1269927|Coagulation Factor IX (Recombinant) For Inj 1000 Unit
C1269927|Coagulation Factor IX (Recombinant) For Inj 250 Unit
C1269927|Coagulation Factor IX (Recombinant) For Inj 500 Unit
C1269927|coagulation factor IX recombinant intravenous powder for injection
C1269927|Coagulation Factor IX (Recombinant) For Inj 2000 Unit
C1269927|FACTOR IX,RECOMBINANT 1000 UNT/VIL INJ
C1269927|FACTOR IX,RECOMBINANT 1000 UNT/VIL INJ [VA Product]
C1269927|Coagulation Factor IX Recombinant 1 IU Intravenous Powder for Solution
C1269927|Coagulation Factor IX Recombinant Powder for solution for injecti with Alcohol Pad or Swab - IV Administration Set (unspecified) - Filter Spike - Double-Ended Needle - Sterile Water for Injection -
C1269927|Coagulation Factor IX (Recombinant) For Inj 3000 Unit
C1269927|FACTOR IX,RECOMBINANT 3000 UNIT/VIL INJ
C1269927|FACTOR IX,RECOMBINANT 2000 UNIT/VIL INJ
C1269927|FACTOR IX,RECOMBINANT 2000 UNIT/VIL INJ [VA Product]
C1269927|FACTOR IX,RECOMBINANT 3000 UNIT/VIL INJ [VA Product]
C1269927|Coagulation Factor IX (Recomb) (rFIXFc) For Inj 500 Unit
C1269927|Coagulation Factor IX (Recomb) (rFIXFc) For Inj 2000 Unit
C1269927|Coagulation Factor IX Recombinant Lyophilisate for solution for injecti with Vial adapter - Diluent -
C1269927|Coagulation Factor IX (Recomb) (rFIXFc) For Inj 1000 Unit
C1269927|Coagulation Factor IX (Recomb) (rFIXFc) For Inj 3000 Unit
C1269927|Coagulation Factor IX (Recombinant) For Inj 1500 Unit
C1269927|FACTOR IX,RECOMBINANT (THR148) 1500 UNIT/VIL INJ [VA Product]
C1269927|FACTOR IX,RECOMBINANT (THR148) 1000 UNIT/VIL INJ
C1269927|FACTOR IX,RECOMBINANT (THR148) 500 UNIT/VIL INJ
C1269927|FACTOR IX,RECOM(THR148) 1000UNIT/VIL INJ
C1269927|FACTOR IX,RECOM(THR148) 1500UNIT/VIL INJ
C1269927|FACTOR IX,RECOM(THR148) 500UNIT/VIL INJ
C1269927|FACTOR IX,RECOMBINANT (THR148) 1500 UNIT/VIL INJ
C1269927|FACTOR IX,RECOMBINANT (THR148) 500 UNIT/VIL INJ [VA Product]
C1269927|FACTOR IX,RECOMBINANT (THR148) 1000 UNIT/VIL INJ [VA Product]
C1269927|coagulation factor IX (recombinant human) 1 UNT Injection
C1269927|Recombinant coagulation factor IX 1000iu injection (pdr for recon)+solvent
C1269927|Recombinant coagulation factor IX 1000iu powder and solvent for injection solution vial (product)
C1269927|Recombinant coagulation factor IX 1000iu powder and solvent for injection solution vial
C1269927|Recombinant coagulation factor IX 250iu injection (pdr for recon)+solvent
C1269927|Recombinant coagulation factor IX 250iu powder and solvent for injection solution vial (product)
C1269927|Recombinant coagulation factor IX 250iu powder and solvent for injection solution vial
C1269927|Recombinant coagulation factor IX 500iu injection (pdr for recon)+solvent
C1269927|Recombinant coagulation factor IX 500iu powder and solvent for injection solution vial (product)
C1269927|Recombinant coagulation factor IX 500iu powder and solvent for injection solution vial
C1269927|Recombinant coagulation factor IX 1000iu injection (pdr for recon)+solvent (product)
C1269927|Recombinant coagulation factor IX 1000iu injection (pdr for recon)+solvent (substance)
C1269927|Recombinant coagulation factor IX 250iu injection (pdr for recon)+solvent (product)
C1269927|Recombinant coagulation factor IX 250iu injection (pdr for recon)+solvent (substance)
C1269927|Recombinant coagulation factor IX 500iu injection (pdr for recon)+solvent (product)
C1269927|Recombinant coagulation factor IX 500iu injection (pdr for recon)+solvent (substance)
C1269927|Recombinant coagulation factor IX 1000iu powder for injection solution vial (product)
C1269927|Recombinant coagulation factor IX 1000iu powder for injection solution vial
C1269927|Recombinant coagulation factor IX 250iu powder for injection solution vial (product)
C1269927|Recombinant coagulation factor IX 250iu powder for injection solution vial
C1269927|Recombinant coagulation factor IX 500iu powder for injection solution vial (product)
C1269927|Recombinant coagulation factor IX 500iu powder for injection solution vial
C0724584|factor IX (human)
C0724584|coagulation factor IX human
C0724584|factor IX, human
C0724584|Factor 9
C0724584|Plasma Thromboplastic Component
C0724584|Plasma Thromboplastin Component
C0724584|PTC
C0724584|coagulation factor IX, human
C0724584|Christmas Factor
C0724584|Factor IX
C0724584|Coagulation Factor IX
C0724584|EC 3.4.21.22
C0724584|F9
C0313501|Coagulation factor IX variant (substance)
C0313501|Coagulation factor IX variant
C0313501|Coagulation factor IX variant, NOS
C1273037|Nonacog alfa
C1273037|Recombinant coagulation factor IX
C1273037|Coagulation Factor IX Recombinant
C1273037|Nonacog alfa (substance)
C1273037|Nonacog alfa (product)
C1273037|Recombinant coagulation factor IX (substance)
C1273037|Recombinant coagulation factor IX preparation (product)
C1273037|Recombinant coagulation factor IX preparation
C1815181|Konyne 80
C1815181|Konyne 80 (obsolete)
C0631906|factor IX Seattle(2)
C0631906|factor IX Seattle2
C0633767|Factor IX GLA-peptide
C0636372|Factor IX Vancouver
C0636589|factor IX Niigata
C0636589|blood coagulation factor IX Niigata
C0636589|Niigata factor IX
C0637620|factor IX San Dimas
C0637620|San Dimas factor IX
C0638162|factor IX Troed-y-Rhiw
C0638164|factor IX Kawachinagano
C0638164|factor IX KWC
C0639016|factor IX BM Nagoya
C0639016|IX Nagoya
C0640832|factor IX Chongqing
C0641637|factor IX Alabama
C0641676|factor IX Deventer
C0641677|factor IX Bergamo
C0641681|factor IX Novara
C0641682|factor IX Milano
C0643142|Factor IX Hollywood
C0643142|Factor IX (HW)
C0644057|factor IX Lincoln Park
C0645143|factor IX Basel
C0645333|factor IX Nagoya 3
C0660527|factor IX BM Hilo
C0661606|Preconativ
C0383958|factor IX Zutphen
C1121564|factor IX Denver
C2743140|factor IX, factor VII, factor X, prothrombin drug combination
C1394921|clotting factor; deficiency, VIII, with vascular defect
C1394921|deficiency; clotting factor, VIII, with vascular defect
C0200408|factor IX assay
C0200408|factor IX assay (lab test)
C0200408|factor IX level
C0200408|Coagulation factor IX level
C0200408|Clotting; factor IX (PTC or Christmas)
C0200408|Coagulation factor IX measurement
C0200408|CLOTTING FACTOR IX PTC/CHRISTMAS
C0200408|Factor IX Measurement
C0200408|CLOT FACTOR IX PTC/CHRSTMAS
C0200408|Assay for clotting factor IX (PTC)
C0200408|Clotting factor IX (PTC or Christmas) measurement
C0200408|Factor IX assay (procedure)
C0200408|Christmas Factor
C0200408|Factor IX
C0200408|FACTIX
C0200408|Clotting factor IX assay
C0200408|Christmas disease factor assay
C0200408|Hemophilia B assay
C0200408|Plasma thromboplastin component assay
C0200408|Haemophilia B assay
C0200408|Clotting factor IX assay (procedure)
C0200408|Autoprothrombin II assay
C1277707|Factor IX related antigen level
C1277707|Factor IX related antigen level (procedure)
C1277707|Factor IX related antigen measurement (procedure)
C1277707|Factor IX related antigen measurement
C2238119|factor IX antigen measurement
C2238119|factor IX antigen measurement (lab test)
C1394911|clotting factor; deficiency, IX (congenital) (functional) (hereditary) (with functional defect)
C1394911|deficiency; clotting factor, IX (congenital) (functional) (hereditary) (with functional defect)
C0199967|Clotting factor transfusion
C0199967|Coag factor transfusion
C0199967|Transfusion of coagulation factors
C0199967|Transfusion of coagulation factor
C0199967|Transfusion of coagulation factors (procedure)
C0199968|Antihaemophilic factor transfusion (procedure)
C0199968|Antihemophilic factor transfusion
C0199968|Transfusion of antihemophilic factor
C0199968|Transfusion of antihaemophilic factor
C0199968|Antihaemophilic factor transfusion
C0199968|Transfusion of antihemophilic factor (procedure)
C0199968|Antihemophilic factor transfusion (procedure)
C2242940|plasma fractions, human (treatment)
C2242940|plasma fractions, human
C3161607|plasma fractions, human factor xiii concentrate (human)
C3161607|plasma fractions, human factor xiii concentrate (human) (treatment)
C2064859|plasma fractions, human factor VIII (AHF, AHG)
C2064859|plasma fractions, human factor VIII (AHF, AHG) (treatment)
C2064857|plasma fractions, human albumin, normal serum (treatment)
C2064857|plasma fractions, human albumin, normal serum
C2064858|plasma fractions, factor IX complex (human)
C2064858|human factor IX complex (human)
C2064858|human factor IX complex (human) (treatment)
C2194217|factor VIIa transfusion (treatment)
C2194217|factor VIIa
C2194217|factor VIIa (treatment)
C2069055|plasma fractions, human albumin + globulin (treatment)
C2069055|plasma fractions, human albumin + globulin
C2069056|plasma fractions, antithrombin III (human) (treatment)
C2069056|plasma fractions, antithrombin III (human)
C4064322|plasma fractions, coagulation factor X (human) (treatment)
C4064322|plasma fractions, coagulation factor X (human)
C4064322|plasma fractions, human factor x
C1293889|Coagulation factor IX product administration by intravascular infusion
C1293889|Transfusion of factor IX (procedure)
C1293889|Transfusion of factor IX
C1293888|Coagulation factor VII product administration by intravascular infusion
C1293888|Transfusion of factor VII (procedure)
C1293888|Transfusion of factor VII
C1960763|Transfusion antithrombin III factor (procedure)
C1960763|Transfusion antithrombin III factor
C0854629|Allogenic bone marrow transplantation therapy
C0854630|Autologous bone marrow transplantation therapy
C0005842|Autotransfusion
C0005842|Autotransfusions
C0005842|Blood Transfusion, Autologous
C0005842|Autotransfusion Procedure
C0005842|TRANSFUSION AUTOL BLOOD
C0005842|BLOOD TRANSFUSIONS AUTOL
C0005842|AUTOL BLOOD TRANSFUSIONS
C0005842|TRANSFUSIONS AUTOL BLOOD
C0005842|BLOOD TRANSFUSION AUTOL
C0005842|AUTOL BLOOD TRANSFUSION
C0005842|autotransfusion (treatment)
C0005842|Blood--Transfusion, Autologous
C0005842|Autologous blood transfusion
C0005842|Blood Transfusions, Autologous
C0005842|Autologous Blood Transfusions
C0005842|Transfusion, Autologous Blood
C0005842|Transfusions, Autologous Blood
C0005842|Abt - autologous blood transfusion
C0005842|Autotransfusion (procedure)
C0005842|Autotransfusion, NOS
C0005842|Intravenous autotransfusion each treatment
C0005842|IV autotransfusion ea.Tx
C0854631|Cord blood transplant therapy
C0015236|Exchange Transfusion, Whole Blood
C0015236|blood exchange transfusion
C0015236|Exchange blood transfusion
C0015236|EXCHANGE TRANSFUSION
C0015236|exchange transfusion (treatment)
C0015236|Exchange transfusion of blood
C0015236|Exchange blood transfusion NOS
C0015236|Exchange blood transfusion NOS (procedure)
C0015236|Exchange transfusion, blood
C0015236|Transfusion replacement, total
C0015236|Exsanguination transfusion
C0015236|EBT - Exchange blood transfusion
C0015236|Exchange transfusion (procedure)
C0015236|Transfusion, exsanguination
C0854634|Mismatched donor bone marrow transplantation therapy
C0371803|Exchange transfusion, blood; newborn
C0371803|Neonatal exchange blood transfusion
C0371803|exchange transfusion of newborn (treatment)
C0371803|exchange transfusion of newborn
C0371803|Neonatal exchange transfusion
C0371803|BL EXCHANGE/TRANSFUSE NB
C0371803|EXCHNG TRANSFUSION BLOOD NEWBORN
C0371803|Exchange blood transfusion, newborn
C0371803|Exchange blood transfusion (neonatal)
C0371803|Neonatal exchange transfusion (procedure)
C0199962|packed red blood cell transfusion
C0199962|Transfusion of packed red blood cells
C0199962|Red Blood Cell Transfusion
C0199962|Transfusion of PRBC
C0199962|Intravenous blood transfusion of packed cells
C0199962|Intravenous blood transfusion of packed cells (procedure)
C0199962|Transfusion of packed red blood cells (procedure)
C0199962|PRBC Transfusion
C0199964|Plasma expander transfusion
C0199964|Blood expander transfus
C0199964|Blood expander transfusion
C0199964|Transfusion of blood expander
C0199964|Plasma expander transfusion (procedure)
C0199964|Transfusion of blood expander (procedure)
C0199964|Transfusion of plasma expander
C0199964|Transfusion of blood expander, NOS
C0199964|Transfusion of plasma expander, NOS
C0032134|Plasmaphereses
C0032134|Plasmapheresis
C0032134|Therapeu plasmapheresis
C0032134|Plasmaphoresis
C0032134|Plasma Exchange
C0032134|Plasmapheresis (procedure)
C0032134|therapeutic plasmapheresis
C0032134|Therapeutic Plasma Exchange
C0086818|Platelet Transfusion
C0086818|Platelet Transfusions
C0086818|Transfusion, Platelet
C0086818|Transfusions, Platelet
C0086818|Blood Platelet Transfusions
C0086818|Platelet Transfusion, Blood
C0086818|Platelet Transfusions, Blood
C0086818|Transfusion, Blood Platelet
C0086818|Transfusions, Blood Platelet
C0086818|transfusion of platelets (treatment)
C0086818|transfusion of platelets
C0086818|Platelet transfusion (procedure)
C0086818|Blood platelets--Transfusion
C0086818|Blood Platelet Transfusion
C0086818|Transfusion of thrombocytes
C0086818|Intravenous blood transfusion of platelets
C0086818|Intravenous blood transfusion of platelets (procedure)
C0854635|Unrelated donor bone marrow transplantation therapy
C0677960|T lymphocyte depletion therapy
C0677960|T-cell depletion
C0677960|T-Lymphocyte Depletion Therapy
C0677960|T-Cell Depletion Therapy
C0919689|Donor leukocyte infusion
C0194015|Bone marrow harvest
C0194015|aspiration of bone marrow from donor for transplant
C0194015|aspiration of bone marrow from donor for transplant (treatment)
C0194015|bone marrow collection for transplant (treatment)
C0194015|bone marrow collection for transplant
C0194015|Donor marrow aspiration
C0194015|Bone marrow harvesting
C0194015|Harvest of bone marrow
C0194015|Aspiration of bone marrow from donor for transplant (procedure)
C0023416|Leukaphereses
C0023416|Leukapheresis
C0023416|Leukocytaphereses
C0023416|Leukocytophereses
C0023416|Leukophereses
C0023416|therapeutic leukopheresis (treatment)
C0023416|therapeutic leukopheresis
C0023416|Therapeutc leukopheresis
C0023416|Leukopheresis
C0023416|Leukocytapheresis
C0023416|Leukocytopheresis
C0023416|Leucapheresis
C0023416|Leukopheresis (procedure)
C0023416|Therapeutic leukocytapheresis
C0079186|Cytaphereses
C0079186|Cytapheresis
C0411265|Blood stem cell harvest
C0411265|Stem cell harvesting
C0411265|Harvest of stem cells
C0411265|Harvest of stem cells (procedure)
C0411265|Harvesting of stem cells (procedure)
C0411265|Harvesting of stem cells
C0948144|Peripheral blood stem cell apheresis
C0948145|Erythrocytapheresis
C0948145|Erythrocytapheresis (procedure)
C0949035|Low density lipoprotein apheresis (procedure)
C0949035|Low density lipoprotein apheresis
C0949035|LDL apheresis
C0032202|Blood Plateletphereses
C0032202|Plateletphereses
C0032202|Plateletphereses, Blood
C0032202|Plateletpheresis
C0032202|Plateletpheresis, Blood
C0032202|Thrombocytaphereses
C0032202|Thrombocytophereses
C0032202|Therapeutic plateletpheresis
C0032202|cellular apheresis for platelets (treatment)
C0032202|therapeutic plateletpheresis (treatment)
C0032202|cellular apheresis for platelets
C0032202|apheresis for platelets
C0032202|Therapeu plateltpheresis
C0032202|THERAPEUTIC APHERESIS PLATELETS
C0032202|Mechanical separation of platelet cells from blood
C0032202|Therapeutic apheresis for platelets
C0032202|Therapeutic apheresis; for platelets
C0032202|Blood Plateletpheresis
C0032202|Thrombocytapheresis
C0032202|Thrombocytopheresis
C0032202|Platelet apheresis
C0032202|Plateletpheresis (procedure)
C0032202|APHERESIS PLATELETS
C0948460|Vascular catheter specimen collection
C0524864|Hematopoietic Stem Cell Mobilization
C0524864|Mobilization, Stem Cell
C0524864|Haematopoietic stem cell mobilisation
C0524864|Hematopoietic stem cell mobilisation
C0524864|Stem cell mobilisation
C0524864|Stem cell mobilization
C0005791|Aphereses
C0005791|Blood Component Removal
C0005791|Blood Component Removals
C0005791|Component Removal, Blood
C0005791|Component Removals, Blood
C0005791|Phereses
C0005791|Removal, Blood Component
C0005791|Removals, Blood Component
C0005791|Apheresis (procedure)
C0005791|Apheresis
C0005791|Apheresis.therapeutic
C0005791|Therapeutic apheresis (procedure)
C0005791|Therapeutic apheresis
C0005791|Pheresis
C0005791|Collection, Apheresis/Leukapheresis
C0005791|Apheresis NOS
C0005791|Hemapheresis
C0005791|Apheresis procedure
C0005791|Apheresis - action (qualifier value)
C0005791|Apheresis - action
C0005791|Therapeutic apheresis, NOS
C0206373|Photopheresis
C0206373|Extracorporeal Photochemotherapies
C0206373|Photochemotherapies, Extracorporeal
C0206373|Photopheresis, Extracorporeal
C0206373|extracorporeal photophoresis
C0206373|EXTRACORPOREAL PHOTOCHEMOTHER
C0206373|PHOTOCHEMOTHER EXTRACORPOREAL
C0206373|Extracorporeal Photopheresis
C0206373|photopheresis (treatment)
C0206373|Photophoresis
C0206373|Therapeutc photopheresis
C0206373|PHOTOPHERESIS EXTRACORPOREAL
C0206373|Extracorporeal Photochemotherapy
C0206373|Photochemotherapy, Extracorporeal
C0206373|Extracorporeal photopheresis (procedure)
C0206373|Therapeutic photopheresis
C1879316|Transfusion
C1879316|Transfusion (procedure)
C1879316|transfusions
C1879316|transfusions (treatment)
C1879316|Transfusion, NOS
C0852255|Blood and blood product treatment
C4049189|Immunoadsorption therapy
