C3828565|PHQ-9: total score
C1718207|PHQ-9 interpretation
C4283755|Patient Health Questionnaire Nine Item score
C1718917|Patient Health Questionnaire PHQ-9 administration
C4083201|Patient Health Questionnaire 9 Item
C3641315|PHQ-9 Questionnaire Question
C1715519|Patient health questionnaire 9 item total score:Score:Pt:^Patient:Qn:Reported.PHQ
C3828565|PHQ01-Total Score
C3828565|PHQ-9 - Total Score
C3828565|PHQ0111
C3828565|questionnaires phq-9 total score
C3828565|PHQ-9: total score
C3828565|PHQ-9: total score (procedure)
C1976603|PHQ-9 quick depression assessment panel
C1976603|questionnaires phq-9 quick depression assessment panel
C1976603|PHQ-9: quick depression assessment panel (procedure)
C1976603|PHQ-9: quick depression assessment panel
C3641512|PHQ-9 - Feeling Down, Depressed, or Hopeless
C3641512|PHQ01-Feeling Down Depressed or Hopeless
C3641512|PHQ0102
C3641518|PHQ-9 - Moving or Speaking Slowly or the Opposite being Fidgety or Restless
C3641518|PHQ01-Moving Slowly or Fidgety/Restless
C3641518|PHQ0108
C3641514|PHQ-9 - Feeling Tired or Having Little Energy
C3641514|PHQ0104
C3641514|PHQ01-Feeling Tired or Little Energy
C3641515|PHQ-9 - Poor Appetite or Overeating
C3641515|PHQ0105
C3641515|PHQ01-Poor Appetite or Overeating
C3641516|PHQ-9 - Feeling Bad About Yourself
C3641516|PHQ01-Feeling Bad About Yourself
C3641516|PHQ0106
C3641511|PHQ-9 - Little Interest or Pleasure in Doing Things
C3641511|PHQ0101
C3641511|PHQ01-Little Interest/Pleasure in Things
C3641520|PHQ01-Difficult to Work/Take Care Things
C3641520|PHQ-9 - How Difficult have Problems Made it for You to Work, Take Care of Things, or Get Along with Other People
C3641520|PHQ0110
C3641519|PHQ-9 - Thoughts That You Would be Better Off Dead
C3641519|PHQ01-Thoughts You Be Better Off Dead
C3641519|PHQ0109
C3641513|PHQ-9 - Trouble Falling or Staying Asleep, or Sleeping Too Much
C3641513|PHQ01-Trouble Falling or Staying Asleep
C3641513|PHQ0103
C3641517|PHQ-9 - Trouble Concentrating on Things
C3641517|PHQ01-Trouble Concentrating on Things
C3641517|PHQ0107
C1715519|Patient Health Questionnaire 9 item (PHQ-9) total score [Reported]
C1715519|Patient health questionnaire 9 item total score:Score:Point in time:^Patient:Quantitative:Reported.PHQ
C1715519|Patient health questionnaire 9 item total score:Score:Pt:^Patient:Qn:Reported.PHQ
