C0333106|Bleeding varices
C3837381|gastric variceal procedures
C4288030|Variceal Banding
C0192331|Ligation of esophageal varices
C0192558|Stapling of gastric varices
C0852804|Oesophageal variceal injection
C1739112|Gastrooesophageal variceal haemorrhage prophylaxis
C2062316|acute bleeding of esophageal varices
C2065631|esophagoscopy rigid variceal sclerotherapy
C2960232|Banding of varix of stomach
C3837654|esophagus variceal surgery
C3888799|Gastric variceal injection
C3888800|Gastric variceal ligation
C4272078|Sugiura variceal procedure
C3694764|esophagoscopy transoral flexible with variceal sclerotherapy
C0547715|Follow protocol for vasopressin or nitroglycerine therapy of variceal hemorrhage
C0333106|Bleeding varicose vein
C0333106|Varicose vein hemorrhage
C0333106|Varicose vein haemorrhage
C0333106|Bleeding varices
C0333106|Bleeding varices (morphologic abnormality)
C3837379|gastric surgery variceal stapling (treatment)
C3837379|gastric surgery variceal stapling
C2960232|Banding of varix of stomach (procedure)
C2960232|Banding of gastric varices
C2960232|Banding of varix of stomach
C2960232|gastric surgery variceal banding
C2960232|Banding of gastric varices (treatment)
C3837380|gastric surgery variceal ligation
C3837380|gastric surgery variceal ligation (treatment)
C0192331|ligation of esophageal varices (treatment)
C0192331|ligation of esophageal varices
C0192331|Oesophageal variceal ligation
C0192331|Ligation esoph varix
C0192331|Local ligation of oesophageal varices (procedure)
C0192331|Local ligation of esophageal varices
C0192331|Local ligation of oesophageal varices
C0192331|Ligation of oesophageal varices
C0192331|Esophageal variceal ligation
C0192331|Ligation of esophageal varices (procedure)
C0372009|Ligation, direct, esophageal varices
C0372009|LIGATION DIRECT ESOPHAGEAL VARICES
C0372009|Direct ligation of esophageal varices
C0372009|LIGATE ESOPHAGUS VEINS
C0852804|Oesophageal variceal injection
C0852804|Esophageal variceal injection
C0852804|Injection of esophageal varices
C0852804|Injection of oesophageal varices
C1739112|Gastrooesophageal variceal haemorrhage prophylaxis
C1739112|Gastrooesophageal variceal hemorrhage prophylaxis
C1739112|Gastroesophageal variceal hemorrhage prophylaxis
C1739112|Prophylaxis of gastrooesophageal variceal bleeding
C1739112|Prophylaxis of gastroesophageal variceal bleeding
C0472988|Endoscopic injection sclerotherapy to varices of esophagus using rigid esophagoscope
C0472988|Endoscopic injection sclerotherapy to varices of oesophagus using rigid oesophagoscope
C0472988|Rigid esophagoscopy and injection sclerotherapy of varices
C0472988|Rigid oesophagoscopy and injection sclerotherapy of varices
C0472988|Rigid esophagoscopy and injection sclerotherapy of varices (procedure)
C2959927|Oesophagogastroduodenoscopy and banding of gastric varices
C2959927|Endoscopy of upper gastrointestinal tract and banding of varix of stomach
C2959927|Endoscopy of upper gastrointestinal tract and banding of gastric varices
C2959927|Endoscopy of upper gastrointestinal tract and banding of varix of stomach (procedure)
C2959927|Esophagogastroduodenoscopy and banding of gastric varices
C0472950|Oesoph. varices opn.
C0472950|Operation on oesophageal varices
C0472950|Varices - oesoph.- opn.
C0472950|Operation on esophageal varices
C0472950|Operation on esophageal varices (procedure)
C3888799|Gastric variceal injection
C3888800|Gastric variceal ligation
