C0193388|Biopsy of liver (procedure)
C3174660|Pathology biopsy report:Find:Pt:Liver:Nar
C1524299|Guidance for biopsy:Find:Pt:Abdomen>Liver:Doc:RF
C1628488|CT and biopsy of liver
C1635159|US scan and biopsy of liver
C1955790|Transjugular biopsy of liver
C1955791|Transvenous liver biopsy
C2021366|liver biopsy iron (ug/100 mg of dry weight)
C3836930|liver biopsy with fluoroscopic guidance
C3863012|liver biopsy, transjugular approach
C3880782|Liver biopsy procedure kit
C0193388|Biopsy of liver (procedure)
C0193388|Biopsy of liver
C0193388|Liver biopsy
C0193390|Wedge biopsy of liver
C0521264|Laparoscopic biopsy of liver
C0558534|Percutaneous liver biopsy
C0581276|Needle biopsy of liver
C0842769|Percutaneous [closed] liver biopsy
C0860886|Ultrasound guided liver biopsy
C1261294|Percutaneous needle biopsy liver
C1548877|Consent Type - Liver Biopsy
C1955790|Transjugular biopsy of liver
C1955791|Transvenous liver biopsy
C3522275|Exploration for congenital atresia of bile duct with liver biopsy
C3550399|Increased iron deposition seen on liver biopsy
C0860886|Ultrasound guided liver biopsy
C0372191|Biopsy of liver, needle; when done for indicated purpose at time of other major procedure (List separately in addition to code for primary procedure)
C0372191|NEEDLE BIOPSY LIVER ADD-ON
C0372191|BX LVR NDL DONE PURPOSE TM OTH MAJOR PX
C0176879|Closed liver biopsy
C0176879|Closed (percutaneous) [needle] biopsy of liver
C1955790|Transjugular liver biopsy
C1955790|Transjugular biopsy of liver (procedure)
C1955790|Transjugular biopsy of liver
C1955790|Transjugular liver bx
C2314979|Transjugular biopsy of liver using fluoroscopic guidance
C2314979|Transjugular biopsy of liver using fluoroscopic guidance (procedure)
C0193388|Biopsy of liver
C0193388|Liver Biopsy
C0193388|liver biopsy (procedure)
C0193388|Biopsy liver
C0193388|Biopsy of liver (procedure)
C0193388|Biopsy of liver, NOS
C2121176|a liver biopsy when done for indicated purpose at time of other major procedure
C2121176|liver biopsy when done for indicated purpose at time of other major procedure
C2121176|liver biopsy when done for indicated purpose at time of other major procedure (procedure)
C2021366|liver biopsy iron (ug/100 mg of dry weight) (procedure)
C2021366|liver biopsy iron (ug/100 mg of dry weight)
C2021366|liver biopsy iron
C1261294|Biopsy of liver, needle; percutaneous
C1261294|Percutaneous needle biopsy liver
C1261294|Percutaneous needle biopsy of liver
C1261294|Percutaneous needle biopsy liver (procedure)
C1261294|Percutaneous needle biopsy of liver (procedure)
C1261294|percutaneous needle liver biopsy (procedure)
C1261294|percutaneous needle liver biopsy
C1261294|BIOPSY LIVER NEEDLE PERCUTANEOUS
C1261294|Needle biopsy of liver, accessed through the skin
C1261294|NEEDLE BIOPSY OF LIVER
C0193390|Biopsy of liver, wedge
C0193390|Wedge Biopsy of Liver
C0193390|wedge liver biopsy
C0193390|wedge liver biopsy (procedure)
C0193390|BIOPSY LIVER WEDGE
C0193390|Wedge biopsy of liver (procedure)
C2368137|aspiration of hepatic cyst (procedure)
C2368137|aspiration of hepatic cyst
C0193393|Percutaneous core needle biopsy of liver
C0193393|Percutaneous core needle biopsy of liver (procedure)
C0193389|Open liver biopsy
C0193389|Open biopsy of liver
C0193389|Open biopsy of liver (procedure)
C0193394|Percutaneous fine needle biopsy of liver
C0193394|Percutaneous fine needle aspiration biopsy of liver
C0193394|Percutaneous fine needle biopsy of liver (procedure)
C0581276|Needle Biopsy of Liver
C0581276|Biopsy of liver, needle
C0581276|Needle biopsy of liver (procedure)
C0521264|Laparoscopic liver biopsy
C0521264|Laparoscopic liver bx
C0521264|Laparoscopic biopsy of liver (procedure)
C0521264|Laparoscopic biopsy of liver
C0521264|Laparoscopic biopsy of liver, NOS
C0400397|Diagnostic endoscopic examination of liver and biopsy of lesion of liver using laparoscope
C0400397|Diagnostic endoscopic examination of liver and biopsy of lesion of liver using laparoscope (procedure)
C0400418|Biopsy of liver NEC (procedure)
C0400418|Biopsy of liver NEC
C3836930|liver biopsy with fluoroscopic guidance
C3836930|liver biopsy with fluoroscopic guidance (procedure)
C3863012|liver biopsy, transjugular approach
C3863012|liver biopsy transjugular approach
C3863012|liver biopsy, transjugular approach (procedure)
C4031824|biopsy liver location (procedure)
C4031824|biopsy liver location
C4031823|biopsy liver specimen no. ______
C4031823|biopsy liver specimen no. ______ (procedure)
C4030893|biopsy of liver malignant neoplasm (procedure)
C4030893|biopsy of liver malignant neoplasm
C4030863|biopsy of liver showed carcinoma in situ
C4030863|biopsy of liver showed carcinoma in situ (procedure)
C4030863|bx liver showed carcinoma in situ
C4030881|biopsy of liver showed benign neoplasm
C4030881|biopsy of liver showed benign neoplasm (procedure)
C0400419|Biopsy of liver lesion
C0400419|Biopsy of liver lesion (procedure)
C0558534|Percutaneous Liver Biopsy
C0558534|Percutaneous liver biopsy (procedure)
C0558560|Surgical biopsy of liver (procedure)
C0558560|Surgical biopsy of liver
C0558560|Liver: surgical biopsy (procedure)
C0558560|Liver: surgical biopsy
C1628488|CT and biopsy of liver
C1628488|Computed tomography and biopsy of liver (procedure)
C1628488|Computed tomography and biopsy of liver
C1635159|US scan and biopsy of liver
C1635159|Ultrasound scan and biopsy of liver (procedure)
C1635159|Ultrasound scan and biopsy of liver
C0193392|Open fine needle biopsy of liver (procedure)
C0193392|Open fine needle biopsy of liver
C0193392|Open fine needle aspiration biopsy of liver
C0193392|Open fine needle aspiration biopsy of liver (procedure)
C0193392|Open fine needle biopsy of liver (procedure) [Ambiguous]
C3174660|Pathology biopsy report:Find:Pt:Liver:Nar
C3174660|Liver Path Bx report
C3174660|Pathology biopsy report:Finding:Point in time:Liver:Narrative
C3174660|Liver Pathology biopsy report
C1524299|Fluoroscopy Guidance for biopsy of Liver
C1524299|Liver Flr Bx guid
C1524299|Guidance for biopsy:Finding:Point in time:Liver:Document:XR.fluor
C1524299|Guidance for biopsy:Find:Pt:Liver:Doc:XR.fluor
C2585711|Biopsy of liver using ultrasound guidance (procedure)
C2585711|Biopsy of liver using ultrasound guidance
C1960013|Endoscopic ultrasound examination of liver and biopsy of lesion of liver (procedure)
C1960013|Endoscopic ultrasound examination of liver and biopsy of lesion of liver
C3863011|liver biopsy transjugular approach with fluoroscopic guidance
C3863011|liver biopsy, transjugular approach with fluoroscopic guidance (procedure)
C3863011|liver biopsy, transjugular approach with fluoroscopic guidance
C0400423|Open wedge biopsy of lesion of liver
C0400423|Open wedge biopsy of lesion of liver (procedure)
C0585492|Laparoscopic biopsy of liver lesion
C0585492|Laparoscopic biopsy of liver lesion (procedure)
C2315061|Percutaneous transjugular biopsy of liver using fluoroscopic guidance (procedure)
C2315061|Percutaneous transjugular biopsy of liver using fluoroscopic guidance
C2733386|Percutaneous biopsy of liver using ultrasound guidance (procedure)
C2733386|Percutaneous biopsy of liver using ultrasound guidance
C0400422|Percutaneous transvascular biopsy of lesion of liver
C0400422|Percutaneous transvascular biopsy of lesion of liver (procedure)
C2317400|Fine needle aspiration biopsy of liver
C2317400|Fine needle aspiraton biopsy of liver
C2317400|Fine needle aspiration biopsy of liver (procedure)
C2317400|Fine needle aspiraton biopsy of liver (procedure)
C0554070|Needle biopsy of liver NEC
C0554070|Needle biopsy of liver NEC (procedure)
C0193391|Open core needle biopsy of liver
C0193391|Open core needle biopsy of liver (procedure)
C0554069|Menghini needle biopsy of liver
C0554069|Menghini needle biopsy of liver (procedure)
C0554071|Sheeba needle biopsy of liver
C0554071|Sheeba needle biopsy of liver (procedure)
C2732498|Percutaneous needle biopsy of liver using fluoroscopic guidance (procedure)
C2732498|Percutaneous needle biopsy of liver using fluoroscopic guidance
C3836502|percutaneous needle liver biopsy with fluoroscopic guidance
C3836502|percutaneous needle liver biopsy with fluoroscopic guidance (procedure)
C3862599|percutaneous needle liver biopsy fine needle aspiration (procedure)
C3862599|percutaneous needle liver biopsy fine needle aspiration
