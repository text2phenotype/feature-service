Anatomy|abdomen|abdom||abdominal|
Anatomy|abdomen|lapar||laparoscopic|
Anatomy|arm|brachi||brachial|
Anatomy|artery|aort/o||aortography|aorta
Anatomy|artery|arteri/o||arteriostenosis|artery
Anatomy|back|dors||dorsalgia|
Anatomy|bladder|vesic||vesicular|
Anatomy|blood|angi/o||angiorrhexis|blood vessels
Anatomy|blood|sangui|||
Anatomy|blood|hemat||hematometra|
Anatomy|blood|haemat||haematemesis|
Anatomy|blood_vessel|vas||vascular|
Anatomy|blood_vessel|vascul||vascular|
Anatomy|body|somat|||
Anatomy|body|som|||
Anatomy|bone|oste||osteoporosis|
Anatomy|bone|ossi||ossification|
Anatomy|brain|encephal||encephalopathy|
Anatomy|brain|cerebr||cerebral|
Anatomy|breast|mast||mastectomy|
Anatomy|breast|mamm/o||mammogram|
Anatomy|cells||blast|osteoblast|embryonic, immature
Anatomy|cells||cyte|hematocyte|cell
Anatomy|cells||cytes|lymphocytes|cells
Anatomy|chest||thorax|hemothorax|chest, pleural cavity
Anatomy|chest|steth||stethoscopes|
Anatomy|chest|pector||pectoris|
Anatomy|colorectal|proct||proctology|anus, rectum
Anatomy|colorectal|rect||rectum|rectal, rectum
Anatomy|cyst|cyst||cystoid|
Anatomy|digit|dactyl|||
Anatomy|digit|digit||| 
Anatomy|ear|tympan/o||tympanocentesis|drum, eardrum
Anatomy|ear||cusis|paracusis|hearing
Anatomy|eye|irid||iridectomy|
Anatomy|eye|opthalm/o||opthalmologist|
Anatomy|eye|optic/o||opticochemical|
Anatomy|eye|ocul/o||oculocerebrorenal|
Anatomy|fat|lip/o||lipomatosis|
Anatomy|fat|adip/o||adipose|
Anatomy|fat|ather/o||atherosclerosis|
Anatomy|gallbladder|cholecyst/o||cholecystography|
Anatomy|gland||crine|endocrine|
Anatomy|gland|adren||adrenal|
Anatomy|gland|adreno||Adrenochrome|
Anatomy|gland|aden/o||adenocarcinoma| 
Anatomy|gland|hormon||hormone|hormone
Anatomy|glucose|gluc||glucose|sugar
Anatomy|hand|cheir||| 
Anatomy|hand|manu||| 
Anatomy|hand|chir||| 
Anatomy|head|cephal/o||cephalometry| 
Anatomy|heart|cardi||cardiogram|
Anatomy|heart|cordi||| 
Anatomy|heart||cardium|myocardium|
Anatomy|heart|myocard||myocardial|heart
Anatomy|intenstine|entero|||
Anatomy|joint|arthr||arthritis|
Anatomy|joint|articul||articulate|
Anatomy|kidney|nephr/o||nephrosclerosis|
Anatomy|liver|hepat/o||hepatocellular|liver
Anatomy|liver|hepatic|||
Anatomy|lumb|lumb||lumbar|trunk between lowest ribs +pelvis
Anatomy|lung|pneumon||pneumonia|
Anatomy|lung|pulmo/n||pulmonary|
Anatomy|lung|alveol/o||alveolar|alveolus, small sac
Anatomy|lung|bronchi/o||bronchiectasis|airways
Anatomy|lymph|lymph||lymphedema|
Anatomy|marrow|myel||myelofibrosis|
Anatomy|marrow|medull||medulla|
Anatomy|mind|ment||| 
Anatomy|mouth|stomat/o|||
Anatomy|muscle|muscul||musculoskeletal|
Anatomy|muscle|myo||myoclonic|
Anatomy|neck|trachel/o|||
Anatomy|neck|cervic|||confuses with cervical (cancer)
Anatomy|nerve|neur/o||neurogenic|
Anatomy|nerve|nerv||nerves|
Anatomy|pelvis|pelv||pelvis|
Anatomy|psych|psych||psychiatry|SEE Anatomy.brain
Anatomy|shoulder|humer||humeral|
Anatomy|sinus|sinus||sinusitis|
Anatomy|skin|dermat/o||dermatoglyphics|
Anatomy|skin|derm||dermabrasion|
Anatomy|skin|cuticul||cuticularia|
Anatomy|skull|crani/o||craniometry|
Anatomy|sperm|sperm||spermatogenesis|sperm, male reproduction
Anatomy|stomach|gastr/o||gastrointestinal|
Anatomy|stomach|ventr/o||| 
Anatomy|testis|orchi|||
Anatomy|throat|trache||trachea|
Anatomy|throat|pharyng||pharyngitis|
Anatomy|thumb|pollic||pollichia|
Anatomy|tissue|histol||histology|tissue
Anatomy|tissue|histi/o||histiocytoma|tissue
Anatomy|tongue|gloss||| 
Anatomy|tongue|glott||| 
Anatomy|tongue|lingu/a||| 
Anatomy|tooth|odont/o||odontogenesis|
Anatomy|tooth|dent||dental|
Anatomy|tumor|cel||| 
Anatomy|tumor|onco||oncology| 
Anatomy|tumor|tum||tumor|
Anatomy|urinary|urethr/a||urethral|
Anatomy|urinary|urin||urine|
Anatomy|uterus|hyster/o||hysterotomy|
Anatomy|uterus|metr/o||| 
Anatomy|uterus|uter||uterine|
Anatomy|vein|ven|||veins, venous blood, vascular system
Anatomy|ventricle|ventricul||ventriculography|
Anatomy|wrist|carp/o|||