C0014544|Epilepsy
C0751495|partial seizure
C0751495|Focal Seizure
C0751495|Seizures, partial, afebrile
C0751495|partial seizure (physical finding)
C0751495|seizure partial (focal)
C0751495|Convulsions local
C0751495|Partial seizures, NOS
C0751495|Focal Seizures
C0751495|Seizure, Focal
C0751495|Seizures, partial
C0751495|Partial seizures
C0751495|Local convulsion
C0751495|Partial seizure (finding)
C0751495|Local convulsion (disorder)
C0751495|Seizures, focal
C0751495|Partial seizures NOS
C0751495|Focal fits
C0751495|Local seizure
C0751495|Partial seizure (disorder)
C0751495|Focal seizure, NOS
C0234533|generalized seizure
C0234533|Generalized seizures
C0234533|generalized convulsions (symptom)
C0234533|generalized convulsions
C0234533|generalized seizure (physical finding)
C0234533|seizure generalized
C0234533|Seizure, Generalized
C0234533|Seizures, generalized
C0234533|Generalized convulsion
C0234533|Generalised convulsion
C0234533|Generalized convulsion (finding)
C0234533|Convulsions generalized
C0234533|Convulsions generalised
C0234533|Generalised seizure
C0234533|Generalised fit
C0234533|Generalized fit
C0234533|Generalized seizure (finding)
C0234533|convulsions; generalized
C0234533|generalized; convulsions
C0234533|Generalized convulsion, NOS
C0014544|Epilepsies
C0014544|Epilepsy
C0014544|Epilepsy, unspecified
C0014544|Epileptic Seizure
C0014544|Seizure, Epileptic
C0014544|Seizure disorder NOS
C0014544|Seizure disorder
C0014544|SEIZURE DIS
C0014544|epilepsia
C0014544|epilepsy (diagnosis)
C0014544|seizure disorder (diagnosis)
C0014544|Seizure Disorders
C0014544|Epileptic convulsions NOS
C0014544|Epileptic fits NOS
C0014544|Epilepsy NOS
C0014544|Epileptic seizures NOS
C0014544|Epilepsy [Disease/Finding]
C0014544|Epileptic Seizures
C0014544|Seizures, Epileptic
C0014544|Seizure;epileptic
C0014544|Epileptic attack
C0014544|Epilepsy NOS (disorder)
C0014544|(Epilepsy) or (epileptic attack) (disorder)
C0014544|(Epilepsy) or (epileptic attack)
C0014544|Attack - epileptic
C0014544|Epileptic fit
C0014544|EF - Epileptic fit
C0014544|EP - Epilepsy
C0014544|Epileptic
C0014544|Epilepsy (disorder)
C0014544|Epileptic convulsions
C0014544|Epileptic disorder
C0014544|Epileptic fits
C0014544|Epileptic seizure (finding)
C0014544|Seizure disorder (disorder)
C0014544|caducus; morbus
C0014544|cerebral; epileptic
C0014544|convulsions; epileptic
C0014544|epilepsy; cerebral
C0014544|epilepsy; cortical
C0014544|epilepsy; fit
C0014544|epilepsy; seizure
C0014544|epileptic; convulsions
C0014544|epileptic; syndrome
C0014544|fit; epileptic
C0014544|morbus; caducus
C0014544|seizure; epileptic
C0014544|syndrome; epileptic
C0014544|Epilectic attack, NOS
C0014544|Epilepsy, NOS
C0014544|Epileptic convulsions, NOS
C0014544|Epileptic disorder, NOS
C0014544|Epileptic fits, NOS
C0014544|Epileptic seizures, NOS
C0014544|Epileptic attack, NOS
C0270850|Generalized idiopathic epilepsy and epileptic syndromes
C0270850|IGE
C0270850|EIG
C0270850|EPILEPSY, IDIOPATHIC GENERALIZED
C0270850|Idiopathic generalized epilepsy
C0270850|Generalized idiopathic epilepsy and epileptic syndromes NOS
C0270850|Idiopathic generalised epilepsy
C0270850|epilepsy generalized idiopathic
C0270850|epilepsy generalized idiopathic (diagnosis)
C0270850|Primary generalised epilepsy
C0270850|Primary generalized epilepsy
C0270850|Idiopathic generalized epilepsy (disorder)
C0270850|epilepsy; generalized, idiopathic
C0270850|epilepsy; idiopathic, generalized
C0270850|epilepsy; syndrome, generalized, idiopathic
C0270850|generalized; epileptic, idiopathic
C0270850|syndrome; epileptic, generalized, idiopathic
C0270850|Idiopathic generalized epilepsy, NOS
C0494475|Grand mal seizures, unspecified (with or without petit mal)
C0494475|Generalized Tonic-Clonic Seizure
C0494475|Grand Mal Seizure
C0494475|Grand Mal
C0494475|Grand-Mal Seizure
C0494475|Generalized tonic clonic seizures
C0494475|Generalized tonic-clonic seizures
C0494475|Seizures, generalized tonic-clonic
C0494475|Generalized clonic-tonic seizures
C0494475|Seizures, tonic-clonic
C0494475|Generalized tonic-clonic seizures (GTCS)
C0494475|Generalised tonic-clonic seizures
C0494475|Seizure, Tonic-Clonic
C0494475|Seizures, Tonic Clonic
C0494475|Tonic-Clonic Seizure
C0494475|Tonic-Clonic Seizures
C0494475|Seizures, clonic-tonic
C0494475|Seizure;tonic-clonic
C0494475|Grand mal seizures
C0494475|Grand mal seizure NOS
C0494475|Seizures, generalized tonic-clonic (GTCS)
C0494475|Grand mal seizure (disorder)
C0494475|Grand mal convulsion
C0494475|Grand mal seizure (finding)
C0494475|Generalised tonic-clonic seizure
C0494475|Seizures, Grand-Mal
C0494475|Grand-Mal Seizures
C0494475|Seizures, generalized, tonic-clonic
C0494475|Grand mal epileptic fit
C0494475|Grand mal fit
C0494475|Seizure grand mal
C0494475|tonic-clonic seizure (physical finding)
C0494475|seizure generalized tonic-clonic
C0494475|tonic-clonic convulsion
C0494475|tonic-clonic convulsions
C0494475|Tonic-clonic seizure (finding)
C0494475|Tonic - clonic seizures
C0494475|grand mal; seizure
C0494475|haut mal
C0494475|seizure; grand mal
C0475521|Localization-related (focal) (partial) idiopathic epilepsy and epileptic syndromes with seizures of localized onset
C0475521|Localization-related (focal) (partial) idiopathic epilepsy and epileptic syndromes with seizures of localized onset NOS
C0475521|Localization-related(focal)(partial)idiopathic epilepsy and epileptic syndromes with seizures of localised onset
C0475521|Localization-related(focal)(partial)idiopathic epilepsy and epileptic syndromes with seizures of localized onset
C0475521|Localization-related(focal)(partial)idiopathic epilepsy and epileptic syndromes with seizures of localized onset (disorder)
C0494472|Localization-related (focal) (partial) symptomatic epilepsy and epileptic syndromes with complex partial seizures
C0494472|Localization-related (focal) (partial) symptomatic epilepsy and epileptic syndromes with complex partial seizures NOS
C0494471|Localization-related (focal) (partial) symptomatic epilepsy and epileptic syndromes with simple partial seizures
C0494471|Localization-related (focal) (partial) symptomatic epilepsy and epileptic syndromes with simple partial seizures NOS
C0477371|Other forms of epilepsy
C0477371|Other epilepsy
C0477371|Other epilepsy NOS
C0477371|Other forms of epilepsy NOS (disorder)
C0477371|Other forms of epilepsy (disorder)
C0477371|Other forms of epilepsy NOS
C0477371|[X]Other epilepsy
C0477371|[X]Other epilepsy (disorder)
C0477370|Other generalized epilepsy and epileptic syndromes
C0477370|Other generalized epilepsy and epileptic syndromes NOS
C0477370|[X]Other generalized epilepsy and epileptic syndromes (disorder)
C0477370|[X]Other generalized epilepsy and epileptic syndromes
C0477370|[X]Other generalised epilepsy and epileptic syndromes
C0477370|syndrome; epileptic, generalized
C0014553|Absence Epilepsy
C0014553|Epilepsy, Absence
C0014553|Petit Mal Epilepsies
C0014553|Pyknolepsies
C0014553|Seizure, Absence
C0014553|Absence Seizure
C0014553|Absence seizures
C0014553|Petit mal, unspecified, without grand mal seizures
C0014553|Petit Mal Seizure
C0014553|Petit Mal
C0014553|Petit-Mal Seizure
C0014553|Seizures, absence
C0014553|ABSENCE SEIZURE DIS
C0014553|SEIZURE DIS ABSENCE
C0014553|pyknolepsy
C0014553|epilepsy generalized nonconvulsive pykno-epilepsy (diagnosis)
C0014553|epilepsy generalized nonconvulsive pykno-epilepsy
C0014553|generalized nonconvulsive petit mal seizure
C0014553|petit mal seizure (diagnosis)
C0014553|pykno-epilepsy
C0014553|Petit mal epilepsy
C0014553|Absence Seizure Disorders
C0014553|Seizure Disorders, Absence
C0014553|Convulsion, Petit Mal
C0014553|Minor Epilepsies
C0014553|Minor Epilepsy
C0014553|Pykno Epilepsy
C0014553|Pykno-Epilepsies
C0014553|Childhood absence seizures
C0014553|Epilepsy, Minor
C0014553|Epilepsy, Absence [Disease/Finding]
C0014553|Juvenile Absence Epilepsy
C0014553|Childhood Absence Epilepsy
C0014553|Absence Seizure Disorder
C0014553|Epilepsy, Petit Mal
C0014553|Petit Mal Convulsion
C0014553|Seizure Disorder, Absence
C0014553|Seizure;absence
C0014553|Typical absence seizure
C0014553|Typical absence seizure (disorder)
C0014553|Epilepsy Juvenile Absences
C0014553|Juvenile Absences, Epilepsy
C0014553|Juvenile Absence, Epilepsy
C0014553|Juvenile absence epilepsy (disorder)
C0014553|Absence seizure (finding)
C0014553|Childhood absence epilepsy (disorder)
C0014553|Petit mal (disorder)
C0014553|Epilepsy Juvenile Absence
C0014553|Petit-Mal Seizures
C0014553|Seizures, Petit-Mal
C0014553|Petit mal seizures
C0014553|Typical absence seizures
C0014553|Convulsion petit mal
C0014553|Epilepsy petit mal
C0014553|seizure generalized absence
C0014553|absence seizure (physical finding)
C0014553|childhood absence seizure (diagnosis)
C0014553|juvenile absence seizure (diagnosis)
C0014553|juvenile absence seizure
C0014553|childhood absence seizure
C0014553|Childhood - juvenile - absence epilepsy
C0014553|Petit-mal epilepsy
C0014553|Absence seizure (disorder)
C0014553|epilepsy; absence
C0014553|epilepsy; minor
C0014553|epilepsy; petit mal
C0014553|absence; epileptic
C0014553|absences; epileptic
C0014553|petit mal; epilepsy
C0014553|Absence Epilepsies, Childhood
C0014553|Absence Epilepsy, Childhood
C0014553|Childhood Absence Epilepsies
C0014553|Epilepsies, Childhood Absence
C0014553|Epilepsy, Childhood Absence
C0014553|Absence Epilepsies, Juvenile
C0014553|Absence Epilepsy, Juvenile
C0014553|Epilepsies, Juvenile Absence
C0014553|Epilepsy, Juvenile Absence
C0014553|Juvenile Absence Epilepsies
C0014553|Absences, typical
C0014553|absence of seizure
C0494474|Special epileptic syndromes
C0494474|epilepsy; syndrome, special
C0494474|epileptic; syndrome, special
C0494474|syndrome; epileptic, special
C0009952|Febrile convulsion
C0009952|Convulsion, Febrile
C0009952|Febrile Convulsions
C0009952|Febrile Seizure
C0009952|Seizures, Febrile
C0009952|Seizure, Febrile
C0009952|Febrile convulsions (simple), unspecified
C0009952|Febrile seizures NOS
C0009952|[D]Convulsions, febrile (context-dependent category)
C0009952|Seizures, generalized, associated with fever
C0009952|Seizures, febrile, in early childhood
C0009952|Febrile seizures
C0009952|febrile convulsion (diagnosis)
C0009952|Febrile Convulsion Seizures
C0009952|Seizure, Febrile Convulsion
C0009952|Seizures, Febrile Convulsion
C0009952|Convulsion, Fever
C0009952|Convulsions, Fever
C0009952|Fever Convulsions
C0009952|Convulsion, Pyrexial
C0009952|Convulsions, Pyrexial
C0009952|Pyrexial Convulsions
C0009952|Febrile Fits
C0009952|Fit, Febrile
C0009952|Fits, Febrile
C0009952|Fever Seizures
C0009952|Seizure, Fever
C0009952|Seizures, Fever
C0009952|Pyrexial Seizures
C0009952|Seizure, Pyrexial
C0009952|Seizures, Pyrexial
C0009952|Febrile convulsions NOS
C0009952|Febrile seizure NOS
C0009952|Febrile convulsion NOS
C0009952|Febrile Fit
C0009952|Fever Seizure
C0009952|Pyrexial Seizure
C0009952|Convulsions, Febrile
C0009952|Febrile Convulsion Seizure
C0009952|Seizures, Febrile [Disease/Finding]
C0009952|Fever Convulsion
C0009952|Pyrexial Convulsion
C0009952|Convulsions;febrile
C0009952|Seizure;febrile
C0009952|[D]Convulsions, febrile (situation)
C0009952|[D]Convulsions, febrile
C0009952|Febrile seizure (from fever)
C0009952|[D]Pyrexial convulsion
C0009952|Febrile convulsions (finding)
C0009952|Convulsion febrile
C0009952|Pyrexial fit
C0009952|Febrile convulsion (finding)
C0009952|convulsions; febrile
C0009952|febrile; convulsions
C0009952|febrile; seizures
C0009952|seizure; febrile
C0014547|Epilepsies, Focal
C0014547|Epilepsies, Localization-Related
C0014547|Epilepsies, Partial
C0014547|Focal Epilepsies
C0014547|Focal Epilepsy
C0014547|Localization-Related Epilepsies
C0014547|Localization-Related Epilepsy
C0014547|Partial Epilepsies
C0014547|FOCAL SEIZURE DIS
C0014547|PARTIAL SEIZURE DIS
C0014547|SEIZURE DIS PARTIAL
C0014547|EPILEPSY LOCALIZATION RELAT
C0014547|SEIZURE DIS FOCAL
C0014547|Localization-related epilepsy -RETIRED-
C0014547|Localisation-related epilepsy -RETIRED-
C0014547|Disorders, Focal Seizure
C0014547|Focal Seizure Disorders
C0014547|Seizure Disorders, Focal
C0014547|Disorders, Partial Seizure
C0014547|Partial Seizure Disorders
C0014547|Seizure Disorders, Partial
C0014547|Epilepsies, Partial [Disease/Finding]
C0014547|Epilepsy, Partial
C0014547|Focal Seizure Disorder
C0014547|Seizure Disorder, Focal
C0014547|Epilepsy, Focal
C0014547|Epilepsy, Localization-Related
C0014547|Seizure Disorder, Partial
C0014547|Partial Epilepsy
C0014547|Partial Seizure Disorder
C0014547|Localisation-related epilepsy
C0014547|Localisation-related epilepsy (disorder)
C0014547|Localization-related epilepsy (disorder)
C0014547|Localisation related epilepsy
C0014547|Localization related epilepsy
C0014547|Local epilepsy
C0014547|epilepsy; focal
C0014547|epilepsy; localization-related
C0014547|epilepsy; partial
C0014547|focal; epileptic
C0014547|partial; epileptic
C0014547|Focal epilepsy, NOS
C0014547|Localization-related epilepsy, NOS
C0014547|Epilepsy, focal NOS
C0014547|Epilepsy, partial NOS
C0014548|Epilepsies, Generalized
C0014548|Epilepsy, Generalized
C0014548|Generalized Epilepsies
C0014548|Generalized Epilepsy
C0014548|SEIZURE DIS GENERALIZED
C0014548|Generalized Seizure Disorder
C0014548|Generalized Seizure Disorders
C0014548|Seizure Disorders, Generalized
C0014548|Epilepsy, Generalized [Disease/Finding]
C0014548|Seizure Disorder, Generalized
C0014548|epilepsy generalized
C0014548|generalized epilepsy (diagnosis)
C0014548|Generalised epilepsy (disorder)
C0014548|Generalised epilepsy
C0014548|Generalized epilepsy (disorder)
C0014548|epilepsy; generalized
C0014548|epilepsy; syndrome, generalized
C0014548|generalized; epileptic
C0014548|Generalized epilepsy, NOS
C0014548|Generalised epilepsy [Ambiguous]
C0014550|Epilepsies, Myoclonic
C0014550|Epilepsy, Myoclonic
C0014550|Myoclonic Epilepsies
C0014550|Myoclonus Epilepsies
C0014550|Myoclonus Epilepsy
C0014550|Seizures, myoclonic
C0014550|Myoclonic seizures
C0014550|Myoclonic epilepsy
C0014550|MYOCLONIC SEIZURE DIS
C0014550|myoclonia epileptica
C0014550|myoclonic seizure
C0014550|Myoclonic seizure disorder
C0014550|myoclonic epilepsy (diagnosis)
C0014550|generalized convulsive myoclonic seizure
C0014550|Disorder, Myoclonic Seizure
C0014550|Disorders, Myoclonic Seizure
C0014550|Myoclonic Seizure Disorders
C0014550|Seizure Disorder, Myoclonic
C0014550|Seizure Disorders, Myoclonic
C0014550|Epilepsies, Myoclonic [Disease/Finding]
C0014550|Epilepsy, Myoclonus
C0014550|Seizure;myoclonic
C0014550|Myoclonic seizure NOS
C0014550|seizure generalized myoclonic
C0014550|myoclonic seizure (physical finding)
C0014550|Epileptic seizures - myoclonic
C0014550|Epileptic seizures - myoclonic (disorder)
C0014550|Myoclonic seizure (disorder)
C0014550|epilepsy; myoclonus
C0014550|epileptica; myoclonus
C0014550|Epileptic seizures, myoclonic
C0014557|Epilepsies, Post-Traumatic
C0014557|Epilepsies, Traumatic
C0014557|Epilepsy, Post Traumatic
C0014557|Epilepsy, Post-Traumatic
C0014557|Post-Traumatic Epilepsies
C0014557|Post-Traumatic Epilepsy
C0014557|Traumatic Epilepsies
C0014557|Traumatic Epilepsy
C0014557|SEIZURE DIS POST TRAUMATIC
C0014557|POST TRAUMATIC SEIZURE DIS
C0014557|Disorder, Post-Traumatic Seizure
C0014557|Disorders, Post-Traumatic Seizure
C0014557|Post Traumatic Seizure Disorder
C0014557|Post-Traumatic Seizure Disorders
C0014557|Seizure Disorder, Post Traumatic
C0014557|Seizure Disorders, Post-Traumatic
C0014557|Epilepsy, Post-Traumatic [Disease/Finding]
C0014557|Post-Traumatic Seizure Disorder
C0014557|Epilepsy, Traumatic
C0014557|Seizure Disorder, Post-Traumatic
C0014557|Traumatic epilepsy (disorder)
C0014557|PTE - Post-traumatic epilepsy
C0014557|Post-traumatic epilepsy (disorder)
C0014557|epilepsy; traumatic
C0014557|traumatic; epileptic
C0036572|Seizure
C0036572|Convulsions
C0036572|Seizures
C0036572|convulsion
C0036572|[D]Convulsion NOS (context-dependent category)
C0036572|[D]Convulsions (context-dependent category)
C0036572|[D]Fit (context-dependent category)
C0036572|Seizure NOS
C0036572|seizure (physical finding)
C0036572|convulsions (symptom)
C0036572|Fit, NOS
C0036572|Seizure, NOS
C0036572|Convulsion, NOS
C0036572|Unspecified convulsions
C0036572|Fit NOS
C0036572|Seizures [Disease/Finding]
C0036572|Fit(s)
C0036572|Fits - convulsions
C0036572|[D]Convulsions
C0036572|[D]Convulsions (situation)
C0036572|[D]Fit (situation)
C0036572|[D]Fit
C0036572|[D]Convulsion NOS
C0036572|Fits - convulsions (disorder)
C0036572|[D]Convulsion NOS (situation)
C0036572|[D]Seizure NOS
C0036572|Fit - convulsion (finding)
C0036572|Fit
C0036572|Fit - convulsion
C0036572|Convulsion (disorder)
C0036572|Fitting
C0036572|Convulsion (NOS)
C0036572|Fits NOS
C0036572|Convulsions NOS
C0036572|Seizure (finding)
C0036572|fits
C0038220|Status Epilepticus
C0038220|Status epilepticus, unspecified
C0038220|Generalized Status Epilepticus
C0038220|Status Epilepticus [Disease/Finding]
C0038220|Status Epilepticus, Generalized
C0038220|[X]Status epilepticus, unspecified (disorder)
C0038220|[X]Status epilepticus, unspecified
C0038220|Status epilepticus (disorder)
C0038220|epilepsy; status
C0038220|epilepticus; status
C0038220|status; epilepticus
C0038220|status; epileptic
C0038220|Status epilepticus NOS
C0282512|Acquired Epileptic Aphasia
C0282512|Acquired Epileptic Aphasias
C0282512|Epileptic Aphasia, Acquired
C0282512|Epileptic Aphasias, Acquired
C0282512|Landau Kleffner Syndrome
C0282512|Landau-Kleffner Syndrome
C0282512|Syndrome, Landau-Kleffner
C0282512|Acquired aphasia with epilepsy [Landau-Kleffner]
C0282512|LKS
C0282512|ACQUIRED CHILDHOOD APHASIA WITH CONVULSIVE DIS
C0282512|Acquired Childhoood Aphasia with Convulsive Disorder
C0282512|Aphasia, Epileptic, Acquired
C0282512|Landau-Kleffner Acquired Epileptiform Aphasia
C0282512|Aphasia, Acquired Epileptic
C0282512|Landau-Kleffner Syndrome [Disease/Finding]
C0282512|Acquired Epileptiform Aphasias
C0282512|Epileptiform Aphasias, Acquired
C0282512|Epileptiform Aphasia, Acquired
C0282512|Acquired Aphasia with Convulsive Disorder
C0282512|Acquired Epileptiform Aphasia
C0282512|Landau Kleffner Acquired Epileptiform Aphasia
C0282512|Aphasia, Acquired, With Convulsive Disorder
C0282512|Acquired aphasia with epilepsy
C0282512|Acquired epileptic aphasia (disorder)
C0282512|Acquired epileptic aphasia (diagnosis)
C0282512|developmental disorder - speech acquired epileptic aphasia
C0270857|Epilepsies, Reflex
C0270857|Epilepsy, Reflex
C0270857|Reflex Epilepsies
C0270857|Reflex Epilepsy
C0270857|Epilepsy, Reflex [Disease/Finding]
C0270857|Epilepsy associated with specific stimuli
C0270857|Sensory-induced epilepsy
C0270857|Reflex epilepsy (disorder)
C0270857|epilepsy; reflex
C0270857|Epilepsy, sensory-induced
C0270851|Benign Neonatal Convulsion
C0270851|Convulsion, Benign Neonatal
C0270851|Convulsions, Benign Neonatal
C0270851|Neonatal Convulsion, Benign
C0270851|Benign Neonatal Epilepsies
C0270851|Epilepsies, Benign Neonatal
C0270851|Epilepsy, Benign Neonatal
C0270851|Neonatal Epilepsies, Benign
C0270851|Neonatal Epilepsy, Benign
C0270851|Benign Neonatal Epilepsy
C0270851|Neonatal Convulsions, Benign
C0270851|Benign Neonatal Convulsions
C0270851|Epilepsy, Benign Neonatal [Disease/Finding]
C0270851|Benign neonatal seizures
C0270851|Benign neonatal seizures (disorder)
C0270851|Benign neonatal convulsions (disorder)
C0270851|Benign neonatal seizures [Ambiguous]
C1856931|EPILEPSY, PHOTOGENIC, WITH SPASTIC DIPLEGIA AND MENTAL RETARDATION
C1856930|EPILEPSY WITH BILATERAL OCCIPITAL CALCIFICATIONS
C1856930|Epilepsy occipital calcifications
C1856930|Bilateral occipital calcifications with epilepsy
C1856930|Familial unilateral and bilateral occipital calcifications and epilepsy
C2584947|Anoxic epileptic seizure
C2584947|Anoxic epileptic seizure (finding)
C0270853|juvenile myoclonic epilepsy
C0270853|generalized convulsive myoclonic seizure, juvenile
C0270853|juvenile myoclonic epilepsy (diagnosis)
C0270853|Adolescent Myoclonic Epilepsies
C0270853|Epilepsies, Adolescent Myoclonic
C0270853|Epilepsy, Adolescent Myoclonic
C0270853|Myoclonic Epilepsies, Adolescent
C0270853|Epilepsies, Juvenile Myoclonic
C0270853|Epilepsy, Juvenile Myoclonic
C0270853|Juvenile Myoclonic Epilepsies
C0270853|Myoclonic Epilepsies, Juvenile
C0270853|Myoclonic Epilepsy, Juvenile
C0270853|Syndrome, Janz
C0270853|EJM
C0270853|JME
C0270853|EPILEPSY, MYOCLONIC JUVENILE
C0270853|Adolescent Myoclonic Epilepsy
C0270853|Janz Juvenile Myoclonic Epilepsy
C0270853|Epilepsy, Myoclonic, Juvenile
C0270853|Myoclonic Epilepsy, Juvenile [Disease/Finding]
C0270853|Impulsive Petit Mal, Janz
C0270853|Janz Syndrome
C0270853|Myoclonic Epilepsy, Adolescent
C0270853|Petit Mal, Impulsive, Janz
C0270853|Juvenile Myoclonic Epilepsy of Janz
C0270853|Impulsive Petit Mal Epilepsy
C0270853|JME (Juvenile Myoclonic Epilepsy)
C0270853|Janz Impulsive Petit Mal
C0270853|Petit Mals, Impulsive
C0270853|Myoclonic Epilepsy, Juvenile, 1
C0270853|Petit Mal, Impulsive
C0270853|JMEs (Juvenile Myoclonic Epilepsy)
C0270853|Impulsive petit mal of Janz
C0270853|Impulsive petit-mal epilepsy
C0270853|Myoclonic epilepsy of adolescence
C0270853|JME - Juvenile myoclonic epilepsy
C0270853|Juvenile myoclonic epilepsy (disorder)
C0270853|impulsive; petit mal
C0270853|myoclonic; epileptic, juvenile
C1848137|EFMR
C1848137|EPILEPSY, FEMALE-RESTRICTED, WITH MENTAL RETARDATION (disorder)
C1848137|EPILEPTIC ENCEPHALOPATHY, EARLY INFANTILE, 9
C1848137|EIEE9
C1848137|Convulsive Disorder and Mental Retardation
C1848137|Epilepsy, Female-Restricted, with Mental Retardation
C1848137|JUBERG-HELLMAN SYNDROME
C2875138|Epilepsy, unspecified, not intractable
C2875141|Epilepsy, unspecified, intractable
C2919602|Epileptic seizure witnessed by provider of history other than subject
C2919602|Witnessed epileptic seizure
C2919602|Epileptic seizure witnessed by provider of history other than subject (finding)
C1096063|Intractable epilepsy
C1096063|Refractory epilepsy (disorder)
C1096063|Refractory epilepsy
C1096063|epilepsy intractable
C1096063|epilepsy intractable (diagnosis)
C1096063|Epilepsies, Drug Resistant
C1096063|Intractable Epilepsies
C1096063|Epilepsies, Drug Refractory
C1096063|Resistant Epilepsy, Drug
C1096063|Medication Resistant Epilepsies
C1096063|Resistant Epilepsies, Medication
C1096063|Epilepsy, Medication Resistant
C1096063|Refractory Epilepsy, Drug
C1096063|Drug Resistant Epilepsy
C1096063|Epilepsies, Intractable
C1096063|Drug Resistant Epilepsies
C1096063|Resistant Epilepsies, Drug
C1096063|Epilepsies, Medication Resistant
C1096063|Drug Refractory Epilepsies
C1096063|Resistant Epilepsy, Medication
C1096063|Refractory Epilepsies, Drug
C1096063|Epilepsy, Drug Refractory
C1096063|Epilepsy, Drug Resistant
C1096063|Epilepsy, Intractable
C1096063|Drug Refractory Epilepsy
C1096063|Medication Resistant Epilepsy
C1096063|Drug Resistant Epilepsy [Disease/Finding]
C0017332|Generalized nonconvulsive epilepsy
C0017332|GENERALIZED SEIZURE DIS NONCONVULSIVE
C0017332|NONCONVULSIVE SEIZURE DIS GENERALIZED
C0017332|SEIZURE DIS NONCONVULSIVE GENERALIZED
C0017332|GENERALIZED NONCONVULSIVE SEIZURE DIS
C0017332|NONCONVULSIVE GENERALIZED SEIZURE DIS
C0017332|SEIZURE DIS GENERALIZED NONCONVULSIVE
C0017332|generalized nonconvulsive seizure (diagnosis)
C0017332|generalized nonconvulsive seizure
C0017332|Generalised non-convulsive epilepsy
C0017332|Epilepsy, Generalized Nonconvulsive
C0017332|Nonconvulsive Epilepsy, Generalized
C0017332|Generalized nonconvulsive epilepsy (disorder)
C0017332|Generalised non-convulsive epilepsy NOS
C0017332|Generalized non-convulsive epilepsy NOS
C0017332|Generalized non-convulsive epilepsy NOS (disorder)
C0017332|Generalised nonconvulsive epilepsy
C0017332|Generalized non-convulsive epilepsy
C0017332|Seizure Disorder, Nonconvulsive Generalized
C0017332|Seizure Disorder, Generalized Nonconvulsive
C0017332|Generalized Seizure Disorder, Nonconvulsive
C0017332|Nonconvulsive Generalized Seizure Disorder
C0017332|Nonconvulsive Seizure Disorder, Generalized
C0017332|Generalized non-convulsive epilepsy (disorder)
C0017332|epilepsy; generalized, nonconvulsive
C0017332|generalized; epileptic, nonconvulsive
C0017332|Generalized nonconvulsive epilepsy, NOS
C0017332|Generalized Nonconvulsive Seizure Disorder
C0311334|CONVULSIVE GENERALIZED SEIZURE DIS
C0311334|CONVULSIVE SEIZURE DIS GENERALIZED
C0311334|SEIZURE DIS GENERALIZED ONSET
C0311334|SEIZURE DIS CONVULSIVE GENERALIZED
C0311334|SEIZURE DIS GENERALIZED CONVULSIVE
C0311334|GENERALIZED SEIZURE DIS CONVULSIVE
C0311334|GENERALIZED ONSET SEIZURE DIS
C0311334|Convulsive Epilepsies, Generalized
C0311334|Convulsive Epilepsy, Generalized
C0311334|Epilepsies, Generalized Convulsive
C0311334|Epilepsy, Generalized Convulsive
C0311334|Generalized Convulsive Epilepsies
C0311334|Generalized convulsive epilepsy (disorder)
C0311334|Generalized convulsive epilepsy NOS
C0311334|Generalised convulsive epilepsy
C0311334|Generalised convulsive epilepsy NOS
C0311334|Generalized convulsive epilepsy
C0311334|Generalized convulsive epilepsy NOS (disorder)
C0311334|generalized convulsive seizure (diagnosis)
C0311334|generalized convulsive seizure
C0311334|epilepsy generalized convulsive
C0311334|Convulsive Seizure Disorder, Generalized
C0311334|Seizure Disorder, Generalized Onset
C0311334|Seizure Disorder, Generalized, Convulsive
C0311334|Seizure Disorder, Convulsive, Generalized
C0311334|Generalized Seizure Disorder, Convulsive
C0311334|Generalized Onset Seizure Disorder
C0311334|Generalised-onset seizures
C0311334|Generalized-onset seizures (disorder)
C0311334|Generalized-onset seizures
C0311334|epilepsy; generalized, convulsive
C0311334|generalized; epileptic, convulsive
C0311334|Generalized convulsive epilepsy, NOS
C0311334|Generalized-onset seizures, NOS
C0311334|Generalized convulsive epilepsy [dup] (disorder)
C0311334|Convulsive Generalized Seizure Disorder
C0149958|Complex partial seizures
C0149958|seizure partial (focal) complex
C0149958|complex partial seizure
C0149958|complex partial seizure (physical finding)
C0149958|partial complex seizure (diagnosis)
C0149958|partial complex seizure
C0149958|Partial complex seizures
C0149958|Seizures, complex partial
C0149958|Partial complex seizure (disorder)
C0149958|Partial seizures, complex
C0149958|Psychomotor fit
C0234972|Convulsive disorder
C0234972|convulsive disorder (diagnosis)
C0234972|Convulsion disorder
C0234972|Disorder convulsive
C0234972|Convulsive disorder NOS
C0238111|Lennox-Gastaut syndrome
C0238111|Lennox-Gastat syndrome
C0238111|Lennox Gastaut syndrome
C0238111|Gastaut syndrome
C0238111|Lennox-Gastant syndrome
C0238111|Lennox-Gastant syndrome (diagnosis)
C0238111|Lennox-Gastaut syndrome (disorder)
C0238111|Syndrome, Lennox Gastaut
C0238111|Gastaut Syndrome, Lennox
C0238111|Lennox Gastaut Syndromes
C0238111|Gastaut Syndromes, Lennox
C0238111|Syndromes, Lennox Gastaut
C0238111|Lennox Gastaut Syndrome [Disease/Finding]
C0238111|LGS
C0238111|Lennox-Gastaut
C0238111|Lennox-Gastaut syndrome (disorder) [Ambiguous]
C2236802|nonepileptic seizures (diagnosis)
C2236802|nonepileptic seizures
C2080645|photosensitive seizures (diagnosis)
C2080645|photosensitive seizures
C2349436|Migraine triggered seizures
C2349436|migraine triggered seizures (diagnosis)
C2349436|Migraine-Triggered Seizure
C0234974|Epilepsy, partial NOS, without impairment of consciousness
C0234974|Epilepsy, partial, without impairment of consciousness
C0234974|Simple partial seizures
C0234974|Simple partial seizures with consciousness preserved
C0234974|seizure partial (focal) simple
C0234974|simple partial seizure
C0234974|simple partial seizure (physical finding)
C0234974|partial simple seizure (diagnosis)
C0234974|partial simple seizure without impairment of consciousness (diagnosis)
C0234974|partial simple seizure
C0234974|partial simple seizure without impairment of consciousness
C0234974|Partial Seizures, Simple
C0234974|Seizures, Simple Partial
C0234974|Seizure;focal;simple partial
C0234974|Partial epilepsy without mention of impairment of consciousness
C0234974|Partial epilepsy without mention of impairment of consciousness (disorder)
C0234974|Simple partial seizure (disorder)
C0234974|Partial epilepsy without mention of impairment of consciousness NOS (disorder)
C0234974|Partial epilepsy without mention of impairment of consciousness NOS
C0234974|Focal seizures without impairment of consciousness or awareness
C0234974|Partial Seizures, Simple, Consciousness Preserved
C0234974|Simple partial seizure, consciousness not impaired
C0234974|Simple partial seizure, consciousness not impaired (disorder)
C0234974|seizure; epileptic, simple, partial
C0234974|simple partial seizures; epileptic
C0234974|Simple partial seizure, consciousness not impaired (finding)
C0234974|simple partial focal seizure
C0234974|Partial epilepsy, without mention of impairment of consciousness
C0270823|Status, Petit Mal
C0270823|Petit mal status
C0270823|Petit mal status epilepticus
C0270823|petit mal epilepsy status
C0270823|petit mal epilepsy status (diagnosis)
C0270823|Status, Absence
C0270823|Status epilepticus;Petit mal
C0270823|Petit mal status, epileptic
C0270823|Status epilepticus petit mal
C0270823|Absence Status
C0270823|Epileptic absence status
C0270823|Epilepsia minoris continua
C0270823|Petit-mal status
C0270823|Prolonged epileptic twilight state
C0270823|Status pyknolepticus
C0270823|Non-convulsive status epilepticus with impaired consciousness
C0270823|Spike wave stupor
C0270823|Petit mal status (disorder)
C0270823|confusional; state, epileptic
C0270823|epilepsy; status, absence
C0270823|epilepsy; status, petit mal
C0270823|epilepticus; status, petit mal
C0270823|absence; status
C0270823|petit mal; status
C0270823|state; confusional, epileptic
C0270823|status; absences
C0270823|status; absence
C0270823|status; epileptic, absence
C0270823|status; epileptic, petit mal
C0270823|status; epilepticus, petit mal
C0270823|status; petit mal
C0270823|twilight state; epileptic
C0270823|Epileptic confusional state
C0270823|Epileptic twilight state
C0311335|Grand mal status epilepticus
C0311335|grand mal epilepsy status
C0311335|grand mal epilepsy status (diagnosis)
C0311335|Grand mal status
C0311335|Status epilepticus;Grand mal
C0311335|Grand mal status, epileptic
C0311335|Convulsive status epilepticus
C0311335|Status epilepticus grand mal
C0311335|Status Epilepticus, Grand Mal
C0311335|Generalized Convulsive Status Epilepticus
C0311335|Status Epilepticus, Generalized Convulsive
C0311335|Grand mal status (disorder)
C0311335|epilepsy; status, grand mal
C0311335|epilepticus; status, grand mal
C0311335|grand mal; status
C0311335|status; epileptic, grand mal
C0311335|status; epilepticus, grand mal
C0311335|status; grand mal
C0751777|progressive familial myoclonic epilepsy
C0751777|progressive familial myoclonic epilepsy (diagnosis)
C0751777|Familial Progressive Myoclonic Epilepsy
C0751777|myoclonic; epileptic, progressive (familial)
C0751783|Disease, Lafora
C0751783|Lafora Disease
C0751783|Lafora's disease
C0751783|LBD
C0751783|MYOCLONIC EPILEPSY OF LAFORA
C0751783|EPM2A
C0751783|LAFORA DIS
C0751783|LAFORA BODY DIS
C0751783|Lafora body disease (diagnosis)
C0751783|Lafora body disease
C0751783|Disease, Lafora Body
C0751783|Lafora Type Progressive Myoclonic Epilepsy
C0751783|Epilepsy, Progressive Myoclonic, Lafora
C0751783|Progressive Myoclonic Epilepsy, Lafora Type
C0751783|Lafora Disease [Disease/Finding]
C0751783|Progressive Myoclonic Epilepsy, Lafora
C0751783|Lafora Progressive Myoclonic Epilepsy
C0751783|Disorder, Lafora Body
C0751783|Lafora Myoclonic Epilepsy
C0751783|Lafora Body Disorder
C0751783|Epilepsy Progressive Myoclonic 2
C0751783|Lafora's myoclonic epilepsy
C0751783|Lafora Progressive Myoclonus Epilepsy
C0751783|Progressive Myoclonus Epilepsy, Lafora Type
C0751783|Progressive Myoclonic Epilepsy Type 2
C0751783|Epilepsy, Progressive Myoclonic 2A
C0751783|EPILEPSY, PROGRESSIVE MYOCLONIC, 2A
C0751783|MELF
C0751783|EPM2
C0751783|Lafora disease (disorder)
C0751783|Lafora
C0037769|Infantile spasms
C0037769|Infantile Spasm
C0037769|Spasms, Infantile
C0037769|Syndrome, West
C0037769|infantile spasms (diagnosis)
C0037769|Attack, Lightning
C0037769|Attacks, Lightning
C0037769|Lightning Attack
C0037769|West syndrome
C0037769|Spasms, Infantile [Disease/Finding]
C0037769|Lightning Attacks
C0037769|Seizure;infant spasms
C0037769|West's syndrome
C0037769|West syndrome (disorder)
C0037769|Infantile spasms NOS
C0037769|West syndrome (finding)
C0037769|Infantile spasms NOS (disorder)
C0037769|Infantile spasms - hypsarrythmia
C0037769|Infantile spasms - hypsarrhythmia
C0037769|Lightning spasms
C0037769|West
C0037769|infantile; spasm
C0037769|lightning; spasm
C0037769|spasm; infantile
C0037769|spasm; lightning
C0270819|Cursive epilepsy
C0270819|cursive seizure (diagnosis)
C0270819|cursive seizure
C0270819|Epilepsies, Cursive
C0270819|Epilepsy, Cursive
C0270819|Reflex Epilepsies, Cursive (Running)
C0270819|Cursive Reflex Epilepsies (Running)
C0270819|Cursive Reflex Epilepsy (Running)
C0270819|Epilepsy, Cursive Reflex (Running)
C0270819|Running epilepsy
C0270819|Cursive (running) epilepsy
C0270819|Cursive (running) epilepsy (disorder)
C0270819|Cursive seizure (disorder)
C0270819|Reflex Epilepsy, Cursive (Running)
C0270819|Epilepsy, running
C0270820|Gelastic epilepsy
C0270820|gelastic seizure
C0270820|gelastic seizure (diagnosis)
C0270820|Epilepsies, Gelastic
C0270820|Gelastic Epilepsies
C0270820|Gelastic seizures
C0270820|Gelastic seizure (disorder)
C0270820|Epilepsy, gelastic
C0085543|Epilepsia Partialis Continua
C0085543|Syndrome, Kojewnikow's
C0085543|Syndrome, Kozhevnikov's
C0085543|Epilepsy, Kojevnikov's
C0085543|epilepsia partialis continua (diagnosis)
C0085543|Kojevnikov Epilepsy
C0085543|Epilepsy, Kojewnikov's
C0085543|Kojewnikov Epilepsy
C0085543|Syndrome, Kojewnikow
C0085543|Syndrome, Kozhevnikov
C0085543|Kojevnikov's Epilepsy
C0085543|Kojewnikow Syndrome
C0085543|Kojewnikow's Syndrome
C0085543|Kozhevnikov's Syndrome
C0085543|Kojewnikov's Epilepsy
C0085543|Epilepsia Partialis Continua [Disease/Finding]
C0085543|Kozhevnikov Syndrome
C0085543|Kojevnikov's Epilepsies
C0085543|Epilepsies, Kojevnikov's
C0085543|Kojevnikov's epilepsy (disorder)
C0085543|Focal status epilepticus
C0085543|Motor simple partial status
C0085543|Epilepsia partialis continua (disorder)
C0796133|RAMON SYNDROME
C0796133|Gingival fibromatosis combined with cherubism
C0796133|CHERUBISM, GINGIVAL FIBROMATOSIS, EPILEPSY, MENTAL DEFICIENCY, HYPERTRICHOSIS, AND STUNTED GROWTH
C1856929|EPILEPSY-TELANGIECTASIA
C1856929|Epilepsy telangiectasia
C0270709|RUD SYNDROME
C0270709|RUDS
C0270709|Ichthyosis hypogonadism mental retardation epilepsy syndrome
C0270709|Ichthyosis mental retardation-epilepsy hypogonadism syndrome
C0270709|Rud's syndrome
C0270709|Neuroichthyosis hypogonadism syndrome
C0270709|Dwarfism ichthyosiform erythroderma mental deficiency syndrome
C0270709|Ichthyosis oligophrenia epilepsy syndrome
C0270709|Ichthyosis male hypogonadism syndrome
C0270709|Dwarfism-ichthyosiform erythroderma-mental deficiency syndrome
C0270709|Rud's syndrome (disorder)
C1849508|EPILEPSY, PYRIDOXINE-DEPENDENT
C1849508|PDE
C1849508|EPD
C1849508|Pyridoxine dependency with seizures
C1849508|Pyridoxine-dependent epilepsy
C1849508|Pyridoxine dependency
C1849508|Aasa Dehydrogenase Deficiency
C1849508|Pyridoxine-Dependent Seizures
C1849508|Vitamin B6-Dependent Seizures
C0795900|Dwarfism, lean spastic type
C0795900|Coffin syndrome 1
C0795900|Lean spastic dwarfism
C0265339|BFLS
C0265339|BORJ
C0265339|BORJESON-FORSSMAN-LEHMANN SYNDROME
C0265339|Borjeson Syndrome
C0265339|Mental deficiency, epilepsy and endocrine disorders
C0265339|MRXSBFL
C0265339|Mental Deficiency, Epilepsy, And Endocrine Disorders
C0265339|Borjeson-Forssman-Lehmann syndrome (diagnosis)
C0265339|MENTAL RETARDATION, EPILEPSY, AND ENDOCRINE DISORDERS
C0265339|MENTAL RETARDATION, X-LINKED, SYNDROMIC, BORJESON-FORSSMAN-LEHMANN TYPE
C0265339|Borjeson-Forssman-Lehmann syndrome (disorder)
C0796202|Wittwer syndrome
C0265328|ALOPECIA-EPILEPSY-OLIGOPHRENIA SYNDROME OF MOYNAHAN
C0265328|Moynahan's syndrome (diagnosis)
C0265328|Moynahan's syndrome
C0265328|Moynahan syndrome
C0265328|Alopecia epilepsy oligophrenia syndrome of Moynahan
C0265328|Moynahan alopecia syndrome
C0265328|Progressive cardiomyopathic lentiginosis
C0265328|Moynahan's syndrome (disorder)
C1863090|ALOPECIA, PSYCHOMOTOR EPILEPSY, PYORRHEA, AND MENTAL SUBNORMALITY
C1863090|Congenital universal alopecia, epilepsy, mental subnormality and pyorrhea
C1863090|Alopecia, epilepsy, pyorrhea, mental subnormality
C1863090|Shokeir syndrome
C0406740|KOHLSCHUTTER-TONZ SYNDROME
C0406740|Epilepsy dementia amelogenesis imperfecta
C0406740|Epilepsy and yellow teeth
C0406740|Kohlschutter syndrome
C0406740|Kohlschutter Tonz syndrome
C0406740|Epilepsy, Dementia, And Amelogenesis Imperfecta
C0406740|KTZS
C0406740|Kohlschutter's syndrome
C0406740|disorders of central nervous system kohlschutter's syndrome
C0406740|Kohlschutter's syndrome (diagnosis)
C0406740|Amelocerebrohypohidrotic syndrome
C0406740|Epilepsy, dementia and amelogenesis imperfecta
C0406740|Epilepsy, mental deterioration and yellow teeth
C0406740|Kohlschutter's syndrome (disorder)
C2931451|Sandhaus Ben-Ami syndrome
C2931451|Patella hypoplasia skeletal malformations
C2931495|Arthrogryposis multiplex congenita with epileptic seizures and migrational brain disorder
C2931495|Arthrogryposis epileptic seizures migrational brain disorder
C1846278|MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, AND OBESITY
C1846278|MEHMO
C1846278|MENTAL RETARDATION, EPILEPTIC SEIZURES, HYPOGONADISM AND HYPOGENITALISM, MICROCEPHALY, AND OBESITY (disorder)
C1846278|MEHMO syndrome
C1846278|X-linked MEHMO syndrome
C1846278|MRXS20
C1846278|MRXS25
C1846278|MENTAL RETARDATION, X-LINKED, SYNDROMIC 25
C1846278|MENTAL RETARDATION, X-LINKED, SYNDROMIC 20
C0796046|GURRIERI SYNDROME
C0796046|Skeletal dysplasia epilepsy short stature
C0796046|Gurrieri Sammito Bellussi syndrome
C2931579|Battaglia Neri syndrome
C0796010|KIFAFA SEIZURE DISORDER
C0796010|Complex familial seizure disorder
C0796010|Vitsala
C2931668|Boudhina Yedes Khiari syndrome
C1838491|Pachygyria, mental retardation and epilepsy
C1838491|Pachygyria with mental retardation and seizures
C1838491|Kuzniecky syndrome
C1838491|PACHYGYRIA WITH MENTAL RETARDATION, SEIZURES, AND ARACHNOID CYSTS
C3472688|Single epileptic seizure (finding)
C3472688|Single epileptic seizure
C0751111|Epilepsy, Awakening
C0751111|Awakening Epilepsy
C0751110|Seizure, Single
C0751110|Seizures, Single
C0751110|Single Seizures
C0751110|Single seizure
C0751110|Single seizure (finding)
C0086237|Cryptogenic Epilepsies
C0086237|Cryptogenic Epilepsy
C0086237|Epilepsies, Cryptogenic
C0086237|Epilepsy, Cryptogenic
C0586323|ALCOHOL WITHDRAWAL IND SEIZURE
C0586323|Alcohol Withdrawal Induced Seizure
C0586323|Alcohol Withdrawal-Induced Seizures
C0586323|Seizure, Alcohol Withdrawal-Induced
C0586323|Seizures, Alcohol Withdrawal-Induced
C0586323|Withdrawal-Induced Seizure, Alcohol
C0586323|Withdrawal-Induced Seizures, Alcohol
C0586323|Alcohol Withdrawal Seizure
C0586323|Alcohol Withdrawal Seizures
C0586323|Seizure, Alcohol Withdrawal
C0586323|Seizures, Alcohol Withdrawal
C0586323|Withdrawal Seizure, Alcohol
C0586323|Withdrawal Seizures, Alcohol
C0586323|Alcoholic Seizure
C0586323|Alcoholic Seizures
C0586323|Seizure, Alcoholic
C0586323|Seizures, Alcoholic
C0586323|Alcohol Withdrawal-Induced Seizure
C0586323|Alcohol Withdrawal Seizures [Disease/Finding]
C0586323|Alcohol-induced epilepsy
C0586323|Alcohol-induced epilepsy (disorder)
C0586323|Rum fits
C0586323|Alcohol withdrawal-induced convulsion
C0586323|Alcohol-related fit
C0586323|Alcohol withdrawal-induced convulsion (disorder)
C0586323|Alcohol-related fit (finding)
C0586323|epilepsy; alcohol
C0586323|Alcohol-induced epilepsy [Ambiguous]
C0553754|Fit (in known epileptic) NOS
C0553754|Fit (in known epileptic) NOS (disorder)
C0553754|Fit (in known epileptic)
C1827389|Epilepsy, not refractory (disorder)
C1827389|Epilepsy, not refractory
C1827389|Epilepsy, not intractable
C1827389|epilepsy not intractable
C1827389|Epilepsy, not intractable (diagnosis)
C3649195|epilepsy, not intractable, with status epilepticus
C3649195|epilepsy not intractable with status epilepticus
C3649195|epilepsy, not intractable, with status epilepticus (diagnosis)
C3646244|seizures related to external causes (diagnosis)
C3646244|seizures related to external causes
C0472349|Localization-related symptomatic epilepsy
C0472349|epilepsy localization-related symptomatic
C0472349|Localization-related symptomatic epilepsy (diagnosis)
C0472349|Localisation-related symptomatic epilepsy
C0472349|Localization-related symptomatic epilepsy (disorder)
C0472349|epilepsy; localization-related, symptomatic
C0472348|epilepsy localization-related idiopathic (diagnosis)
C0472348|epilepsy localization-related idiopathic
C0472348|Localisation-related idiopathic epilepsy
C0472348|Localization-related idiopathic epilepsy
C0472348|Localization-related idiopathic epilepsy (disorder)
C0472348|epilepsy; idiopathic, localization-related
C0472348|epilepsy; localization-related, idiopathic
C3662042|Seizure disorder as sequela of stroke
C3662042|Seizure disorder as sequela of stroke (disorder)
C0751124|Atypical absence epilepsy
C0751124|Atypical absence epilepsy (disorder)
C0751124|Epilepsy, Absence, Atypical
C0086236|Atonic Epilepsies
C0086236|Atonic Epilepsy
C0086236|Epilepsies, Atonic
C0086236|Atonic epilepsy (disorder)
C0086236|Epilepsy, Atonic
C0086236|Epileptic seizures - atonic
C0086236|Epileptic seizures - atonic (finding)
C0393730|Self-induced non-photosensitive epilepsy
C0393730|Self-induced non-photosensitive epilepsy (diagnosis)
C0393730|epilepsy self-induced non-photosensitive
C0393730|Factitious epilepsy
C0393730|Self-induced non-photosensitive epilepsy (disorder)
C0393715|Drug-induced epilepsy (diagnosis)
C0393715|epilepsy drug-induced
C0393715|Drug-induced epilepsy
C0393715|Drug-induced epilepsy (disorder)
C3697594|Post-cerebrovascular accident epilepsy (disorder)
C3697594|Post-cerebrovascular accident epilepsy
C1837530|AICAR TRANSFORMYLASE/IMP CYCLOHYDROLASE DEFICIENCY
C1837530|AICA Ribosuria due to ATIC Deficiency
C1837530|AICAR Transformylase Inosine Monophosphate Cyclohydrolase Deficiency
C1837530|ATIC DEFICIENCY
C1837530|AICA-RIBOSURIA DUE TO ATIC DEFICIENCY
C1845343|EPILEPSY, X-LINKED, WITH VARIABLE LEARNING DISABILITIES AND BEHAVIOR DISORDERS
C1849416|RETINAL DEGENERATION AND EPILEPSY
C1845102|EPILEPTIC ENCEPHALOPATHY, EARLY INFANTILE, 8
C1845102|EIEE8
C1845102|Hyperekplexia and Epilepsy
C2751195|EPILEPSY, BENIGN NEONATAL, 1, AND/OR MYOKYMIA
C2751195|Epilepsy, Benign Neonatal, 1, And-Or Myokymia
C1845543|MRXSH
C1845543|MRXE
C1845543|MENTAL RETARDATION, X-LINKED, SYNDROMIC, HEDERA TYPE
C1845543|Mental Retardation, X-Linked, with Epilepsy
C1836824|AMISH INFANTILE EPILEPSY SYNDROME
C1836824|GM3 Synthase Deficiency
C1836824|Epilepsy Syndrome, Infantile-Onset Symptomatic
C1836824|SALT AND PEPPER MENTAL RETARDATION SYNDROME
C1843852|SPINOCEREBELLAR ATAXIA WITH EPILEPSY
C1843852|SCAE
C1843852|Myoclonic epilepsy myopathy sensory ataxia
C1843852|Myoclonic epilepsy myopathy sensory ataxia (disorder)
C1843852|MEMSA - myoclonic epilepsy myopathy sensory ataxia
C1970203|PMSE
C1970203|POLYHYDRAMNIOS, MEGALENCEPHALY, AND SYMPTOMATIC EPILEPSY
C1970203|PMSE SYNDROME
C1832437|MENTAL RETARDATION, MICROCEPHALY, EPILEPSY, AND COARSE FACE
C1853564|DEND
C1853564|DEVELOPMENTAL DELAY, EPILEPSY, AND NEONATAL DIABETES
C1853623|FRYNS-AFTIMOS SYNDROME
C1853623|Cerebrooculofacial Lymphatic Syndrome
C1853623|Pachygyria, Mental Retardation, Epilepsy, and Characteristic Facies
C1853623|Mental Retardation with Epilepsy and Characteristic Facies
C1853623|COFL SYNDROME
C2678194|MENTAL RETARDATION, X-LINKED, SYNDROMIC, CHRISTIANSON TYPE
C2678194|MRXSCH
C2678194|Mental Retardation, Microcephaly, Epilepsy, and Ataxia Syndrome
C2678194|Angelman-Like Syndrome, X-Linked
C2678194|christianson syndrome (diagnosis)
C2678194|christianson syndrome
C2678194|Intellectual Deficit, X-Linked, South African Type
C2678194|X-linked mental retardation syndrome, Christianson type (disorder)
C2678194|X-linked intellectual deficit, South African type
C2678194|X-linked mental retardation syndrome, Christianson type
C3837709|epilepsy, not intractable, without status epilepticus
C3837709|epilepsy not intractable without status epilepticus
C3837709|epilepsy, not intractable, without status epilepticus (diagnosis)
C3826393|Epilepsy in pregnancy
C3826393|Epilepsy in mother complicating pregnancy (disorder)
C3826393|Epilepsy in mother complicating pregnancy
C3840267|Epilepsy in childbirth
C3840267|Epilepsy in mother complicating childbirth
C3840267|Epilepsy in mother complicating childbirth (disorder)
C0751122|SMEI
C0751122|Infantile Severe Myoclonic Epilepsy
C0751122|EIEE6
C0751122|Syndromes, Dravet
C0751122|Dravet Syndromes
C0751122|Syndrome, Dravet
C0751122|Dravet syndrome
C0751122|Severe myoclonic epilepsy of infancy
C0751122|EPILEPTIC ENCEPHALOPATHY, EARLY INFANTILE, 6
C0751122|Severe Infantile Myoclonic Epilepsy
C0751122|Severe Myoclonic Epilepsy, Infantile
C0751122|Epilepsy, Myoclonic, Infantile, Severe
C0751122|Myoclonic Epilepsy, Infantile, Severe
C0751122|Myoclonic Epilepsy, Severe, Of Infancy
C0751122|Myoclonic Epilepsy, Severe Infantile
C0751122|Severe myoclonic epilepsy in infancy
C0751122|Severe myoclonic epilepsy in infancy (disorder)
C2363129|BECTS
C2363129|CENTRALOPATHIC EPILEPSY
C2363129|ECT
C2363129|Benign Rolandic Epilepsy
C2363129|Epilepsies, Centrotemporal
C2363129|Epilepsy, Centralopathic
C2363129|Rolandic Epilepsy, Benign
C2363129|Epilepsy, Benign Rolandic
C2363129|Epilepsies, Centralopathic
C2363129|Centrotemporal Epilepsies
C2363129|Centralopathic Epilepsies
C2363129|Benign Childhood Epilepsy With Centro Temporal Spikes
C2363129|Benign childhood epilepsy with centrotemporal spike (disorder)
C2363129|Benign childhood epilepsy with centrotemporal spike
C2363129|BENIGN EPILEPSY OF CHILDHOOD WITH CENTROTEMPORAL SPIKES
C2363129|Benign Childhood Epilepsy With Centrotemporal Spikes
C2363129|BRE
C2363129|TEMPORAL-CENTRAL FOCAL EPILEPSY
C2363129|CENTROTEMPORAL EPILEPSY
C2363129|BCECTS
C2363129|Benign Rolandic Epilepsy of Childhood
C2363129|Epilepsy, Centrotemporal
C2363129|Benign Childhood Epilepsy With Centro-Temporal Spikes
C2363129|Benign Epilepsy With Centrotemporal Spikes
C2363129|Benign Rolandic epilepsy (disorder)
C3889476|Benign Familial Neonatal Seizures
C3889476|Benign Familial Convulsions
C3889476|Benign Familal Neonatal Seizures
C3889476|Benign Familial Convulsion
C1846385|FOCAL CORTICAL DYSPLASIA OF TAYLOR
C1846385|FCDT
C1846385|CDT
C1846385|Cortical dysplasia of Taylor
C1846385|Focal cortical dysplasia, type 2
C1846385|Focal Cortical Dysplasia, Type II
C4064621|migraine triggered seizures without intractable migraine w/o status migrainosus
C4064621|migraine triggered seizures without intractable migraine without status migrainosus
C4064621|migraine triggered seizures without intractable migraine without status migrainosus (diagnosis)
C4064624|migraine triggered seizures with intractable migraine without status migrainosus
C4064624|migraine triggered seizures with intractable migraine without status migrainosus (diagnosis)
C4064623|migraine triggered seizures without intractable migraine (diagnosis)
C4064623|migraine triggered seizures without intractable migraine
C4064622|migraine triggered seizures without intractable migraine with status migrainosus (diagnosis)
C4064622|migraine triggered seizures without intractable migraine with status migrainosus
C0270825|Visceral epilepsy
C0270825|Visceral epilepsy (disorder)
C0270825|epilepsy; visceral
C0270825|visceral; epileptic
C0270825|Epilepsy, visceral
C0270824|visual partial simple seizure (diagnosis)
C0270824|visual partial simple seizure
C0270824|Seizure, Visual
C0270824|Visual Seizure
C0270824|Visual Seizures
C0270824|Seizures, Visual
C0270824|Visual epilepsy
C0270824|Visual epilepsy (disorder)
C0270824|epilepsy; visual
C0270824|visual; epileptic
C0270824|Epilepsy, visual
C0347873|Psychosensory epilepsy
C0347873|Psychosensory epilepsy (disorder)
C0347873|epilepsy; psychosensory
C0347873|psychosensory; epileptic
C0347873|Epilepsy, psychosensory
C0347874|Somatosensory epilepsy
C0347874|Somatosensory epilepsy (disorder)
C0347874|epilepsy; somatosensory
C0347874|somatosensory; epileptic
C0347874|Epilepsy, somatosensory
C0014549|Epilepsies, Tonic-Clonic
C0014549|Epilepsy, Tonic Clonic
C0014549|Epilepsy, Tonic-Clonic
C0014549|Grand Mal Epilepsy
C0014549|Tonic-Clonic Epilepsies
C0014549|Tonic-Clonic Epilepsy
C0014549|TONIC CLONIC CONVULSION DIS
C0014549|MAJOR MOTOR SEIZURE DIS
C0014549|SEIZURE DIS TONIC CLONIC
C0014549|TONIC CLONIC SEIZURE DIS
C0014549|GRAND MAL SEIZURE DIS
C0014549|SEIZURE DIS GRAND MAL
C0014549|SEIZURE DIS MAJOR MOTOR
C0014549|generalized convulsive tonic-clonic seizure
C0014549|generalized convulsive grand mal seizure
C0014549|tonic-clonic epilepsy (diagnosis)
C0014549|Convulsion Disorder, Tonic-Clonic
C0014549|Convulsion Disorders, Tonic-Clonic
C0014549|Disorder, Tonic-Clonic Convulsion
C0014549|Disorders, Tonic-Clonic Convulsion
C0014549|Tonic Clonic Convulsion Disorder
C0014549|Tonic-Clonic Convulsion Disorders
C0014549|Convulsion Syndrome, Tonic-Clonic
C0014549|Convulsion Syndromes, Tonic-Clonic
C0014549|Syndrome, Tonic-Clonic Convulsion
C0014549|Syndromes, Tonic-Clonic Convulsion
C0014549|Tonic Clonic Convulsion Syndrome
C0014549|Tonic-Clonic Convulsion Syndromes
C0014549|Convulsion, Tonic Clonic
C0014549|Convulsions, Tonic Clonic
C0014549|Tonic Clonic Convulsion
C0014549|Disorder, Tonic-Clonic Seizure
C0014549|Disorders, Tonic-Clonic Seizure
C0014549|Seizure Disorder, Tonic-Clonic
C0014549|Seizure Disorders, Tonic-Clonic
C0014549|Tonic Clonic Seizure Disorder
C0014549|Tonic-Clonic Seizure Disorders
C0014549|Seizure Syndrome, Tonic-Clonic
C0014549|Seizure Syndromes, Tonic-Clonic
C0014549|Syndrome, Tonic-Clonic Seizure
C0014549|Syndromes, Tonic-Clonic Seizure
C0014549|Tonic Clonic Seizure Syndrome
C0014549|Tonic-Clonic Seizure Syndromes
C0014549|Convulsion, Grand Mal
C0014549|Grand Mal Convulsion
C0014549|Grand Mal Convulsions
C0014549|Major Epilepsies
C0014549|Major Epilepsy
C0014549|Major Motor Seizure Disorder
C0014549|Tonic-Clonic Convulsion Syndrome
C0014549|Epilepsy, Tonic-Clonic [Disease/Finding]
C0014549|Tonic Clonic Convulsions
C0014549|Epilepsy, Major
C0014549|Tonic-Clonic Convulsion Disorder
C0014549|Seizure Disorder, Grand Mal
C0014549|Tonic-Clonic Seizure Syndrome
C0014549|Epilepsy, Grand Mal
C0014549|Grand Mal Seizure Disorder
C0014549|Seizure Disorder, Major Motor
C0014549|Convulsions, Grand Mal
C0014549|Seizure Disorder, Tonic Clonic
C0014549|Tonic-Clonic Seizure Disorder
C0014549|Epilepsy;grand mal
C0014549|Tonic-clonic convulsion
C0014549|Clonic-tonic convulsions
C0014549|Grand mal
C0014549|Convulsion grand mal
C0014549|Major convulsion
C0014549|Convulsions grand mal
C0014549|Epilepsy grand mal
C0014549|Tonic/ clonic convulsions
C0014549|grand mal seizure
C0014549|grand mal seizure (diagnosis)
C0014549|Tonic-clonic epilepsy (disorder)
C0014549|epilepsy; grand mal
C0014549|epilepsy; major
C0014549|grand mal; epilepsy
C0014549|major; epileptic
C0014549|Epileptic seizures, tonic-clonic
C0472355|Epilepsy undetermined whether focal or generalised
C0472355|Epilepsy undetermined whether focal or generalized
C0472355|Epilepsy undetermined whether focal or generalized (disorder)
C0438419|Unilateral epilepsy (situation)
C0438419|Unilateral epilepsy (disorder)
C0438419|Unilateral epilepsy
C0477372|Other status epilepticus
C0477372|[X]Other status epilepticus
C0477372|[X]Other status epilepticus (disorder)
C0270822|Centerncephalic epilepsy
C0270822|Centrencephalic epilepsy (disorder)
C0270822|Centrencephalic epilepsy
C0270822|Centrencephalic absence
C0270822|Centerncephalic absence
C0347869|akinetic epilepsy
C0347869|Akinetic Epilepsies
C0347869|Epilepsies, Akinetic
C0347869|Akinetic seizures
C0347869|Epilepsy, Akinetic
C0347869|Epileptic seizures - akinetic
C0347869|Epileptic seizures - akinetic (finding)
C0347869|epilepsy; akinetic
C0347869|akinetic; epileptic
C0347869|akinetic; seizures
C0347869|seizure; akinetic
C0347869|Seizures, akinetic
C0347870|Epileptic seizures - clonic
C0347870|Epileptic seizures - clonic (finding)
C0347870|Epileptic seizures, clonic
C0086241|Epilepsies, Tonic
C0086241|Tonic Epilepsies
C0086241|Tonic Epilepsy
C0086241|Epileptic seizures - tonic
C0086241|Epileptic seizures - tonic (finding)
C0086241|epilepsy; tonic
C0086241|tonic; epileptic
C0086241|Epilepsy, Tonic
C0086241|Epileptic seizures, tonic
C0422855|Seizure, Vertiginous
C0422855|Vertiginous Seizure
C0422855|Vertiginous Seizures
C0422855|Seizure, Vestibular
C0422855|Vestibular Seizure
C0422855|Vestibular Seizures
C0422855|Vertiginous seizure (disorder)
C0422855|Seizures, Vertiginous
C0422855|Seizures, Vestibular
C0422855|Epileptic vertigo
C0422855|Vertiginous epilepsy
C0422855|Epileptic vertigo (disorder)
C0422855|epileptic; vertigo
C0422855|vertigo; epileptic
C0422855|Vertiginous seizure (finding)
C0159020|Convulsions of newborn
C0159020|convulsions in newborn (diagnosis)
C0159020|convulsions in newborn
C0159020|Convulsion neonatal
C0159020|Convulsions in newborn (disorder)
C0159020|Neonatal Seizure
C0159020|Neonatal convulsion
C0159020|Neonatal fit
C0159020|Neonatal seizures
C0159020|Convulsions neonatal
C0159020|Convulsions in the newborn
C0159020|Fits in the newborn
C0159020|Seizures in the newborn
C0159020|Fits in newborn
C0159020|Neonatal convulsions
C0159020|Seizures in newborn
C0159020|Convulsions in the newborn (disorder)
C0159020|convulsions; neonatal
C0159020|convulsions; newborn
C0159020|fit; newborn
C0159020|neonatal; convulsions
C0159020|newborn; convulsions
C0159020|newborn; fit
C0270826|Unclassified epileptic seizures
C0270826|Unclassified epileptic seizures (disorder)
C0393707|Situation-related seizures
C0393707|Situation-related seizures (disorder)
C1299598|Seizures due to metabolic disorder (disorder)
C1299598|Seizures due to metabolic disorder
C0871737|Experimental Epilepsy
C0857345|Late onset epilepsy
C1328935|nocturnal focal lobe epilepsy
C0700438|Headache, Sick
C0700438|Headaches, Sick
C0700438|Sick Headaches
C0700438|"Sick" headaches
C0700438|Sick Headache
C0700438|Sick headache (disorder)
C0553587|Epilepsy, partial, with impairment of consciousness
C0553587|Partial epilepsy with impairment of consciousness NOS
C0553587|Partial epilepsy with impairment of consciousness NOS (disorder)
C0553587|Partial epilepsy, with impairment of consciousness
C0553587|Partial epilepsy with impairment of consciousness
C0553587|Partial epilepsy with impairment of consciousness (disorder)
C0544645|Focal Sensory Seizures
C0544645|Seizure, Focal Sensory
C0544645|Seizures, Focal Sensory
C0544645|Sensory Seizure, Focal
C0544645|Sensory Seizures, Focal
C0544645|Partial Sensory Seizures
C0544645|Seizure, Partial Sensory
C0544645|Seizures, Partial Sensory
C0544645|Sensory Seizure, Partial
C0544645|Sensory Seizures, Partial
C0544645|Partial Sensory Seizure
C0544645|Focal Sensory Seizure
C0270854|Epilepsy, Symptomatic Generalized
C0270854|Generalized Epilepsy, Symptomatic
C0270854|Symptomatic Generalized Epilepsy
C0270854|Symptomatic generalised epilepsy
C0270854|Symptomatic generalized epilepsy (disorder)
C0270854|Symptomatic generalized epilepsy, NOS
C0154721|Epilepsy, unspecified, without mention of intractable epilepsy
C0154721|Epilep NOS w/o intr epil
C0154722|Epilepsy, unspecified, with intractable epilepsy
C0154722|Epilepsy NOS w intr epil
C1395129|dementia; epilepsy (etiology)
C1395129|dementia; epilepsy (manifestation)
C1395129|epilepsy; dementia (etiology)
C1395129|epilepsy; dementia (manifestation)
C1387228|postictal in epilepsy; amnesia
C1387228|amnesia; postictal in epilepsy
C1392243|cerebral; dysrhythmia
C1394140|cortical; dysrhythmia
C1395970|dysrhythmia; cerebral or cortical
C0391957|epilepsy; idiopathic
C0391957|idiopathic; epileptic
C1397835|fugue; postictal in epilepsy
C1397835|postictal in epilepsy; fugue
C0751778|Epilepsies, Progressive Myoclonic
C0751778|Myoclonic Epilepsies, Progressive
C0751778|Progressive Myoclonic Epilepsies
C0751778|Epilepsy, Progressive Myoclonic
C0751778|Myoclonic epilepsy, progressive
C0751778|Epilepsies, Progressive Myoclonus
C0751778|Epilepsy, Progressive Myoclonus
C0751778|Myoclonus Epilepsies, Progressive
C0751778|Progressive Myoclonus Epilepsy
C0751778|Progressive myoclonic epilepsy
C0751778|Myoclonic Epilepsies, Progressive [Disease/Finding]
C0751778|Progressive Myoclonus Epilepsies
C0751778|Progressive myoclonic epilepsy (disorder)
C0751778|Progressive myoclonic epilepsy (disorder) [Ambiguous]
C0852977|Epilepsy aggravated
C0852977|Aggravated Epilepsy
C0854109|Epilepsy congenital
C0854109|Congenital Epilepsy
C0270849|Extratemporal epilepsy
C0270849|Extratemporal epilepsy (disorder)
C1332300|Anosognostic Epilepsy
C1857575|CONVULSIVE DISORDER, FAMILIAL, WITH PRENATAL OR EARLY ONSET
