T131|SNOMEDCT_US|Hazardous or Poisonous Substance|allergy
T046|SNOMEDCT_US|Pathologic Function|allergy
T195|RXNORM|Antibiotic|allergy,medication

T061|SNOMEDCT_US|Therapeutic or Preventive Procedure|immunization,procedure,treatment

T109|RXNORM|Organic Chemical|medication,allergy,lab,?
T121|RXNORM|Pharmacologic Substance|medication,lab,diagnosis?,?
T196|RXNORM|Element, Ion, or Isotope|medication,lab,physical_exam

T123|LNC|Biologically Active Substance|medication,lab,?

T184|SNOMEDCT_US|Sign or Symptom|problem
T047|SNOMEDCT_US|Disease or Syndrome|diagnosis,problem
T037|SNOMEDCT_US|Injury or Poisoning|diagnosis,problem,allergy
T190|SNOMEDCT_US|Anatomical Abnormality|diagnosis,problem

T127|SNOMEDCT_US|Vitamin|lab,?

T025|LNC|Cell|lab
T126|LNC|Enzyme|lab
T116|LNC|Amino Acid, Peptide, or Protein|lab
T034|LNC|Laboratory or Test Result|lab,physical_exam
T059|LNC|Laboratory Procedure|lab,physical_exam,procedure
T060|LNC|Diagnostic Procedure|lab,physical_exam,procedure

T023|SNOMEDCT_US|Body Part, Organ, or Organ Component|physical_exam
T029|SNOMEDCT_US|Body Location or Region|physical_exam
T040|SNOMEDCT_US|Organism Function|physical_exam
