C0009170|Cocaine
C0085163|Crack Cocaine
C0002763|Central Nervous System Stimulants
C2203924|methylphenidate abuse
C1456332|Stimulant abuse
C3509122|stimulant abuse with stimulant-induced disorder
C2874625|Other stimulant abuse
C2874626|Other stimulant abuse, uncomplicated
C2874631|Other stimulant abuse with intoxication, unspecified
C3494717|Catha edulis abuse
C3509117|stimulant abuse - uncomplicated
C3509118|stimulant abuse with intoxication
C3509119|stimulant abuse with intoxication - uncomplicated
C3509120|stimulant abuse with intoxication delirium
C3662831|Nondependent amphetamine abuse
C4481000|other stimulant abuse in remission
C2874632|Other stimulant abuse with stimulant-induced mood disorder
C2874636|Other stimulant abuse with stimulant-induced psychotic disorder, unspecified
C2874637|Other stimulant abuse with other stimulant-induced disorder
C2874638|Other stimulant abuse with stimulant-induced anxiety disorder
C2874639|Other stimulant abuse with stimulant-induced sexual dysfunction
C2874640|Other stimulant abuse with stimulant-induced sleep disorder
C2874641|Other stimulant abuse with unspecified stimulant-induced disorder
C3509123|stimulant abuse with stimulant-induced anxiety disorder
C3509124|stimulant abuse with stimulant-induced sexual function
C3509125|stimulant abuse with stimulant-induced sleep disorder
C3509126|stimulant abuse with stimulant-induced mood disorder
C3509127|stimulant abuse with stimulant-induced psychotic disorder
C3509128|stimulant abuse with stimulant-induced psychotic disorder with delusions
C3509129|stimulant abuse with stimulant-induced psychotic disorder with hallucinations
C0553808|Nondependent amphetamine or other psychostimulant abuse
C2874628|Other stimulant abuse with intoxication, uncomplicated
C2874629|Other stimulant abuse with intoxication delirium
C3509121|stimulant abuse with intoxication with perceptual disturbance
C3836657|nondependent intravenous amphetamine abuse
C2874634|Other stimulant abuse with stimulant-induced psychotic disorder with delusions
C2874635|Other stimulant abuse with stimulant-induced psychotic disorder with hallucinations
C0338682|Nondependent amphetamine or psychostimulant abuse, continuous
C0338683|Nondependent amphetamine or psychostimulant abuse, episodic
C0338684|Nondependent amphetamine or psychostimulant abuse in remission
C2874630|Other stimulant abuse with intoxication with perceptual disturbance
C0085163|Cocaine, Crack
C0085163|Crack Cocaine
C0085163|free base cocaine
C0085163|Crack Cocaine [Chemical/Ingredient]
C0085163|Crack
C0085163|Cocaine freebase
C0085163|Rocks - cocaine
C0085163|Cocaine freebase (substance)
C0009169|Coca
C0009169|Erythroxylum coca Lam.
C0009169|Cocas
C0009169|Erythroxylons
C0009169|Erythroxylon
C0009169|Coca plant
C0009169|Cocaine plant
C0009169|Erythroxylum coca
C0009169|Erythroxylum coca (organism)
C0009169|hayo
C0975799|COCAINE HCL PWDR
C0975799|Cocaine HCl Powder
C0975799|COCAINE HCL PWDR [VA Product]
C0009170|Cocaine
C0009170|8-Azabicyclo(3.2.1)octane-2-carboxylic acid, 3-(benzoyloxy)-8-methyl-, methyl ester, (1R-(exo,exo))-
C0009170|(1R,2R,3S,5S)-2-Methoxycarbonyltropan-3-yl Benzoate
C0009170|Cocaine [Chemical/Ingredient]
C0009170|cocaine (Schedule I substance)
C0009170|Blow
C0009170|C
C0009170|Snow
C0009170|Coke
C0009170|Coca
C0009170|Cocaine product
C0009170|Cocaine (product)
C0009170|Cocaine (substance)
C2315434|Nasal form cocaine (product)
C2315434|Nasal form cocaine
C2315442|Ophthalmic form cocaine (product)
C2315442|Ophthalmic form cocaine
C2316909|Oropharyngeal form cocaine (product)
C2316909|Oropharyngeal form cocaine
C2316959|Oral form cocaine
C2316959|Oral form cocaine (product)
C0282108|Cocaine Hydrochloride
C0282108|Hydrochloride, Cocaine
C0282108|cocaine hydrochloride (medication)
C0282108|Methyl 3-beta-hydroxy-1-alpha-H,5-alpha-H-tropan-2-beta-carboxylate, benzoate (ester) HCl
C0282108|Cocaine Hydrochloride [Chemical/Ingredient]
C0282108|Cocaine HCl
C0282108|HCl, Cocaine
C0282108|Cocaine hydrochloride (substance)
C0171681|RTI-82
C0171681|8-Azabicyclo(3.2.1)octane-2-carboxylic acid, 3-(4-chlorophenyl)-8-methyl-, 2-(4-azido-3-iodophenyl)ethyl ester, (exo,exo)-
C0171681|RTI 82
C0532637|trimethylstannyl-(2-carbomethoxy-3-(4-phenyl)tropane)
C0532637|trimethylstannyl-beta-CT
C3472752|C-Topical
C0991509|Flake
C0991509|Flake Dosage Form
C0991509|Flake Dose Form
C0991509|Flakes
C0991509|Flakes (product)
C0991509|Oral Flakes
C0991509|Oral Flakes [Dose Form]
C0350656|Morphine + cocaine elixir
C0350656|Morphine + cocaine elixir (product)
C0350656|Morphine + cocaine elixir (substance)
C0359982|Cocaine Hydrochloride Powder
C0359982|Cocaine hydrochloride powder BP
C0359982|Cocaine hydrochloride powder (product)
C0359982|Cocaine hydrochloride powder BP (product)
C0359982|Cocaine hydrochloride powder BP (substance)
C0359981|Cocaine powder BP (product)
C0359981|Cocaine powder BP
C0359981|Cocaine powder BP (substance)
C0350555|Cocaine [no drugs here] (product)
C0350555|Cocaine [no drugs here]
C0350555|Cocaine [no drugs here] (substance)
C1985612|Cocaine &#x7C; urine
C1985611|Cocaine &#x7C; unknown substance
C0082060|benzoylecgonine ethyl ester
C0082060|coca-ethylene
C0082060|cocaethylene
C0082060|ethylcocaine
C0082060|Cocaethylene (substance)
C0053258|benzoyl ecgonine
C0053258|benzoylecgonine
C0053258|Benzoylecgonine (substance)
C1985608|Cocaine &#x7C; meconium
C1985609|Cocaine &#x7C; saliva
C1985613|Cocaine &#x7C; vitreous fluid
C0058917|ecgonine methyl ester
C0058917|methyl ecgonine
C1985610|Cocaine &#x7C; stool
C1985607|Cocaine &#x7C; hair
C1985606|Cocaine &#x7C; gastric fluid
C1455816|Cocaine metabolites
C1455816|Cocaine metabolite
C1455816|Cocaine metabolite (substance)
C1985605|Cocaine &#x7C; bld-ser-plas
C1985604|Cocaine &#x7C; bile fluid
C0250237|3-hydroxybenzoylecgonine
C0250237|m-hydroxybenzoylecgonine
C1985614|Cocaine &#x7C; XXX
C1624743|Cocaine+Benzoylecgonine
C0212482|RTI-121
C0212482|8-Azabicyclo(3.2.1)octane-2-carboxylic acid, 3-(4-iodophenyl)-8-methyl-, 1-methylethyl ester, (1R-(exo,exo))-
C0212482|RTI 121
C0909999|3-2-FTCAME
C0909999|3-4-FTCAME
C0909999|3beta-(2(18F)-fluoromethylphenyl)tropane-2beta-carboxylic acid methyl ester
C0909999|3beta-(2-fluoromethylphenyl)tropane-2beta-carboxylic acid methyl ester
C0068973|8-Azabicyclo(3.2.1)oct-8-yloxy, 3-(benzoyloxy)-2-(methoxycarbonyl)-, (1R-(exo,exo))-
C0068973|norcocaine nitroxide
C1611404|6-methyl-3-(4-iodo)phenyltropane-2-carboxylic acid methyl ester
C1611404|6-methyl-IPTCAME
C0676235|3-((2'-hydroxy-4'-iodobenzoyl)oxy)-8-methyl-8-azabicyclo(3.2.1)octane-2-carboxylic acid isopropyl ester
C0676235|3-HIO-MAOCA iProp
C0656790|3-(4-iodophenyl)tropan-2beta-carboxylic acid phenyl ester
C0656790|8-Azabicyclo(3.2.1)octane-2-carboxylic acid, 3-(4-iodophenyl)-8-methyl-, phenyl ester, (1R-(exo,exo))-
C1256547|(1R-(exo,exo))-3-(4-fluorophenyl)-8-methyl-8- azabicyclo(3.2.1)octane-2-carboxylic acid, methyl ester
C2352975|2-carbomethoxy-3-(3'-iodophenyl)tropane
C0655454|norcocaethylene
C0254083|N-nor-3-(4'-iodophenyl)tropane-2-carboxylic acid methyl ester
C0254083|N-nor-CIT
C0254083|nor-beta-CIT
C0386427|noranhydroecgonine
C0909543|tropoxene
C0140997|RTI-COC 32
C0140997|RTI-COC-32
C0140997|RTI 32
C0140997|RTI-32
C0244553|4'-hydroxybenzoylecgonine methyl ester
C0244553|4'-hydroxycocaine
C0244553|p-hydroxycocaine
C0620835|3'-hydroxy-4'-methoxycocaine
C0650345|methyl 8-benzoyl-3-hydroxy-8-azabicyclo(3.2.1)octane-2-carboxylate
C0650345|N-benzoylnormethylecgonine
C1308577|2-propanoyl-3-(2-naphthyl)-tropane
C0131123|methyl 3-benzoyloxy-8-formyl-8-azabicyclo(3.2.1)octane-2-carboxylate
C0131123|N-formylnorcocaine
C0531553|2-carbomethoxy-3-(4-fluorophenyl)-N-(1-iodoprop-1-en-3-yl)nortropane
C0531553|N-iodoallyl-2-carbomethoxy-3-(4-fluorophenyl)tropane
C0531553|IACFT
C3492805|benzoylecgonine isopropyl ester
C3492416|3-(4-fluorobenzoyloxy)tropane
C3492416|fluorotropacocaine
C3492416|3-pseudotropyl 4-fluorobenzoate
C0649823|3-iodo-4-azidococaine
C0649823|IACoc
C0103379|anhydroecgonine methyl ester
C0103379|anhydromethylecgonine
C0103379|methylecgonidine
C0909656|4'-isopropylnortropane-2-beta-carboxylic acid methyl ester
C0620837|4'-hydroxy-3'-methoxybenzoylecgonine methyl ester
C0620837|4'-hydroxy-3'-methoxycocaine
C0909360|8-oxa-norcocaine
C0909360|8-oxanorcocaine
C1452804|N-(2-fluoroethyl)-3beta-(4-iodophenyl)-8-methyl-8-azabicyclo(3.2.1)octane-2alpha-carboxamide
C1452804|N-F-IMA-OC
C1872843|AIMAOC methyl ester
C1872843|3-(4'-azido-3'-iodobiphenyl-4-yl)-8-methyl-8-azabicyclo(3.2.1)octane-2-carboxylic acid methyl ester
C0620844|3'-hydroxybenzoylecgonine methyl ester
C0620844|3'-hydroxycocaine
C1699433|8-((E)-4-fluoro-but-2-enyl)-3beta-p-tolyl-8-aza-bicyclo(3.2.1)octane-2beta-carboxylic acid methyl ester
C0530288|4'-phenylcocaine
C0964123|4-hydroxybenzoylecgonine
C0964123|p-OHBZE
C3657183|6-(3-(benzoyloxy)-8-methyl-8-azabicyclo(3.2.1)octane-2-carboxoamido)hexanoic acid
C3657183|GNE compound
C0077387|2-methoxycarbonyl-3-phenyltropane
C0077387|troparil
C0140994|RTI 55
C0140994|RTI-55
C0055761|cinnamoylcocaine
C0256893|2-carbomethoxy-3-(bis(4-fluorophenyl)methoxy)tropane
C0256893|difluoropine
C0910000|3-FTCAME
C0910000|3beta-(4(18F)-fluoromethylphenyl)tropane-2beta-carboxylic acid methyl ester
C0910000|3beta-(4-fluoromethylphenyl)tropane-2beta-carboxylic acid methyl ester
C0909657|(4'-isopropenyl-phenyl)nortropane-2-beta-carboxylic acid methylester
C0758316|RTI-113
C0967017|8-methyl-3-(4-methylphenyl)tropane--2-carboxylic acid N-methyl-N-(4-nitrobenzo-2-oxa-1,3-diazol-7-yl)ethanolamine ester
C0249751|methyl 3-benzoyloxy-7-methoxy-8-methyl-8-azabicyclo(3.2.1)octane-2-carboxylate
C0249751|methyl BMAOC
C0254073|N-nor-3-(4'-ethylphenyl)tropane-2-carboxylic acid methyl ester
C0254073|NETCME
C0531551|2-carbomethoxy-3-(3,4-dichlorophenyl)tropane
C0531551|CDCT cpd
C0531551|dichloropane
C0058916|3 beta-hydroxy-2 beta-tropanecarboxylic acid
C0058916|ecgonine
C0058916|Ecgonine (product)
C0058916|Ecgonine (substance)
C0669003|3-(4-ethyl-3-iodophenyl)nortropane-2-carboxylic acid methyl ester
C0669003|EINCA methyl ester
C0659449|ethylecgonine
C0659449|ethyl ecgonine
C3713617|SNC-rCTB vaccine
C0252165|4'-fluorococaine
C0540637|RTI 352
C0540637|RTI-352
C1610300|7-methyl IPTCAME
C1610300|7-methyl-3-(4-iodo)phenyltropane-2-carboxylic acid methyl ester
C0094945|3-(4-chlorophenyl)tropane-2-carboxylic acid methyl ester
C2974274|methyl-8-((2-(fluoromethyl)cyclopropyl)methyl)-3-phenyl-8-azabicyclo(3.2.1)octane-2-carboxylate
C2974274|PR17.MZ
C0077383|benzoyltropeine
C0077383|exo-8-methyl-8-azabicyclo(3.2.1)octan-3-ol, benzoate (ester)
C0077383|tropacocaine
C1142737|anhydroecgonine methyl ester N-oxide
C0050097|8-hydroxynorcocaine
C0534033|RTI 130
C0534033|RTI-130
C0171107|cocaine methiodide
C0255561|2-PTT
C0255561|2-propanoyl-3-(4-toluyl)tropane
C0255561|2-propanoyl-3-(4-tolyl)tropane
C0081740|benzoylnorecgonine
C0081740|norbenzoylecgonine
C1452515|cocaine N-oxide
C1570541|3-(3-fluoro-4-methylphenyl)nortropane-2-carboxylic acid methyl ester
C1570541|3-FMNCA methyl ester
C1741593|4,5,6,7,8,9,10,11,13,17a,18,19,20,21,22,22a-hexadecahydro-23-methyl-14,17-etheno-19,22-imino-1H-cyclohept(c)(1,9)oxaazacyclononadecine-3,12-dione
C1741593|hexadecahydro-MEICOD
C0676233|4'-iodococaine
C0909655|3-beta-(4'-n-propyl)nortropane-2-beta-carboxylic acid methyl ester
C0631334|3-(benzyloxy)-2-carbomethoxy-2-tropene
C0631334|2,3-dehydrococaine
C0300695|2'-fluoroethyl 8-methyl-3-(4-chlorophenyl)-8-azabicyclo(3.2.1)octane-2-carboxylate
C0300695|FECT-4ClP
C0612504|N-allylnorcocaine
C0909646|RTI 117
C0909646|RTI-117
C0300693|2'-fluoroethyl 8-methyl-3-(4-methylphenyl)-8-azabicyclo(3.2.1)octane-2-carboxylate
C0300693|FETT-4MP
C0608545|exo-8-azabicyclo(3.2.1)octan-3-ol, benzoate (ester)
C0608545|nortropacocaine
C1740172|5,6,7,8,10,14a,15,16,17,18,19,19a-dodecahydro-20-methyl-11,14-etheno-16,19-iminocyclohept(c)(1,9)oxaazacyclohexadecine-3,9(1H,4H)-dione
C1740172|dodecahydro-MEIOD
C0068972|norcocaine
C3847743|Cocaine+Metabolites &#x7C; Saliva
C3849705|8-(2-fluoroethyl)-3-(4-iodophenyl)-8-azabicyclo(3.2.1)octane-2-carboxylic acid methyl ester
C3849705|FE-beta-CIT
C3883790|FE@IPCIT
C3883790|2-fluoroethyl 8-(3-iodoprop-2-en-1-yl)-3-(4-iodophenyl)-8-azabicyclo(3.2.1)octane-2-carboxylate
C0359988|Cocaine 100 MG/ML Nasal Solution
C0359988|cocaine 10 % Nasal Solution
C0359988|Cocaine 10% nasal drops
C0359988|Cocaine 10% nasal drops (product)
C0359988|Cocaine 10% nasal drops (substance)
C0359989|Cocaine 0.1 MG/MG Paste
C0359989|cocaine 10 % Paste
C0359989|Cocaine 10% paste
C0359989|Cocaine 10% paste (product)
C0359989|Cocaine 10% paste (substance)
C0359985|Cocaine 200 MG/ML Ophthalmic Solution
C0359985|cocaine 20 % Ophthalmic Solution
C0359985|Cocaine 20% eye drops
C0359985|Cocaine 20% eye drops (product)
C0359985|Cocaine 20% eye drops (substance)
C0357721|Cocaine 40 MG/ML Ophthalmic Solution
C0357721|cocaine 4 % Ophthalmic Solution
C0357721|Cocaine 4% preservative-free eye drops
C0357721|Cocaine hydrochloride 4% eye drops
C0357721|Cocaine 4% preservative-free eye drops (product)
C0357721|Cocaine hydrochloride 4% eye drops (product)
C0357721|Cocaine 4% preservative-free eye drops (substance)
C0357721|Cocaine hydrochloride 4% eye drops (substance)
C0359984|Cocaine 50 MG/ML Ophthalmic Solution
C0359984|cocaine 5 % Ophthalmic Solution
C0359984|Cocaine 5% eye drops
C0359984|Cocaine 5% eye drops (product)
C0359984|Cocaine 5% eye drops (substance)
C0359987|Cocaine hydrochloride 10% single-use solution
C0359987|Cocaine hydrochloride 10% single-use solution (product)
C0359987|Cocaine hydrochloride 10% single-use solution (substance)
C0359986|Cocaine hydrochloride 2.5% single-use solution
C0359986|Cocaine hydrochloride 2.5% single-use solution (product)
C0359986|Cocaine hydrochloride 2.5% single-use solution (substance)
C0359958|Cocaine / homatropine
C0359958|Cocaine+homatropine
C0359958|Cocaine+homatropine (product)
C0359958|Cocaine+homatropine (substance)
C0975796|Cocaine Hydrochloride 100 MG/ML Topical application Solution
C0975796|Cocaine Hydrochloride 10% Topical solution
C0975796|Cocaine HCl Soln 10%
C0975796|COCAINE HCL 10% SOLN,TOP
C0975796|COCAINE HCL 10% SOLN,TOP [VA Product]
C0975796|COCAINE HCL 10% TOP SOLN
C0975796|Cocaine Hydrochloride 100 MG/ML Topical Solution
C0975796|COCAINE HYDROCHLORIDE 100 mg in 1 mL TOPICAL SOLUTION
C0975796|Cocaine hydrochloride 10% topical solution (product)
C0975796|cocaine HCl 10 % Topical Solution
C0975796|Cocaine viscous 10% topical solution (product)
C0975796|Cocaine viscous 10% topical solution
C0975796|Cocaine Hydrochloride, 10% topical solution
C0975796|cocaine topical 10% topical solution
C0975798|Cocaine Hydrochloride 40 MG/ML Topical application Solution
C0975798|Cocaine Hydrochloride 4% Topical solution
C0975798|Cocaine HCl Soln 4%
C0975798|COCAINE HCL 4% SOLN,TOP
C0975798|COCAINE HCL 4% SOLN,TOP [VA Product]
C0975798|Cocaine Hydrochloride 40 MG/ML Topical Solution
C0975798|COCAINE HYDROCHLORIDE 40 mg in 1 mL TOPICAL SOLUTION
C0975798|cocaine hydrochloride 4 % Topical Solution
C0975798|Cocaine hydrochloride 4% topical solution (product)
C0975798|COCAINE HCL 4% TOP SOLN
C0975798|Cocaine viscous 4% topical solution (product)
C0975798|Cocaine viscous 4% topical solution
C0975798|Cocaine Hydrochloride, 4% topical solution
C0975798|cocaine topical 4% topical solution
C0359957|Cocaine / Epinephrine
C0359957|Cocaine+adrenaline
C0359957|Cocaine+epinephrine (product)
C0359957|Cocaine+epinephrine
C0359957|Cocaine+adrenaline (product)
C0359957|Cocaine+adrenaline (substance)
C0565790|Cocaine - non-pharmaceutical
C0565790|Cocaine - non-pharmaceutical (substance)
C1644725|Cocaine - pharmaceutical (substance)
C1644725|Cocaine - pharmaceutical
C0072534|pseudococaine
C0075888|8-Azabicyclo(3.2.1)octane-2-carboxylic acid, 3-(benzoyloxy)-8-methyl-, methyl ester, (1R-(exo,exo))-, mixt. with 2-(dimethylamino)ethyl 4-(butylamino)benzoate and (R)-4-(1-hydroxy-2-(methylamino)ethyl)-1,2-benzenediol
C0075888|TAC combination
C0075888|TEC solution
C0621633|Baker's cocktail
C0621633|aluminum hydroxide - cimetidine - cocaine - hydroxyzine - morphine
C0621633|aluminum hydroxide, cimetidine, cocaine, hydroxyzine, morphine drug combination
C0621633|Baker's mixture
C0053928|Bonain's liquid
C0056054|cocaine-dipicrylaminate
C0056054|cocaine - dipicrylaminate
C0056054|cocaine, dipicrylaminate drug combination
C0757327|cocaine benzoyl thioester
C0770042|ecgonidine
C1827575|Morphine + cocaine
C1827575|Morphine + cocaine (product)
C1827575|Cocaine + Morphine
C0009950|Convulsants
C0009950|convulsant
C0006644|Caffeine
C0006644|1H-Purine-2,6-dione, 3,7-dihydro-1,3,7-trimethyl-
C0006644|1,3,7-trimethylxanthine
C0006644|3,7-Dihydro-1,3,7-trimethyl-1H-purine-2,6-dione
C0006644|CAF
C0006644|Caffeine product
C0006644|caffeine (medication)
C0006644|caffeine as diuretic (medication)
C0006644|caffeine as diuretic
C0006644|Caffeine [Chemical/Ingredient]
C0006644|Methyltheobromine
C0006644|Theine
C0006644|Trimethylxanthine
C0006644|Caffeine (product)
C0006644|Caffeine (substance)
C0006644|Caffeine, NOS
C0006644|Caffeine product (product)
C0006644|Caffeine product (substance)
C0025810|Methylphenidate
C0025810|2-Piperidineacetic acid, alpha-phenyl-, methyl ester
C0025810|alpha-Phenyl-2-piperidineacetic Acid Methyl Ester
C0025810|Methylphenidate [Chemical/Ingredient]
C0025810|methylphenidate (medication)
C0025810|cns stimulants methylphenidate
C0025810|Methylphenidate (product)
C0025810|Methylphenidate (substance)
C0025810|d-methylphenidate
C0031890|Picrotoxin
C0031890|3,6-Methano-8H-1,5,7-trioxacyclopenta(ij)cycloprop(a)azulene-4,8(3H)-dione, hexahydro-2a-hydroxy-9-(1-hydroxy-1-methylethyl)-8b-methyl-, (1aR-(1aalpha,2abeta,3beta,6beta,6abeta,8aS*,8bbeta,9S*))-, compd. with (1aR-(1aalpha,2abeta,3beta,6beta,6abeta,8aS*,8bbeta,9R*))-hexahydro-2a-hydroxy-8b-methyl-9-(1-methylethenyl)-3,6-methano-8H-1,5,7-trioxacyclopenta(ij)cycloprop(a)azulene-4,8(3H)-dione (1:1)
C0031890|3,6-Methano-8H-1,5,7-trioxacyclopenta(ij)cycloprop(a)azulene-4,8(3H)-dione, hexahydro-2a-hydroxy-9-(1-hydroxy-1-methylethyl)-8b-methyl-, (1aR-(1aalpha,2abeta,3beta,6beta,6abeta,8aS*,8bbeta,9S*))-, compd. with (1aR-(1aalpha,2abeta,3beta,6beta,6abeta,8aS*,8
C0031890|Picrotoxin [Chemical/Ingredient]
C0031890|Picrotoxin (substance)
C0039763|Theobromine
C0039763|1H-Purine-2,6-dione, 3,7-dihydro-3,7-dimethyl-
C0039763|theobromine (medication)
C0039763|vasodilators general theobromine
C0039763|Theobromine [Chemical/Ingredient]
C0039763|3,7-Dimethylxanthine
C0039763|3,7-Dihydro-3,7-Dimethyl-1H-Purine-2,6-Dione
C0039763|Theobromine (substance)
C0002658|Amphetamine
C0002658|dl-Amphetamine
C0002658|Benzeneethanamine, alpha-methyl-, (+-)-
C0002658|Desoxynorephedrine
C0002658|Amfetamine
C0002658|amphetamine (medication)
C0002658|Phenopromin
C0002658|Amphetamine [Chemical/Ingredient]
C0002658|Desoxynorephedrin
C0002658|Phenamine
C0002658|Amphetamine (substance)
C0002658|1-phenylpropan-2-amine
C0002658|d,1-alpha- Methylphenethylamine
C0002658|Phenylaminopropane
C0002658|dl-alpha-methylphenethylamine
C0002658|1-phenylpropan-2-amine (substance)
C0002658|cns stimulants amphetamine (medication)
C0002658|cns stimulants amphetamine
C0002658|Amphetamine (product)
C0002658|Amphetamine, NOS
C0002658|Amphetamine [dup] (substance)
C0002658|Amphetamine (dl-)
C0009014|Clonidine
C0009014|1H-Imidazol-2-amine, N-(2,6-dichlorophenyl)-4,5-dihydro-
C0009014|N-(2,6-Dichlorophenyl)-4,5-dihydro-1H-imidazol-2-amine
C0009014|clonidine (medication)
C0009014|Clonidine [Chemical/Ingredient]
C0009014|Klofenil
C0009014|Clofenil
C0009014|Clonidine (product)
C0009014|Clonidine (substance)
C0024977|Mazindol
C0024977|3H-Imidazo(2,1-a)isoindol-5-ol, 5-(4-chlorophenyl)-2,5-dihydro-
C0024977|mazindol (discontinued) (medication)
C0024977|mazindol (discontinued)
C0024977|anorexics mazindol (discontinued)
C0024977|Mazindole
C0024977|Mazindol [Chemical/Ingredient]
C0024977|Mazindol (product)
C0024977|Mazindol (substance)
C0028128|Monoxide, Nitrogen
C0028128|Nitrate Vasodilator, Endogenous
C0028128|Nitric Oxide
C0028128|Oxide, Nitric
C0028128|Vasodilator, Endogenous Nitrate
C0028128|Endothelium-Derived Nitric Oxide
C0028128|Nitric Oxide, Endothelium Derived
C0028128|Nitrogen oxide (NO)
C0028128|endothelial cell derived relaxing factor
C0028128|Nitric oxide gas
C0028128|Monoxide, Mononitrogen
C0028128|vasodilators pulmonary nitric oxide
C0028128|nitric oxide (medication)
C0028128|Mononitrogen Monoxide
C0028128|Nitric Oxide, Endothelium-Derived
C0028128|Endogenous Nitrate Vasodilator
C0028128|Nitric Oxide [Chemical/Ingredient]
C0028128|Nitrogen Monoxide
C0028128|EDRF
C0028128|NO
C0028128|Nitrogen Oxide
C0028128|NO - Nitric oxide
C0028128|Nitric oxide (substance)
C0028128|Nitric oxide (product)
C0028128|Endothelium-Derived Relaxing Factor
C0030511|Parasympathetic Blocking Agents
C0030511|Parasympatholytics
C0030511|Agents, Parasympathetic-Blocking
C0030511|Agents, Parasympatholytic
C0030511|Drugs, Parasympatholytic
C0030511|PARASYMPATHETIC BLOCK AGENTS
C0030511|parasympatholytic agent
C0030511|[AU350] PARASYMPATHOLYTICS
C0030511|Parasympatholytic
C0030511|Parasympatholytic (product)
C0030511|Parasympatholytic agents
C0030511|Parasympathetic-Blocking Agents
C0030511|Parasympatholytic Drugs
C0030511|Parasympatholytic drug
C0030511|Parasympatholytic drug, NOS
C0030511|Parasympatholytic (substance)
C0030800|Pemoline
C0030800|4(5H)-Oxazolone, 2-amino-5-phenyl-
C0030800|2-Imino-4-keto-5-phenyltetrahydrooxazole
C0030800|5-Phenylisohydantion
C0030800|pemoline (medication)
C0030800|Pemoline [Chemical/Ingredient]
C0030800|Phenoxazole
C0030800|Phenylisohydantoin
C0030800|PIO
C0030800|Pemoline (product)
C0030800|Pemoline (substance)
C0030903|Pentylenetetrazole
C0030903|5H-Tetrazolo(1,5-a)azepine, 6,7,8,9-tetrahydro-
C0030903|PTZ
C0030903|pentylenetetrazol
C0030903|pentylenetetrazol (medication)
C0030903|Leptazole
C0030903|Pentetrazole
C0030903|Pentylenetetrazole [Chemical/Ingredient]
C0030903|Pentamethylenetetrazole
C0030903|Pentetrazol
C0030903|Pentylenetetrazol (substance)
C0030903|Pentylenetetrazol [dup] (substance)
C0043318|Xanthines
C0043318|xanthines (medication)
C0043318|Xanthines [Chemical/Ingredient]
C0031974|pipradrol
C0031974|pyridrol
C0031974|pipradol
C0031974|Pipradrol (substance)
C0701400|Nicorette
C0028040|Nicotine
C0028040|Pyridine, 3-(1-methyl-2-pyrrolidinyl)-, (S)-
C0028040|beta-Pyridyl-alpha-N-methylpyrrolidine
C0028040|(S)-3-(1-Methyl-2-pyrrolidinyl)pyridine
C0028040|1-Methyl-2-(3-pyridyl)pyrrolidine
C0028040|NIC
C0028040|Nicotine product
C0028040|nicotine (medication)
C0028040|Nicotine [Chemical/Ingredient]
C0028040|(-)-Nicotine
C0028040|Nicotine - chemical
C0028040|Nicotine (product)
C0028040|Nicotine (substance)
C0028040|Nicotine agent (substance)
C0028040|Nicotine agent
C0028040|Nicotine product (product)
C0028040|Nicotine product (substance)
C0733634|AN448
C0733634|AN-448
C0030802|Magnesium, Pemoline
C0030802|Pemoline Magnesium
C0031977|Piracetam
C0031977|1-Pyrrolidineacetamide, 2-oxo-
C0031977|Piracetam [Chemical/Ingredient]
C0031977|Pirazetam
C0031977|Pyramem
C0031977|2-Pyrrolidone-N-Acetamide
C0031977|Pyracetam
C0031977|piracetam (medication)
C0031977|Piracetam (product)
C0031977|Piracetam (substance)
C0004960|Bemegride
C0004960|2,6-Piperidinedione, 4-ethyl-4-methyl-
C0004960|Methetharimide
C0004960|Bemegride [Chemical/Ingredient]
C0004960|Ethylmethylglutarimide
C0004960|Bemegride (substance)
C0005096|Benzphetamine
C0005096|Benzeneethanamine, N,alpha-dimethyl-N-(phenylmethyl)-, (S)-
C0005096|Benzphetamine [Chemical/Ingredient]
C0005096|Benzfetamine
C0005096|Benzphetamine (product)
C0005096|Benzphetamine (substance)
C0011812|Dextroamphetamine
C0011812|d Amphetamine
C0011812|d-Amphetamine
C0011812|dextro Amphetamine
C0011812|Benzeneethanamine, alpha-methyl-, (S)-
C0011812|AMPHETAMINE A D
C0011812|(+)-Amphetamine
C0011812|Dextroamphetamine [Chemical/Ingredient]
C0011812|Dexamfetamine
C0011812|Dexamphetamine
C0011812|dextro-Amphetamine
C0011812|Dexamfetamine (substance)
C0011812|psychostimulants dextroamphetamine
C0011812|dextroamphetamine (medication)
C0011812|Dextroamphetamine (product)
C0011812|Dextroamphetamine (substance)
C0011812|Amphetamine (d-)
C0013084|Doxapram
C0013084|2-Pyrrolidinone, 1-ethyl-4-(2-(4-morpholinyl)ethyl)-3,3-diphenyl-
C0013084|Doxapram [Chemical/Ingredient]
C0013084|Doxapram (product)
C0013084|Doxapram (substance)
C0014479|Ephedrine
C0014479|[R-(R*,S*)]-alpha-[1-(Methylamino)ethyl]benzenemethanol
C0014479|(-)-Ephedrine
C0014479|(1R,2S)-2-methylamino-1-phenyl-propan-1-ol
C0014479|Ephedrine Erythro Isomer
C0014479|ephedrine (medication)
C0014479|Ephedrine [Chemical/Ingredient]
C0014479|Erythro Isomer of Ephedrine
C0014479|antiasthmatics ephedrine (medication)
C0014479|antiasthmatics ephedrine
C0014479|Ephedrine (product)
C0014479|Ephedrine (substance)
C0018602|Harmaline
C0018602|3H-Pyrido(3,4-b)indole, 4,9-dihydro-7-methoxy-1-methyl-
C0018602|Harmaline [Chemical/Ingredient]
C0018602|Dihydroharmine
C0018602|Harmidine
C0018602|Harmaline (substance)
C0025611|Methamphetamine
C0025611|N Methylamphetamine
C0025611|Benzeneethanamine, N,alpha-dimethyl-, (S)-
C0025611|Desoxyephedrine
C0025611|deoxyephedrine
C0025611|decongestants desoxyephedrine
C0025611|desoxyephedrine (medication)
C0025611|methamphetamine preparations
C0025611|anorexics amphetamines methamphetamine preparations
C0025611|methamphetamine preparations (medication)
C0025611|Metamfetamine
C0025611|Methamphetamine [Chemical/Ingredient]
C0025611|Methylamphetamine
C0025611|N-Methylamphetamine
C0025611|Speed
C0025611|Tina
C0025611|Ice
C0025611|Glass
C0025611|Crystal
C0025611|Chalk
C0025611|Meth
C0025611|Desoxyephedrine (substance)
C0025611|anorexics amphetamines methamphetamine
C0025611|methamphetamine (medication)
C0025611|Methamphetamine (product)
C0025611|Methamphetamine (substance)
C0028089|Diethylamide, Nicotinic
C0028089|Nikethamide
C0028089|3-Pyridinecarboxamide, N,N-diethyl-
C0028089|nikethamide (medication)
C0028089|Corethamid
C0028089|Nicotinic Diethylamide
C0028089|Nizethamid
C0028089|Nicethamide
C0028089|Nikethamide [Chemical/Ingredient]
C0028089|Diethylnicotinamid
C0028089|Nikethamide (product)
C0028089|Nikethamide (substance)
C0031411|Phenmetrazine
C0031411|Morpholine, 3-methyl-2-phenyl-
C0031411|Fenmetrazin
C0031411|Phenmetraline
C0031411|Oxazimedrine
C0031411|Phenmetrazine [Chemical/Ingredient]
C0031411|Defenmetrazin
C0031411|Phenmetrazine (product)
C0031411|Phenmetrazine (substance)
C0031447|Phentermine
C0031447|Benzeneethanamine, alpha,alpha-dimethyl-
C0031447|Phentermine [Chemical/Ingredient]
C0031447|1,1-Dimethyl-2-phenylethylamine
C0031447|2-Phenyl-tert-butylamine
C0031447|2-Amino-2-methyl-1-phenylpropane
C0031447|Phenyl-tertiary-butylamine
C0031447|Phentermine (product)
C0031447|Phentermine (substance)
C0003567|Aphrodisiacs
C0003567|Aphrodisiac (substance)
C0003567|Aphrodisiac
C0003567|Aphrodisiac, NOS
C0376447|Appetite Stimulants
C0376447|Appetite Stimulating Drugs
C0376447|Drugs, Appetite-Stimulating
C0376447|Stimulants, Appetite
C0376447|Appetite-Stimulating Drugs
C0002763|Central Nervous System Stimulants
C0002763|Stimulants, Central
C0002763|CNS stimulant
C0002763|CNS STIMULANTS
C0002763|central nervous system stimulant
C0002763|central nervous system stimulants (medication)
C0002763|Analeptic Agent
C0002763|Analeptics
C0002763|[CN800] CNS STIMULANTS
C0002763|Stimulants
C0002763|stimulant
C0002763|Central Stimulants
C0002763|Central stimulant
C0002763|Central stimulant (product)
C0002763|Central stimulant (substance)
C0002763|Central nervous system stimulant, NOS
C0002763|Central stimulant, NOS
C0002763|CNS Stimulating Drugs
C0002763|Stimulants of CNS
C0012201|Diethylpropion
C0012201|1-Propanone, 2-(diethylamino)-1-phenyl-
C0012201|Amfepramone
C0012201|2-Diethylaminopropiophenone
C0012201|Diethylpropion [Chemical/Ingredient]
C0012201|Amfepramon
C0012201|Phepranon
C0012201|Diethylpropion (product)
C0012201|Diethylpropion (substance)
C0795571|AMPHETAMINE/DEXTROAMPHETAMINE
C0795571|amphetamine + dextroamphetamine (medication)
C0795571|anorexics amphetamine + dextroamphetamine
C0795571|amphetamine + dextroamphetamine
C0795571|amphetamine-dextroamphetamine
C0795571|Amphetamine / Dextroamphetamine
C0795571|dextroamphetamine-amphetamine
C0795571|SLI381
C0795571|D,L-amphetamine
C0795571|Amphetamine+dextroamphetamine (product)
C0795571|Amphetamine+dextroamphetamine
C0066677|benzhydrylsulfinylacetamide
C0066677|modafinil
C0066677|modafinil (medication)
C0066677|modafinil [Chemical/Ingredient]
C0066677|2-((diphenylmethyl)sulfinyl)acetamide
C0066677|Modafinil (product)
C0066677|Modafinil (substance)
C0994515|7-acetyl-5-(4-aminophenyl)-8,9-dihydro-8-methyl-7H-1,3-dioxolo(4,5-h)benzodiazepine
C0994515|(R)-(-)-1-(4-Aminophenyl)-3-acetyl-4-methyl-7,8-methylenedioxy-3,4-dihydro-5H-2,3-benzodiazepine
C0994515|talampanel
C0994515|1-(4'-aminophenyl)-3-acetyl-4-methyl-3,4-dihydro-7,8-methylenedioxy-5H-2,3-benzodiazepine
C0282133|Diethylpropion Hydrochloride
C0282133|Hydrochloride, Diethylpropion
C0282133|1-phenyl-2-diethyl-amino-1-propanone Hydrochloride
C0282133|anorexics diethylpropion hydrochloride
C0282133|diethylpropion hydrochloride (medication)
C0282133|Diethylpropion Hydrochloride [Chemical/Ingredient]
C0282133|Diethylpropion hydrochloride (substance)
C0282133|Diethylpropion hydrochloride (product)
C0282133|Amfepramone hydrochloride
C0282133|Diethylpropion hydrochloride [dup] (substance)
C0767825|Irampanel
C0767825|dimethyl-(2-(2-(3-phenyl-(1,2,4)oxadiazol-5-yl)phenoxy)ethyl)amine hydrochloride
C0767825|5-(o-(2-(Dimethylamino)ethoxy)phenyl)-3-phenyl-1,2,4-oxadiazole
C1565316|(S)-N-(2-(1,6,7,8-tetrahydro-2H-indeno-(5,4)furan-8-yl)ethyl)propionamide
C1565316|ramelteon
C1565316|ramelteon (medication)
C1565316|ramelteon [Chemical/Ingredient]
C1565316|Ramelteon (product)
C1565316|Ramelteon (substance)
C2699993|Endomide
C2698084|Amfetaminil
C0051684|2,4-diamino-5-phenylthiazole
C0051684|amiphenazole
C0051684|Amiphenazole (substance)
C0034295|Pyrithioxin
C0034295|pyritinol (medication)
C0034295|pyritinol
C0034295|4-Pyridinemethanol, 3,3'-(dithiobis(methylene))bis(5-hydroxy-6-methyl- )
C0034295|Pyrithioxin [Chemical/Ingredient]
C0034295|Pyrithioxine
C0034295|Piritinol
C0034295|Dipyridoxolyldisulfide
C0034295|Pyridoxinedisulfide
C0034295|Pyritinol (substance)
C2700197|Flubanilate
C0002164|Almitrine
C0002164|1,3,5-Triazine-2,4-diamine, 6-(4-(bis(4-fluorophenyl)methyl)-1-piperazinyl)-N,N'-di-2-propenyl-
C0002164|2,4-Bis(allylamino)-6-(4-(bis(p-fluorophenyl)methyl)-1-piperazinyl)-s-triazine
C0002164|Almitrin
C0002164|Almitrine [Chemical/Ingredient]
C0002164|Almitrine (substance)
C2699299|Sibopirdine
C2698764|Perampanel
C2698764|3-(2-cyanophenyl)-5-(2-pyridyl)-1-phenyl-1,2-dihydropyridin-2-one
C2698764|perampanel (medication)
C2698764|anticonvulsants perampanel
C2698764|Perampanel (substance)
C2698764|Perampanel (product)
C2698764|E2007
C2698764|Benzonitrile, 2-(1',6'-Dihydro-6'-oxo-1'-phenyl(2,3'-bipyridin)-5'-yl)-
C0068978|cafedrine
C0068978|norephendrinetheophylline
C0068978|7-(2-(1-methyl-2-hydroxy-2-phenylethylamino)ethyl)theophylline
C2699227|Cinoxopazide
C2698105|Ampyzine Sulfate
C0056852|cyprodenate
C0056852|dimethylamino- 2-ethyl-beta-cyclohexylpropionic acid maleate
C0056852|cyprodemanol
C2699566|Deanol Aceglumate
C0057219|2-(dimethylamino)ethanol p-acetamidobenzoate
C0057219|deanol acetamidobenzoate
C2699617|Dextroamphetamine Phosphate
C0059692|etamivan
C0059692|ethamivan
C0059692|Ethamivan (product)
C0059692|Ethamivan (substance)
C0016380|Flurothyl
C0016380|Flurotyl
C0016380|Ethane, 1,1'-oxybis(2,2,2-trifluoro)-
C0016380|Fluorothyl
C0016380|Flurothyl [Chemical/Ingredient]
C0016380|Hexafluorodiethyl ether
C0016380|Flurothyl (substance)
C0016380|Flurothyl [dup] (substance)
C2698810|Pimeclone
C0071957|prethcamide
C1739826|lisdexamfetamine dimesylate
C1739826|Lisdexamfetamine dimesylate (substance)
C1739826|lisdexamfetamine dimesylate (medication)
C1739826|Dimesylate, Lisdexamfetamine
C1739826|Dimesylate, Lis-dexamfetamine
C1739826|Lis dexamfetamine Dimesylate
C1739826|Lisdexamfetamine Dimesylate [Chemical/Ingredient]
C1739826|Lis-dexamfetamine Dimesylate
C1999336|tezampanel
C1999336|(3S,4aR,6R,8aR)-6-(2-(1H-Tetrazol-5-yl)ethyl)decahydroisoquinoline-3-carboxylic Acid Monohydrate
C0050407|aceglutamide
C0050407|N-acetyl-L-glutamine
C0050407|N-acetylglutamine
C2698101|Amphetamine Hydrochloride
C2699365|Clofenciclan
C2699618|Dextrofemine
C2698336|Becampanel
C2698336|((7-Nitro-2,3-dioxo-1,2,3,4-tetrahydroquinoxalin-5-yl)methylamino)methylphosphonic Acid
C2698104|Ampyzine
C2698056|Almitrine Mesylate
C2698056|1,3,5-Triazine-2,4-diamine, 6-(4-(bis(4-fluorophenyl)methyl)-1-piperazinyl)-N,N'-di-2-propenyl-, Dimethanesulfonate
C0000379|3,4 Methylenedioxyamphetamine
C0000379|3,4-Methylenedioxyamphetamine
C0000379|MDA
C0000379|1,3-Benzodioxole-5-ethanamine, alpha-methyl-
C0000379|METHYLENEDIOXYAMPHETAMINE 03 04
C0000379|Alpha-Methyl-1,3-benzodioxole-5-ethanamine
C0000379|Tenamfetamine
C0000379|Methylenedioxyamphetamine
C0000379|3,4-Methylenedioxyamphetamine [Chemical/Ingredient]
C0000379|Methylenedioxyamphetamine (substance)
C2699925|(3S,4aR,6R,8aR)-6-(2-(1H-Tetrazol-5-yl)ethyl)decahydroisoquinoline-3-carboxylic Acid Monohydrate Anhydrous
C2699925|Tezampanel Anhydrous
C0058252|dimephenopan
C0058252|dimethylamphetamine
C0058252|N,N,alpha-trimethylbenzeneethanamine
C0058252|N,N,alpha-trimethylphenethylamine
C0058252|N,N-dimethylamphetamine
C0058252|Dimetamfetamine
C0058252|Dimethamphetamine
C0058252|(S)-N,N,alpha-Trimethylphenethylamine
C0058252|Dimethamphetamine (product)
C0058252|Dimethamphetamine (substance)
C0058252|N-methyl-methamphetamine
C0072127|1-(alpha-propylphenethyl)pyrrolidine
C0072127|phenylpyrrolidinylpentan
C0072127|prolintane
C0072127|Prolintane (product)
C0072127|Prolintane (substance)
C0070549|phendimetrazine
C0070549|phendimetrazine [Chemical/Ingredient]
C0070549|(2S,3S)-3,4-Dimethyl-2-Phenylmorpholine
C0070549|Morpholine, 3,4-Dimethyl-2-Phenyl-, (2s-Trans)-
C0070549|Phendimetrazine (product)
C0070549|Phendimetrazine (substance)
C0289432|Methylergonovine Maleate
C0289432|Ergoline-8-carboxamide, 9,10-didehydro-N-((1S)-1-(hydroxymethyl)propyl)-6-methyl-,(8beta)-,(2Z)-2-butenedioate(1:1)(salt)
C0289432|Maleic Acid, Methyl Ergonovine
C0289432|methylergonovine maleate (medication)
C0289432|oxytocics methylergonovine maleate
C0289432|Methylergonovine Maleate [Chemical/Ingredient]
C0289432|Methylergometrine Maleate
C0289432|Methylergometrine maleate preparation
C0289432|Methylergonovine maleate preparation
C0289432|Methylergonovine maleate (substance)
C0289432|Methylergonovine maleate preparation (product)
C0289432|Methylergonovine maleate preparation (substance)
C0724568|Dextroamphetamine Saccharate
C0724568|dextroamphetamine saccharate (medication)
C0724568|Dextroamphetamine saccharate (product)
C0724568|Dexamfetamine saccharate
C0724568|Dextroamphetamine saccharate (substance)
C0025760|Methylergonovine
C0025760|Ergoline-8-carboxamide, 9,10-didehydro-N-(1-(hydroxymethyl)propyl)-6-methyl-, (8beta(S))-
C0025760|Methylergonovine [Chemical/Ingredient]
C0025760|Methylergometrine
C0025760|Methylergobasin
C0025760|Methylergometrin
C0025760|Methylergometrine preparation
C0025760|Methylergonovine preparation
C0025760|Methylergonovine (substance)
C0025760|Methylergonovine preparation (product)
C0025760|Methylergonovine preparation (substance)
C2825427|Camphramine
C2825427|Camphotamide
C2825428|Cyclazodone
C0059791|ethylamphetamine
C0059791|Etilamfetamine
C0059791|N-ethylamphetamine
C0060167|7-(2-((alpha-methylphenethyl)amino)ethyl)theophylline
C0060167|7-ethyltheophyllineamphetamine
C0060167|fenethylline
C0060167|fenetylline
C0060167|Theophylline ethylamphetamine
C0060167|Fenethylline (substance)
C2825430|Fenethylline Hydrochloride
C0064875|levophacetoperane
C0064875|Levofacetoperane
C2826074|Zylofuramine
C0301388|2-Amino-1,1-diphenylheptamol
C0301388|Hexapradol
C0301388|Alpha-(1-Aminohexyl)benzhydrol
C0301388|Hexapradol (substance)
C0771352|CAFFEINE MONOHYDRATE
C0771352|1,3,7-Trimethyl-3,7-Dihydro-1H-Purine-2,6-Dione Monohydrate
C2827094|Calcium Hopantenate Anhydrous
C0219131|Hexacyclonate Sodium
C0219131|1-(hydroxymethyl)cyclohexaneacetic acid, sodium salt
C2827167|Hexacyclonic Acid
C2827167|Hexacyclonate
C2827167|Cyclohexaneacetic Acid, 1-(Hydroxymethyl)-
C2827167|1-(Hydroxymethyl)Cyclohexaneacetate
C0072777|4'-methyl-2-(1-pyrrolidinyl)valerophenone
C0072777|pyrovalerone
C0072777|1-(4-methylphenyl)-2-pyrrolidin-1-yl-pentan-1-one
C0072777|Pyrovalerone (substance)
C0066048|2-(dimethylamino)propiophenone
C0066048|dimepropion
C0066048|dimethylpropion
C0066048|metamfepramone
C0982017|Amphetamine Adipate
C0108116|calcium hopantenate
C0108116|Calcium Homopantothenate
C0108116|Hopantenate Calcium
C0108116|Hopantenic Acid, Calcium Salt Hemihydrate
C0108116|Calcium D-(+)-4-(2,4-Dihydroxy-3,3-Dimethylbutylamido)Butyrate Hemihydrate
C1170743|Dexmethylphenidate Hydrochloride
C1170743|d-threo-Methylphenidate Hydrochloride
C1170743|2-Piperidineacetic Acid, Alpha-phenyl-, Methyl Ester, Hydrochloride, (alphaR,2R)-
C1170743|dexmethylphenidate hydrochloride (medication)
C1170743|Hydrochloride, Dexmethylphenidate
C1170743|Dexmethylphenidate Hydrochloride [Chemical/Ingredient]
C1170743|Dexmethylphenidate hydrochloride (substance)
C0010725|5'-Diphosphocholine, Cytidine
C0010725|Choline, CDP
C0010725|Choline, Cytidine Diphosphate
C0010725|Cytidine Diphosphate Choline
C0010725|Diphosphate Choline, Cytidine
C0010725|Cytidine 5' Diphosphocholine
C0010725|Cytidine 5'-(trihydrogen diphosphate), P'-(2-(trimethylammonio)ethyl) ester, inner salt
C0010725|citicoline (medication)
C0010725|citicoline
C0010725|Cytidine Diphosphate Choline [Chemical/Ingredient]
C0010725|Cyticholine
C0010725|CDP Choline
C0010725|Citicholine
C0010725|Cidifos
C0010725|Cytidine 5'-Diphosphocholine
C0010725|CDP-choline
C0010725|Cytidine 5-diphosphocholine
C0010725|Cytidine 5'-(trihydrogen Diphosphate), Mono(2-(trimethylammonio)ethyl) Ester, Hydroxide, Inner Salt
C0010725|Citicoline (substance)
C0123163|idebenone
C0123163|Idebenone (product)
C0123163|Idebenone (substance)
C0123163|idebenone (medication)
C0123163|hydroxydecyl ubiquinone
C0123163|noben
C2047880|idebenone + vitamin E (medication)
C2047880|idebenone + vitamin E
C2047880|idebenone / Vitamin E
C2194148|fencamfamine + vitamins (medication)
C2194148|fencamfamine + vitamins
C2081457|pipradrol + B1 + B2 + B3 + B6 + choline + inositol
C2081457|pipradrol + thiamine + riboflavin + niacin + pyridoxine + choline + inositol (medication)
C2081457|pipradrol + thiamine + riboflavin + niacin + pyridoxine + choline + inositol
C2081458|pipradrol + vitamins + minerals
C2081458|pipradrol + vitamins + minerals (medication)
C0771021|prolintane hydrochloride
C0771021|prolintane hydrochloride (medication)
C1701455|Armodafinil
C1701455|Armodafinil (product)
C1701455|Armodafinil (substance)
C1701455|(-)-2-((R)-(Diphenylmethyl)sulfinyl)acetamide
C1701455|2-((R)-(diphenylmethyl)sulfinyl)acetamide
C1701455|armodafinil (medication)
C1701455|cns stimulants armodafinil
C0068722|nicotine polacrilex
C0068722|nicotine polacrilex (medication)
C0068722|nicotine polacrilex [Chemical/Ingredient]
C0068722|Nicotine Polacrilices
C0068722|Polacrilex, Nicotine
C0068722|Polacrilices, Nicotine
C0068722|Nicotine polacrilex (substance)
C0358855|Nicotine Transdermal Patch
C0358855|nicotine patch
C0358855|nicotine transdermal patch (medication)
C0358855|Patch, Nicotine Transdermal
C0358855|Transdermal Patch, Nicotine
C0358855|Patch, Nicotine
C0358855|Nicotine m/r transdermal patch (product)
C0358855|Nicotine m/r transdermal patch
C0358855|Nicotine patches
C0358855|Nicotine patches (product)
C0358855|Nicotine patches (substance)
C0358855|Nicotine Skin Patch
C0002667|Amphetamines
C0002667|amphetamines (medication)
C0002667|anorexics amphetamines
C0002667|[CN801] AMPHETAMINES
C0002667|Amphetamines [Chemical/Ingredient]
C0002667|Amphetamine
C0002667|Amphetamine group
C0002667|Amfetamine group
C1874222|AMPHETAMINE LIKE STIMULANTS
C1874222|[CN802] AMPHETAMINE LIKE STIMULANTS
C0731742|Other central nervous system stimulants
C0731742|CNS STIMULANTS,OTHER
C0731742|[CN809] CNS STIMULANTS,OTHER
C0731742|Other central nervous system stimulants (product)
C0731742|Other central nervous system stimulants (substance)
C2981334|Famiraprinium
C2981334|6-Amino-1-(3-Carboxypropyl)-5-Methyl-3-Phenylpyridazinium
C0916220|Picrotin
C0042674|Vincamine
C0042674|Eburnamenine-14-carboxylic acid, 14,15-dihydro-14-hydroxy-, methyl ester, (3alpha,14beta,16alpha)-
C0042674|Vincamine [Chemical/Ingredient]
C0042674|Vincamine (substance)
C0301353|Alpha-Methyl-N-(2,2,2-Trichloroethylidene)Phenethylamine
C0301353|Amphecloral
C0301353|Amfecloral
C0301353|Benzeneethanamine, Alpha-Methyl-N-(2,2,2-Trichloroethylidene)-
C0301353|Amphechloral
C0301353|Amphechloral (substance)
C0301353|Amfecloral (substance)
C0051574|7-benzyl-1-ethyl-1,4-dihydro-4-oxo-1,8-naphthyridine-3-carboxylic acid
C0051574|amfonelic acid
C2983904|Methamphetamine, DL-
C2987049|(-)-Amphetamine Sulfate
C2987049|Levamphetamine Sulphate
C2987049|L-Amphetamine Sulfate
C2987049|L-Amphetamine Sulphate
C2987049|Benzeneethanamine, Alpha-Methyl-, (R)-, Sulphate (2:1)
C2987049|(-)-Amphetamine Sulphate
C2987049|Levamfetamine Sulfate
C2987049|Levamphetamine Sulfate
C0000477|4 Aminopyridine
C0000477|4-Aminopyridine
C0000477|4-Pyridinamine
C0000477|FAMPRIDINE (4-AMINOPYRIDINE)
C0000477|AMINOPYRIDINE 04
C0000477|FAMPRIDINE
C0000477|dalfampridine
C0000477|Pymadine
C0000477|4-Aminopyridine [Chemical/Ingredient]
C0000477|4-AP
C0000477|dalfampridine (medication)
C0000477|cns stimulants dalfampridine
C0000477|4-Aminopyridine (substance)
C0000477|4-Aminopyridine (product)
C0011064|Deanol
C0011064|Ethanol, 2-(dimethylamino)-
C0011064|N,N Dimethyl 2 hydroxyethylamine
C0011064|Dimethylethanolamine
C0011064|Dimethyl ethanolamine
C0011064|parasympathomimetics deanol
C0011064|deanol (medication)
C0011064|N,N-Dimethyl-N-(2-hydroxyethyl)amine
C0011064|2-Dimethylaminoethanol
C0011064|Dimethylaminoethanol
C0011064|Demanyl
C0011064|Demanol
C0011064|N,N-Dimethyl-2-hydroxyethylamine
C0011064|N,N-Dimethylethanolamine
C0011064|Deanol [Chemical/Ingredient]
C0011064|Dimethyl ethanolamine (substance)
C0011064|Deanol (substance)
C0011064|2 Dimethylaminoethanol
C0242181|Analeptics
C0242181|analeptic
C0242181|Agents, Analeptic
C0242181|Drugs, Analeptic
C0242181|Analeptic agent
C0242181|Analeptic agent (substance)
C0242181|Analeptic Drugs
C0242181|Analeptic Agents
C0242181|Analeptic agent (product)
C0242181|Analeptic agent, NOS
C0056512|cropropamide
C0056512|n-(N'-crotonyl-N'-propyl)amino-N,N-dimethylbutyramide
C0056512|Cropropamide (substance)
C0705972|modafinil 200 MG Oral Tablet
C0705972|MODAFINIL 200MG TAB
C0705972|Modafinil Tab 200 MG
C0705972|MODAFINIL 200MG TAB [VA Product]
C0705972|Modafinil 200mg Oral tablet
C0705972|Modafinil, 200 mg oral tablet
C0705972|MODAFINIL 200 mg ORAL TABLET [Modafinil]
C0705972|Modafinil 200mg tablet
C0705972|Modafinil 200mg tablet (product)
C0876575|Pemoline 37.5 MG Oral Tablet
C0876575|Pemoline 37.5mg Oral tablet
C0876575|PEMOLINE 37.5MG TAB
C0876575|PEMOLINE 37.5MG TAB [VA Product]
C0876575|Pemoline, 37.5 mg oral tablet
C0876575|Pemoline 37.5mg tablet (product)
C0876575|Pemoline 37.5mg tablet
C0350544|Weak central nervous system stimulants (product)
C0350544|Weak central nervous system stimulants
C0350544|Weak central nervous system stimulants (substance)
C1591277|Pemoline 18.75 MG Oral Tablet
C1591277|Pemoline 18.8 MG Oral Tablet
C1591277|Pemoline 18.75mg Oral tablet
C1591277|PEMOLINE 18.75MG TAB
C1591277|PEMOLINE 18.75MG TAB [VA Product]
C1591277|Pemoline, 18.75 mg oral tablet
C1591277|Pemoline 18.75mg tablet (product)
C1591277|Pemoline 18.75mg tablet
C0142928|SODIUM SUCCINATE
C0142928|Sodium succinate (substance)
C0060157|2-ethylamino-3-phenylnorcamphane
C0060157|bicyclo(2.2.1)heptan-2-amine, N-ethyl-3-phenyl-
C0060157|fencamfamine
C0060157|N-ethyl-3-phenylbicyclo(2.2.1)heptan-2-amine
C0060157|Fencamfamin
C0060157|2-Norbornanamine, N-Ethyl-3-Phenyl-
C0060157|3-Phenyl-N-Ethyl-2-Norbornanamine
C0060157|2-Phenyl-3-Ethylaminobicyclo(2.2.1)Heptane
C0060157|2-Ethylamino-3-Phenylnorbornane
C0060157|Fencamfamin (substance)
C0056521|crotetamide
C0056521|crotethamide
C0056521|n-(N'-crotonyl-N'-ethyl)amino- N,N-dimethylbutyramide
C0056521|Crotethamide (substance)
C0361631|Drugs used to treat hyperactivity disorders
C0361631|Drugs used to treat hyperactivity disorders (product)
C0361631|Drugs used to treat hyperactivity disorders (substance)
C0689908|Pemoline 75 MG Oral Tablet
C0689908|Pemoline 75mg Oral tablet
C0689908|PEMOLINE 75MG TAB
C0689908|PEMOLINE 75MG TAB [VA Product]
C0689908|Pemoline, 75 mg oral tablet
C0689908|Pemoline 75mg tablet (product)
C0689908|Pemoline 75mg tablet
C0350545|Weak central nervous system stimulant+vitamins (product)
C0350545|Weak central nervous system stimulant+vitamins
C0350545|Weak central nervous system stimulant+vitamins (substance)
C1569608|varenicline
C1569608|Varenicline (product)
C1569608|Varenicline (substance)
C1569608|7,8,9,10-tetrahydro-6,10-methano-6H-pyrazino(2,3-h)(3)benzazepine (2R,3R)-2,3-dihydroxybutqanedioate
C1569608|cns stimulants varenicline
C1569608|varenicline (medication)
C1569608|6,7,8,9-Tetrahydro-6,10-methano-6H-pyrazino(2,3-h)benzazepine
C1569608|Varenicline [Chemical/Ingredient]
C1873633|Lisdexamfetamine
C1873633|Lisdexamfetamine (product)
C1873633|Lisdexamfetamine (substance)
C1873633|lisdexamfetamine (medication)
C1873633|cns stimulants lisdexamfetamine
C3658225|Wake Promoting Drugs
C3658225|Drugs, Wake-Promoting
C3658225|Substances, Wake-Promoting
C3658225|Drugs, Eugeroic
C3658225|Wakefulness-Promoting Agents
C3658225|Agents, Wakefulness-Promoting
C3658225|Wakefulness Promoting Agents
C3658225|Agents, Wake-Promoting
C3658225|Wake Promoting Agents
C3658225|Wake Promoting Substances
C3658225|Eugeroic Drugs
C3658225|Wake-Promoting Drugs
C3658225|Wake-Promoting Substances
C3658225|Wake-Promoting Agents
C0072732|pyrisuccideanol
C0072732|Pirisudanol
C0072732|Pirisudanol (substance)
C1972380|Pyrovalerone &#x7C; urine
C3534074|Methylenedioxypyrovalerone &#x7C; Urine
C1445631|Amphetamine and derivatives (substance)
C1445631|Amphetamine and derivatives
C1169997|dexmethylphenidate
C1169997|Dexmethylphenidate (product)
C1169997|d-MPH
C1320172|Methylphenidate and derivative (substance)
C1320172|Methylphenidate and derivative
C0047392|3-fluorotyrosine
C0047392|meta-fluorotyrosine
C0047392|3-fluoro-tyrosine
C0070743|4-(2-(methylamino)propyl)phenol
C0070743|4-hydroxy-N-methylamphetamine
C0070743|4-hydroxymethamphetamine
C0070743|p-hydroxymethamphetamine
C0070743|pholedrine
C0070743|pulsotyl
C0070743|1-(p-Hydroxyphenyl)-2-methylaminopropane
C0070743|Pholedrine (substance)
C0074500|mesocarb
C0074500|N-phenylcarbamoyl-3-(beta-phenylisopropyl)sydnonimine
C0074500|sidnocarb
C0074500|sydnocarb
C0050672|Actovegin
C0066815|morphine-3-glucuronide
C0054876|1-propanone, 2-amino-1-phenyl
C0054876|2-amino-1-phenyl-1-propanone
C0054876|2-aminopropiophenone
C0054876|alpha-aminopropiophenone
C0054876|cathinine
C0054876|cathinone
C0058222|dimethyl methylphosphonate
C0058222|dimethyl methanephosphonate
C0058222|dimethylmethylphosphonate
C0290795|Adderall
C0011786|Dexfenfluramine
C0011786|Benzeneethanamine, N-ethyl-alpha-methyl-3-(trifluoromethyl)-, (S)-
C0011786|Dexfenfluramine [Chemical/Ingredient]
C0011786|Dexfenfluramine (product)
C0011786|Dexfenfluramine (substance)
C1641209|Central respiratory stimulant (substance)
C1641209|Central respiratory stimulant
C0054436|caffeine citrate
C0054436|Citrated Caffeine
C0054436|caffeine citrated
C0054436|caffeine citrated (medication)
C0054436|caffeine citrate [Chemical/Ingredient]
C0054436|Caffeine citrate (product)
C0054436|Caffeine citrate (substance)
C0054436|Caffeina Citrata
C1881803|Metazide
C0025380|Mephentermine
C0025380|Benzeneethanamine, N,alpha,alpha-trimethyl-
C0025380|Mephentermine [Chemical/Ingredient]
C0025380|Mephentermine (substance)
C0115471|MDMA
C0115471|Ecstasy
C0115471|N Methyl 3,4 methylenedioxyamphetamine
C0115471|N-Methyl-3,4-methylenedioxyamphetamine
C0115471|1,3-Benzodioxole-5-ethanamine, N,alpha-dimethyl-
C0115471|3,4 methylenedioxymethamphetamine
C0115471|MMDA
C0115471|3-Methoxy-4,5- methylenedioxyamphetamine
C0115471|3,4-methylenedioxymethamphetamine
C0115471|METHYLMETHYLENEDIOXYAMPHETAMINE N 03 04
C0115471|Ecstasy - drug
C0115471|Methylene-dioxymethamphetamine
C0115471|ecstasy (drug)
C0115471|Ecstasy - agent
C0115471|N-Methyl-3,4-methylenedioxyamphetamine [Chemical/Ingredient]
C0115471|Methylenedioxymethamphetamine
C0115471|XTC
C0115471|n-Methyl-3, 4-methylenedioxyamphetamine (substance)
C0115471|E - Ecstasy
C0115471|n-Methyl-3, 4-methylenedioxyamphetamine
C0115471|Ecstasy - agent (substance)
C0115471|Methylene-dioxymethamphetamine (substance)
C0115471|MDM
C0115471|MDMA - Methylenedioxymethamphetamine
C0115471|Methylene-dioxymethamphetamine (product)
C0115471|Methylenedioxymethamphetamine (substance)
C0115471|Ecstasy - drug (substance)
C0115471|Methylenedioxymethamfetamine
C0700545|Hydrochloride, Methylphenidate
C0700545|Methylphenidate Hydrochloride
C0700545|alpha-Phenyl-2-piperidineacetic Acid Methyl Ester Hydrochloride
C0700545|methylphenidate hydrochloride (medication)
C0700545|Methylphenidate Hydrochloride [Chemical/Ingredient]
C0700545|Methylphenidylacetate hydrochloride
C0700545|Methylphenidate hydrochloride (substance)
C0700545|Methylphenidate hydrochloride (product)
C0060187|2-ethylamino-5-phenyl-2-oxazolin-4-one
C0060187|fenozolone
C0771259|Clortermine
C0282152|Doxapram Hydrochloride
C0282152|Hydrochloride, Doxapram
C0282152|Stimulexin
C0282152|3,3-Diphenyl-1-ethyl-4-(2-morpholinoethyl)-2-pyrrolidinone Hydrochloride
C0282152|1-ethyl-4-[2-(4-morpholinyl)ethyl]-3,3-diphenyl-2-pyrrolidinone Monohydrochloride, Monohydrate
C0282152|respiratory stimulants doxapram hydrochloride
C0282152|doxapram hydrochloride (medication)
C0282152|Doxapram Hydrochloride [Chemical/Ingredient]
C0282152|Doxapram HCl [anesthesia] (product)
C0282152|Doxapram HCl [anesthesia]
C0282152|Doxapram hydrochloride [respiratory use] (product)
C0282152|Doxapram hydrochloride [respiratory use]
C0282152|Doxapram HCl [anaesthesia]
C0282152|Doxapram hydrochloride (substance)
C0282152|Doxapram HCl [anesthesia] (substance)
C0282152|Doxapram hydrochloride [respiratory use] (substance)
C1880248|Dapiclermin
C1880248|2-185-Ciliary neurotrophic factor (17-alanine,63-arginine) (human isoform AXOKINE)
C0058284|dimorpholamine
C0724524|Amphetamine Aspartate
C0724524|Amphetamine aspartate (substance)
C0282233|Hydrochloride, Methamphetamine
C0282233|Methamphetamine Hydrochloride
C0282233|d-N-Methyl-beta-phenylisopropylamine Hydrochloride
C0282233|Benzeneethanamine, N,alpha-dimethyl-, Hydrochloride(9CI)
C0282233|N,alpha-Dimethylphenethylamine Hydrochloride
C0282233|N-methyl-1-phenyl-propan-2-amine
C0282233|anorexics amphetamines methamphetamine hydrochloride
C0282233|methamphetamine hydrochloride (medication)
C0282233|Methamphetamine Hydrochloride [Chemical/Ingredient]
C0282233|Metamfetamine hydrochloride
C0282233|Desoxyephedrine hydrochloride
C0282233|Methamphetamine hydrochloride (product)
C0282233|Methamphetamine hydrochloride (substance)
C1880580|Etifelmine
C0011810|d Amphetamine Sulfate
C0011810|Dextroamphetamine Sulfate
C0011810|Sulfate, Dextroamphetamine
C0011810|(S)-alpha-Methylbenzeneethanamine Sulfate
C0011810|dextroamphetamine sulfate (medication)
C0011810|psychostimulants dextroamphetamine sulfate
C0011810|Dextroamphetamine Sulfate [Chemical/Ingredient]
C0011810|d-Amphetamine Sulfate
C0011810|Dextro-Amphetamine Sulfate
C0011810|d-alpha-Methylphenethylamine Sulfate
C0011810|Dextroamphetamine Sulphate
C0011810|d-Amphetamine Sulphate
C0011810|(+)-Alpha-Methylphenethylamine Sulphate (2:1)
C0011810|Benzeneethanamine, Alpha-Methyl-, (S)-, Sulfate (2:1)
C0011810|Dextro Amphetamine Sulfate
C0011810|Dexamphetamine sulfate
C0011810|Dexamphetamine sulphate
C0011810|Dexamfetamine sulphate
C0011810|Dextroamphetamine sulfate (substance)
C0546851|benzphetamine hydrochloride
C0546851|anorexics amphetamines benzphetamine hydrochloride
C0546851|benzphetamine hydrochloride (medication)
C0546851|Benzfetamine hydrochloride
C0546851|Benzphetamine hydrochloride (substance)
C0677453|cigarette
C0677453|CIGARETTES (CONTAINING TOBACCO)
C0677453|Cigarettes
C0600181|Hydrochloride, Chlorphentermine
C0600181|Chlorphentermine Hydrochloride
C0600181|chlorphentermine hydrochloride (discontinued) (medication)
C0600181|chlorphentermine hydrochloride (discontinued)
C0282051|Sulfate, Amphetamine
C0282051|Amphetamine Sulfate
C0282051|Desoxynorephedrine Sulfate
C0282051|Amphetamine Sulfate [Chemical/Ingredient]
C0282051|Amphetamine Sulfate (2:1)
C0282051|Benzeneethanamine, Alpha-Methyl-, Sulphate (2:1), (+/-)-
C0282051|(+-)-Phenisopropylamine Sulfate
C0282051|(+-)-2-Amino-1-phenylpropane Sulfate
C0282051|1-Phenyl-2-aminopropane Sulfate
C0282051|(+/-)-Alpha-Methylphenethylamine Sulfate (2:1)
C0282051|Amfetamine Sulphate
C0282051|(+-)-alpha-Methylphenethylamine Sulfate (2:1)
C0282051|(+-)-Amphetamine Sulfate
C0282051|Astedin
C0282051|dl-Amphetamine Sulfate
C0282051|dl-Amphetamine Sulphate
C0282051|amphetamine sulfate (medication)
C0282051|Amphetamine sulfate (substance)
C0282051|Amphetamine sulphate
C0700556|Hydrochloride, Phenmetrazine
C0700556|Phenmetrazine Hydrochloride
C0700556|phenmetrazine hydrochloride (discontinued) (medication)
C0700556|phenmetrazine hydrochloride (discontinued)
C0700556|Phenmetrazine Hydrochloride [Chemical/Ingredient]
C0700556|Phenmetrazine hydrochloride (product)
C0700556|Phenmetrazine hydrochloride (substance)
C0008283|Chlorphentermine
C0008283|Benzeneethanamine, 4-chloro-alpha,alpha-dimethyl-
C0008283|Chlorphentermine [Chemical/Ingredient]
C0008283|Chlorphentermine (substance)
C0700547|Maleate, Methysergide
C0700547|methysergide maleate
C0700547|Methysergide Maleate [Chemical/Ingredient]
C0700547|Methysergide maleate (substance)
C0700547|Methysergide maleate [dup] (substance)
C0952747|Dimefline Hydrochloride
C0058192|3-methyl-7-methoxy-8-dimethylamino-methylflavone
C0058192|dimefline
C0040329|Tobacco
C0040329|TABACCO
C0040329|TABACCO [VA Product]
C0040329|TOBACCO [VA Product]
C0040329|Tobacco Product
C0040329|Tobacco Products
C0040329|Product, Tobacco
C0040329|Products, Tobacco
C0040329|TOBACCO LEAF
C0040329|Tobacco (substance)
C0040329|Tobacco - substance
C0040329|Tobacco (Drug)
C0148932|phendimetrazine tartrate
C0148932|(2S,3S)-3,4-Dimethyl-2-phenylmorpholine L-(+)-tartrate(1:1)
C0148932|Morpholine, 3,4-dimethyl-2-phenyl-,(2S,3S)-,(2R,3R)-2,3-dihydroxybutanedioate(1:1)
C0148932|phendimetrazine tartrate (medication)
C0148932|anorexics phendimetrazine tartrate
C0148932|Phendimetrazine tartrate (product)
C0148932|Phendimetrazine tartrate (substance)
C0282231|Sulfate, Mephentermine
C0282231|Mephentermine Sulfate
C0282231|Mephentermine Sulfate (2:1)
C0282231|Mephentermine Sulfate [Chemical/Ingredient]
C0282231|Mephentermine sulfate (substance)
C0282231|Mephentermine sulphate
C2348683|Flubanilate Hydrochloride
C0951428|Pyrovalerone Hydrochloride
C0553808|Nondependent amphetamine or other psychostimulant abuse
C0553808|nondependent amphetamine or psychostimulant abuse
C0553808|stimulant abuse nondependent amphetamine or psychostimulant
C0553808|nondependent amphetamine or psychostimulant abuse (diagnosis)
C0553808|Nondependent amphetamine or other psychostimulant abuse (disorder)
C0553808|Nondependent amfetamine or other psychostimulant abuse
C3509117|stimulant abuse - uncomplicated (diagnosis)
C3509117|stimulant abuse - uncomplicated
C3509118|stimulant abuse with intoxication
C3509118|stimulant abuse with intoxication (diagnosis)
C3509119|stimulant abuse with intoxication - uncomplicated (diagnosis)
C3509119|stimulant abuse with intoxication - uncomplicated
C3509120|stimulant abuse with intoxication delirium (diagnosis)
C3509120|stimulant abuse with intoxication delirium
C3509121|stimulant abuse with intoxication with perceptual disturbance
C3509121|stimulant abuse with intoxication with perceptual disturbance (diagnosis)
C3509126|stimulant abuse with stimulant-induced mood disorder (diagnosis)
C3509126|stimulant abuse with stimulant-induced mood disorder
C3509127|stimulant abuse with stimulant-induced psychotic disorder
C3509127|stimulant abuse with stimulant-induced psychotic disorder (diagnosis)
C3509128|stimulant abuse with stimulant-induced psychotic disorder with delusions
C3509128|stimulant abuse with stimulant-induced psychotic disorder with delusions (diagnosis)
C3509129|stimulant abuse with stimulant-induced psychotic disorder with hallucinations
C3509129|stimulant abuse with stimulant-induced psychotic disorder with hallucinations (diagnosis)
C3509122|stimulant abuse with stimulant-induced disorder (diagnosis)
C3509122|stimulant abuse with stimulant-induced disorder
C3509123|stimulant abuse with stimulant-induced anxiety disorder
C3509123|stimulant abuse with stimulant-induced anxiety disorder (diagnosis)
C3509124|stimulant abuse with stimulant-induced sexual function (diagnosis)
C3509124|stimulant abuse with stimulant-induced sexual function
C3509125|stimulant abuse with stimulant-induced sleep disorder (diagnosis)
C3509125|stimulant abuse with stimulant-induced sleep disorder
C1456332|Stimulant abuse (disorder)
C1456332|Stimulant abuse
C1456332|stimulant abuse (diagnosis)
C1456332|Psychostimulant abuse
C1456332|abuse; stimulants
C1456332|stimulants; abuse
C3494717|Miraa abuse
C3494717|Khat abuse
C3494717|Qat abuse
C3494717|Catha edulis abuse (disorder)
C3494717|Gat abuse
C3494717|Catha edulis abuse
C3494717|stimulant abuse catja edulis
C3494717|Catha edulis abuse (diagnosis)
C2874626|Other stimulant abuse, uncomplicated
C2874631|Other stimulant abuse with intoxication
C2874631|Other stimulant abuse with intoxication, unspecified
C2874632|Other stimulant abuse with stimulant-induced mood disorder
C2874636|Other stimulant abuse with stimulant-induced psychotic disorder, unspecified
C2874636|Other stimulant abuse with stimulant-induced psychotic disorder
C2874636|Oth stimulant abuse w stim-induce psychotic disorder, unsp
C2874637|Other stimulant abuse with other stimulant-induced disorder
C2874641|Other stimulant abuse with unspecified stimulant-induced disorder
C2874641|Other stimulant abuse with unsp stimulant-induced disorder
C2874628|Other stimulant abuse with intoxication, uncomplicated
C2874629|Other stimulant abuse with intoxication delirium
C2874630|Other stimulant abuse with intoxication with perceptual disturbance
C2874630|Oth stimulant abuse w intoxication w perceptual disturbance
C3662854|Nondependent intraveous amphetamine abuse (disorder)
C3662854|Nondependent intraveous amphetamine abuse
C3662831|Nondependent amphetamine abuse (disorder)
C3662831|Nondependent amphetamine abuse
C3662831|stimulant abuse nondependent amphetamine
C3662831|Nondependent amphetamine abuse (diagnosis)
C3836657|stimulant abuse nondependent amphetamine intravenous
C3836657|nondependent intravenous amphetamine abuse (diagnosis)
C3836657|nondependent intravenous amphetamine abuse
C2874634|Other stimulant abuse with stimulant-induced psychotic disorder with delusions
C2874634|Oth stimulant abuse w stim-induce psych disorder w delusions
C2874635|Other stimulant abuse with stimulant-induced psychotic disorder with hallucinations
C2874635|Oth stimulant abuse w stim-induce psych disorder w hallucin
C2874638|Other stimulant abuse with stimulant-induced anxiety disorder
C2874638|Oth stimulant abuse with stimulant-induced anxiety disorder
C2874639|Other stimulant abuse with stimulant-induced sexual dysfunction
C2874639|Oth stimulant abuse w stimulant-induced sexual dysfunction
C2874640|Other stimulant abuse with stimulant-induced sleep disorder
C0338685|Nondependent amfetamine or psychostimulant abuse NOS
C0338685|Nondependent amphetamine or psychostimulant abuse, unspecified
C0338685|Nondependent amphetamine or psychostimulant abuse NOS
C0338685|Nondependent amfetamine or psychostimulant abuse, unspecified
C0338685|Nondependent amphetamine or psychostimulant abuse, unspecified (disorder)
C0338685|Nondependent amphetamine or psychostimulant abuse NOS (disorder)
C0338683|stimulant abuse nondependent amphetamine or psychostimulant - episodic
C0338683|nondependent amphetamine or psychostimulant abuse - episodic
C0338683|nondependent amphetamine or psychostimulant abuse - episodic (diagnosis)
C0338683|Nondependent amphetamine or psychostimulant abuse, episodic
C0338683|Nondependent amphetamine or psychostimulant abuse, episodic (life style)
C0338683|Nondependent amfetamine or psychostimulant abuse, episodic
C0338683|Nondependent amphetamine or psychostimulant abuse, episodic (disorder)
C0338683|Nondependent amphetamine or psychostimulant abuse, episodic (finding)
C0338684|Nondependent amphetamine or psychostimulant abuse in remission
C0338684|Nondependent amfetamine or psychostimulant abuse in remission
C0338684|Nondependent amphetamine or psychostimulant abuse in remission (qualifier value)
C0338684|stimulant abuse nondependent amphetamine or psychostimulant - in remission
C0338684|nondependent amphetamine or psychostimulant abuse - in remission
C0338684|nondependent amphetamine or psychostimulant abuse - in remission (diagnosis)
C0338684|Nondependent amphetamine or psychostimulant abuse in remission (life style)
C0338684|Nondependent amphetamine or psychostimulant abuse in remission (disorder)
C0338682|nondependent amphetamine or psychostimulant abuse - continuous
C0338682|nondependent amphetamine or psychostimulant abuse - continuous (diagnosis)
C0338682|stimulant abuse nondependent amphetamine or psychostimulant - continuous
C0338682|Nondependent amphetamine or psychostimulant abuse, continuous
C0338682|Nondependent amphetamine or psychostimulant abuse, continuous (life style)
C0338682|Nondependent amfetamine or psychostimulant abuse, continuous
C0338682|Nondependent amphetamine or psychostimulant abuse, continuous (disorder)
C0338682|Nondependent amphetamine or psychostimulant abuse, continuous (finding)
C2104574|continuous methamphetamine abuse
C2104574|continuous methamphetamine abuse (diagnosis)
C2104575|episodic methamphetamine abuse (diagnosis)
C2104575|episodic methamphetamine abuse
C2104576|methamphetamine abuse in remission (diagnosis)
C2104576|methamphetamine abuse in remission
