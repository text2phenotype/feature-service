C0010054|Coronary Arteriosclerosis
C1956346|Coronary Artery Disease
C0010054|Arterioscleroses, Coronary
C0010054|Coronary Arterioscleroses
C0010054|Coronary Arteriosclerosis
C0010054|Coronary atherosclerosis
C0010054|Atherosclerotic heart disease
C0010054|coronary arteriosclerosis (diagnosis)
C0010054|ASHD - Atherosclerotic heart disease
C0010054|Atherosclerosis of coronary artery
C0010054|Atherosclerosis of coronary artery (disorder)
C0010054|Cardiac sclerosis
C0010054|Coronary (artery) atherosclerosis
C0010054|Coronary (artery) sclerosis
C0010054|Disease;atherosclerotic;heart
C0010054|Atherosclerotic heart disease NOS
C0010054|Atherosclerosis, Coronary
C0010054|Arteriosclerosis, Coronary
C0010054|atherosclerosis of coronary artery (diagnosis)
C0010054|atherosclerosis coronary artery
C0010054|Coronary atherosclerosis (disorder)
C0010054|Coronary sclerosis
C0010054|Arteriosclerotic heart disease
C0010054|ASHD
C0010054|Coronary artherosclerosis
C0010054|Coronary artery sclerosis
C0010054|Coronary artery atherosclerosis
C0010054|Arteriosclerosis coronary artery
C0010054|cardiac; sclerosis
C0010054|coronary; arteriosclerosis
C0010054|coronary; sclerosis
C0010054|disease (or disorder); arteriosclerotic, coronary (artery)
C0010054|disease (or disorder); arteriosclerotic, heart
C0010054|heart; arteriosclerosis
C0010054|sclerosis; cardiac
C0010054|sclerosis; coronary
C0010054|arteriosclerosis; coronary (artery)
C0010054|arteriosclerosis; coronary
C0010054|arteriosclerosis; heart
C0010054|Atheroscleroses, Coronary
C0010054|Coronary Atheroscleroses
C0010054|Coronary arteriosclerosis (disorder)
C0010054|Coronary artery arteriosclerosis
C0002963|Prinzmetal angina
C0002963|Angina Pectoris, Variant
C0002963|Prinzmetals Angina
C0002963|Variant Angina Pectoris
C0002963|Angina, Prinzmetal's
C0002963|Prinzmetal's angina
C0002963|Variant Angina
C0002963|Prinzmental angina
C0002963|Prinzmetal's angina (diagnosis)
C0002963|Angina Pectoris, Variant [Disease/Finding]
C0002963|Angina, Prinzmetal
C0002963|Vasospastic angina
C0002963|Coronary artery spasm angina
C0002963|Prinzmetal angina (disorder)
C0002963|Prinzmetal; angina
C0002963|angina pectoris; variant
C0002963|variant; angina
C0596384|coronary fibrosis
C0178570|coronary occlusion/thrombosis
C0542269|Non-Q wave myocardial infarction NOS
C0542269|Non-Q wave myocardial infarction
C0542269|acute non-Q-wave myocardial infarction
C0542269|acute non-Q-wave myocardial infarction (diagnosis)
C0542269|subendocardial non-Q-wave myocardial infarction acute
C0542269|Non-Q wave myocardial infarction (disorder)
C0542060|Ischemia coronary artery origin
C0542060|Ischaemia coronary artery origin
C0542060|ischemia; coronary
C0856737|Single vessel disease
C0856738|Triple vessel disease
C0856739|Left main stem disease
C0856740|Main stem disease
C0857530|Right main stem disease
C0375265|Cor ath bypass graft NOS
C0375265|Coronary atherosclerosis of unspecified bypass graft
C0375265|Coronary atherosclerosis of unspecified type of bypass graft
C0375265|Coronary atherosclerosis of bypass graft
C0375265|Coronary atherosclerosis of bypass graft NOS
C0340285|3-vessel coronary artery stenosis (diagnosis)
C0340285|3-vessel coronary artery stenosis
C0340285|Triple vessel coronary artery disease (disorder)
C0340285|Triple vessel coronary artery disease
C0340285|Triple vessel disease of the heart
C0340285|arteriosclerosis coronary artery triple vessel disease
C0340285|triple vessel disease of heart
C0340285|triple vessel disease of heart (diagnosis)
C0340285|Triple vessel disease of the heart (disorder)
C2366973|coronary arteriosclerosis due to lipid-rich plaque
C2366973|coronary arteriosclerosis due to lipid-rich plaque (diagnosis)
C2062869|asymptomatic coronary arteriosclerosis (diagnosis)
C2062869|asymptomatic coronary arteriosclerosis
C0685094|calcific coronary arteriosclerosis
C0685094|calcific coronary arteriosclerosis (diagnosis)
C0685094|coronary arteriosclerosis due to calcified coronary lesion
C0685094|coronary arteriosclerosis due to calcified coronary lesion (diagnosis)
C0685094|Calcific coronary arteriosclerosis (disorder)
C2321373|progressive coronary artery disease
C2321373|progressive coronary artery disease (diagnosis)
C2321817|sample template coronary artery disease
C2321817|sample template coronary artery disease (diagnosis)
C1997154|Coronary arteriosclerosis due to radiation
C1997154|coronary arteriosclerosis due to radiation (diagnosis)
C1997154|Coronary arteriosclerosis caused by radiation
C1997154|Coronary arteriosclerosis caused by radiation (disorder)
C1997154|Coronary arteriosclerosis due to radiation (disorder)
C3472163|Coronary arteriosclerosis in native artery (disorder)
C3472163|Coronary arteriosclerosis in native artery
C3472163|arteriosclerosis coronary in native artery
C3472163|Coronary arteriosclerosis in native artery (diagnosis)
C1956346|CAD
C1956346|Coronary artery disease
C1956346|Artery Diseases, Coronary
C1956346|Coronary Artery Diseases
C1956346|Disease, Coronary Artery
C1956346|Artery Disease, Coronary
C1956346|Diseases, Coronary Artery
C1956346|CORONARY ARTERY DIS
C1956346|CAD (coronary artery disease)
C1956346|disorder of coronary arteries (diagnosis)
C1956346|coronary artery disease (diagnosis)
C1956346|disorder of coronary arteries
C1956346|Coronary artery disorders
C1956346|Coronary Disease
C1956346|Coronary Artery Disease [Disease/Finding]
C1956346|Coronary artery disease (disorder)
C1956346|Disease of the coronary arteries
C1956346|CAD - Coronary artery disease
C1956346|coronary heart disease
C1956346|Coronary artery disorder
C1956346|Disease coronary artery
C1956346|Disorder coronary artery
C1956346|Coronary artery disorder (NOS)
C1956346|Coronary artery disease NOS
C1956346|Cardio/pulm: Coronary artery disease
C1956346|coronary (artery); disease
C1956346|disease (or disorder); artery, coronary
C1956346|disease (or disorder); coronary (artery)
C1956346|disease (or disorder); heart, artery, arterial
C1956346|artery; disorder, coronary
C1956346|Coronary artery disease, NOS
C1956346|Disorder of coronary artery (disorder)
C1956346|Disorder of coronary artery
C0948089|Acute Coronary Syndrome
C0948089|Coronary Syndromes, Acute
C0948089|Syndromes, Acute Coronary
C0948089|Acute Coronary Syndromes
C0948089|Syndrome, Acute Coronary
C0948089|Coronary Syndrome, Acute
C0948089|Acute Coronary Syndrome [Disease/Finding]
C0948089|Acute coronary syndrome (disorder)
C0948089|acute coronary syndrome (diagnosis)
C0948089|ACS - Acute coronary syndrome
C0340325|Coronary thrombosis not resulting in myocardial infarction
C0340325|Aborted myocardial infarction
C0340325|MI - Myocardial infarction aborted
C0340325|Aborted myocardial infarction (disorder)
C0340325|Coronary thrombosis not leading to myocardial infarction
C0340325|Coronary thrombosis not resulting in myocardial infarction (disorder)
C0340325|coronary; thrombosis, not resulting in infarction
C0340325|thromboembolism; coronary, not resulting in infarction
C0340325|thrombosis; cardiac, not resulting in infarction
C0340325|thrombosis; coronary, not resulting in infarction
C0002962|Angina Pectoris
C0002962|Stenocardias
C0002962|Angina
C0002962|Angina pectoris, unspecified
C0002962|stenocardia
C0002962|angina pectoris (diagnosis)
C0002962|Anginal syndrome
C0002962|Cardiac angina
C0002962|Angina of effort
C0002962|Ischemic chest pain
C0002962|Angina NOS
C0002962|Angina Pectoris [Disease/Finding]
C0002962|Angor Pectoris
C0002962|Pain;angina
C0002962|Angina pectoris (disorder)
C0002962|Angina (disorder)
C0002962|Angina pectoris NOS
C0002962|Stenocardia (disorder)
C0002962|Angina pectoris NOS (disorder)
C0002962|Ischaemic chest pain
C0002962|Ischaemic chest pain (disorder)
C0002962|Chest pain - cardiac
C0002962|chest pain ischemic
C0002962|Ischemic chest pain (diagnosis)
C0002962|Anginal discomfort
C0002962|Angina syndrome
C0002962|Anginal pain
C0002962|Cardio/pulm: Angina
C0002962|Ischaemic heart disease - angina
C0002962|Ischemic heart disease - angina
C0002962|AP - Angina pectoris
C0002962|Ischemic chest pain (finding)
C0002962|chest; pain, ischemic
C0002962|pain; chest, ischemic
C0002962|syndrome; anginal
C0002962|anginal; syndrome
C0002962|Angina pectoris, NOS
C0002962|Angina, NOS
C0002962|Angina pectoris (disorder) [Ambiguous]
C0002962|Angina, cardiac
C0002962|angina pain
C0264692|Ischemic contracture of left ventricle syndrome
C0264692|Stone heart syndrome
C0264692|Ischaemic contracture of left ventricle syndrome
C0264692|Ischemic contracture of left ventricle syndrome (disorder)
C1510446|Acute ischaemic heart disease, unspecified
C1510446|Acute ischemic heart disease, unspecified
C1510446|acute ischemic heart disease (diagnosis)
C1510446|Acute ischemic heart disease
C1510446|Acute ischemic heart disease (disorder)
C1510446|Acute ischaemic heart disease
C0264684|Arteritis coronary
C0264684|Coronary arteritis
C0264684|Coronary endarteritis
C0264684|Coronary arteritis (disorder)
C0264684|coronary; arteritis
C0264684|arteritis; coronary
C0264684|Coronary artery arteritis or endarteritis
C0264684|Coronary arteritis or endarteritis
C0152107|Dressler's syndrome
C0152107|Postmyocardial infarction syndrome
C0152107|Dressler's syndrome (diagnosis)
C0152107|Post MI syndrome
C0152107|Dresslers syndrome
C0152107|Post myocardial infarction syndrome
C0152107|Postmyocardial infarction pericarditis
C0152107|Post-myocardial infarction syndrome
C0152107|Postmyocardial infarction syndrome (disorder)
C0152107|postmyocardial infarction; syndrome
C0152107|syndrome; postmyocardial infarction
C0152107|Dressler
C0152107|Postmyocardial infarct syndrom
C1279369|Asymptomatic coronary heart disease (disorder)
C1279369|Asymptomatic coronary heart disease
C0264695|Subendocardial ischaemia
C0264695|subendocardial ischemia (diagnosis)
C0264695|subendocardial ischemia
C0264695|Subendocardial ischemia (disorder)
C0264695|ischemia; subendocardial
C0264687|coronary strictire
C0264687|coronary strictire (diagnosis)
C0264687|Coronary stricture
C0264687|Coronary stricture (disorder)
C0264687|coronary; stricture
C0264687|stricture; coronary artery
C0264687|stricture; coronary
C0264687|Coronary artery stricture
C0151744|Disease, Ischemic Heart
C0151744|Diseases, Ischemic Heart
C0151744|Heart Diseases, Ischemic
C0151744|Ischemic Heart Diseases
C0151744|Myocardial Ischemia
C0151744|Ischemias, Myocardial
C0151744|Myocardial Ischemias
C0151744|Ischaemic heart diseases
C0151744|Myocardial ischaemia
C0151744|Ischemic Heart Disease
C0151744|IHD
C0151744|HEART DIS ISCHEMIC
C0151744|ISCHEMIC HEART DIS
C0151744|myocardial ischemia (diagnosis)
C0151744|Heart Disease, Ischemic
C0151744|Ischemia, Myocardial
C0151744|Myocardial Ischemia [Disease/Finding]
C0151744|Disease;ischaemic heart
C0151744|myocardial ischemia/hypoxia
C0151744|Ischemic heart diseases (I20-I25)
C0151744|Ischaemic heart disease (disorder)
C0151744|Cardiac ischaemia
C0151744|Ischaemic heart disease
C0151744|Ischaemic heart disease NOS
C0151744|Ischemic heart disease NOS
C0151744|IHD - Ischemic heart disease
C0151744|Ischemic heart disease NOS (disorder)
C0151744|Myocardial ischaemia (disorder)
C0151744|IHD - Ischaemic heart disease
C0151744|Ischemic heart disease (disorder)
C0151744|Cardiac ischemia
C0151744|Ischaemic heart disease NOS (disorder)
C0151744|ischemic heart disease (diagnosis)
C0151744|Ischaemia myocardial
C0151744|Ischemia myocardial
C0151744|ischemia; heart
C0151744|ischemia; myocardial
C0151744|myocardium; ischemic
C0151744|Ischemic heart disease, NOS
C0151744|Ischaemic heart disease, NOS
C0151744|Myocardial ischemia, NOS
C0151744|Myocardial ischemia (disorder)
C0151744|Disease;ischemic heart
C0340287|Other specified ischaemic heart disease
C0340287|Other specified ischemic heart disease
C0340287|Other specified ischemic heart disease (disorder)
C0349466|myocardial ischemia of newborn
C0349466|myocardial ischemia of newborn (diagnosis)
C0349466|Myocardial ischaemia of newborn
C0349466|Myocardial ischemia of newborn (disorder)
C0340283|Other acute and subacute forms of ischemic heart disease
C0340283|Other acute and subacute forms of ischaemic heart disease
C0340283|Ac ischemic hrt dis NEC
C0340283|Other acute and subacute forms of ischemic heart disease, other
C0340283|Other acute and subacute ischemic heart disease
C0340283|Other acute and subacute ischaemic heart disease
C0340283|Other acute and subacute ischaemic heart disease NOS
C0340283|Other acute and subacute ischemic heart disease (disorder)
C0340283|Other acute and subacute ischaemic heart disease (disorder)
C0340283|Other acute and subacute ischemic heart disease NOS
C0340283|Other acute and subacute ischemic heart disease NOS (disorder)
C1533195|Chronic coronary insufficiency
C0018789|Aneurysms, Cardiac
C0018789|Aneurysms, Heart
C0018789|Cardiac Aneurysms
C0018789|Heart Aneurysm
C0018789|Heart Aneurysms
C0018789|Aneurysm of heart
C0018789|Aneurysm, Cardiac
C0018789|Aneurysm, Heart
C0018789|Cardiac aneurysm
C0018789|Heart Aneurysm [Disease/Finding]
C0018789|Aneurysm;cardiac
C0018789|Aneurysm of heart NOS
C0018789|Aneurysm of heart (disorder)
C0018789|Aneurysm of heart NOS (disorder)
C0018789|cardiac; aneurysm
C0018789|heart; aneurysm
C0018789|aneurysm; cardiac
C0018789|aneurysm; heart
C0018789|Aneurysm of heart, NOS
C0010072|Coronary Thromboses
C0010072|Coronary Thrombosis
C0010072|Thromboses, Coronary
C0010072|Coronary artery thrombosis
C0010072|coronary artery thrombosis (diagnosis)
C0010072|coronary (artery) thrombosis
C0010072|Coronary Thrombosis [Disease/Finding]
C0010072|Thrombosis, Coronary
C0010072|Thrombosis;artery;coronary
C0010072|Coronary artery thrombosis (disorder)
C0010072|CT - Coronary thrombosis
C0010072|Thrombosis - coronary
C0010072|Thrombosis coronary
C0264683|Coronary (artery) atheroma
C0264683|Coronary atheroma
C0264683|coronary artery atheroma (diagnosis)
C0264683|Coronary artery atheroma
C0264683|Atheroma coronary artery
C0264683|Coronary artery atheroma (disorder)
C0264683|atheroma; coronary
C0264683|atheroma; heart
C0264683|coronary; atheroma
C0264683|heart; atheroma
C0155669|Other forms of chronic ischemic heart disease
C0155669|Other forms of chronic ischaemic heart disease
C0155669|Other forms of chronic ischemic heart disease, other
C0155669|Other forms of chronic ischaemic heart disease, other
C0155669|[X]Other forms of chronic ischaemic heart disease
C0155669|[X]Other forms of chronic ischemic heart disease (disorder)
C0155669|Other chronic ischaemic heart disease
C0155669|[X]Other forms of chronic ischemic heart disease
C0155669|Other chronic ischaemic heart disease NOS
C0155669|Other chronic ischemic heart disease NOS
C0155669|Other chronic ischemic heart disease
C0155669|Other chronic ischemic heart disease (disorder)
C0155669|Other chronic ischemic heart disease NOS (disorder)
C0348589|Other current complications following acute myocardial infarction
C0348589|Oth current complications following AMI
C0348589|[X]Other current complications following acute myocardial infarction (disorder)
C0348589|[X]Other current complications following acute myocardial infarction
C0009693|Congenital coronary artery sclerosis
C0009693|Congenital coronary artery sclerosis (disorder)
C0340291|Silent myocardial ischaemia
C0340291|Silent myocardial ischemia
C0340291|silent myocardial ischemia (diagnosis)
C0340291|Silent myocardial ischaemia (disorder)
C0340291|Silent myocardial ischemia (disorder)
C0340291|Asymptomatic ischaemia
C0340291|Asymptomatic ischemia
C0340291|ischemia; myocardial, subclinical
C0581375|2-vessel coronary artery stenosis (diagnosis)
C0581375|2-vessel coronary artery stenosis
C0581375|Two Vessel Coronary Disease
C0581375|Double vessel coronary artery disease
C0581375|Double vessel coronary artery disease (disorder)
C0581375|TWO VESSEL DISEASE
C0581375|Double coronary vessel disease
C0581375|Two coronary vessel disease
C0581375|Double coronary vessel disease (disorder)
C0581374|single vessel coronary artery stenosis
C0581374|single vessel coronary artery stenosis (diagnosis)
C0581374|Single vessel coronary artery disease (disorder)
C0581374|Single vessel coronary artery disease
C0581374|Single coronary vessel disease
C0581374|Single coronary vessel disease (disorder)
C0264696|Microinfarction of heart
C0264696|Microinfarction of heart (disorder)
C0264696|microinfarct of heart (diagnosis)
C0264696|Microinfarct of heart
C0264696|Microinfarct of heart (disorder)
C0264696|microinfarct; heart
C0349780|ischemic myocardial dysfunction (diagnosis)
C0349780|Ischemic myocardial dysfunction
C0349780|Ischaemic myocardial dysfunction
C0349780|Ischemic myocardial dysfunction (disorder)
C0264694|Chronic ischemic heart disease
C0264694|Chronic ischemic heart disease, unspecified
C0264694|Chronic ischaemic heart disease
C0264694|Chronic ischaemic heart disease, unspecified
C0264694|chronic myocardial ischemia
C0264694|chronic myocardial ischemia (diagnosis)
C0264694|Chr ischemic hrt dis NOS
C0264694|Ischemic heart disease (chronic) NOS
C0264694|Ischaemia;myocardial;chronic
C0264694|chronic ischemic heart disease (diagnosis)
C0264694|Chr. ischemic heart dis. NOS
C0264694|Chronic ischaemic heart disease NOS
C0264694|Chronic ischemic heart disease NOS
C0264694|Chronic ischemic heart disease (disorder)
C0264694|Chronic ischemic heart disease NOS (disorder)
C0264694|Chronic myocardial ischaemia
C0264694|Chr. ischaemic heart dis. NOS
C0264694|Chronic myocardial ischaemia (disorder)
C0264694|Chronic ischaemic heart disease NOS (disorder)
C0264694|Chronic myocardial ischemia (disorder)
C0264694|Disease;ischaem heart;chronic
C0264694|Ischemia;myocardial;chronic
C3650149|atherosclerosis of other coronary vessels (diagnosis)
C3650149|atherosclerosis of other coronary vessels
C3650188|atherosclerosis of coronary artery with unstable angina pectoris (diagnosis)
C3650188|atherosclerosis coronary artery with unstable angina pectoris
C3650188|atherosclerosis of coronary artery with unstable angina pectoris
C3650187|atherosclerosis of coronary artery without angina pectoris
C3650187|atherosclerosis of coronary artery without angina pectoris (diagnosis)
C3650187|atherosclerosis coronary artery without angina pectoris
C2882208|Atherosclerosis of other coronary vessels without angina pectoris
C2882208|atherosclerosis of other coronary vessels without angina pectoris (diagnosis)
C3650190|atherosclerosis of coronary artery with angina pectoris
C3650190|atherosclerosis of coronary artery with angina pectoris (diagnosis)
C3650190|atherosclerosis coronary artery with angina pectoris
C3650189|atherosclerosis of coronary artery with angina pectoris with documented spasm
C3650189|atherosclerosis of coronary artery with angina pectoris with documented spasm (diagnosis)
C3650189|atherosclerosis coronary artery with angina pectoris with documented spasm
C2349509|Coronary atherosclerosis due to lipid rich plaque
C2349509|Cor ath d/t lpd rch plaq
C2349509|coronary atherosclerosis due to lipid-rich plaque
C2349509|coronary atherosclerosis due to lipid-rich plaque (diagnosis)
C3161090|Cor ath d/t calc cor lsn
C3161090|Coronary atherosclerosis due to calcified coronary lesion
C3161090|atherosclerosis due calcified coronary lesion
C3161090|coronary atherosclerosis due calcified coronary lesion
C3161090|coronary atherosclerosis due to calcified coronary lesion (diagnosis)
C1867743|Coronary artery disease, premature
C1867743|premature coronary heart disease
C1867743|coronary artery disease premature
C1867743|premature coronary heart disease (diagnosis)
C1867743|Premature coronary artery disease
C1997109|Coronary arteriosclerosis of coronary artery bypass graft
C1997109|Arteriosclerosis in coronary artery bypass graft
C1997109|Arteriosclerosis in coronary artery bypass graft (disorder)
C1997109|Arteriosclerosis of coronary artery bypass graft (disorder)
C1997109|Arteriosclerosis of coronary artery bypass graft
C1997109|arteriosclerosis of coronary artery bypass graft (diagnosis)
C1996973|Recurrent coronary arteriosclerosis after percutaneous transluminal coronary angioplasty (disorder)
C1996973|Recurrent coronary arteriosclerosis after percutaneous transluminal coronary angioplasty
C1996973|Recurrent coronary arteriosclerosis after percutaneous transluminal coronary angioplasty (diagnosis)
C1996973|coronary arteriosclerosis recurrent after percutaneous transluminal angioplasty
C1842247|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT, 1
C1842247|ADCAD1
C1842247|Coronary Artery Disease With Myocardial Infarction
C1842247|CAD autosomal dominant 1 (diagnosis)
C1842247|coronary artery disease autosomal dominant 1
C1842247|CAD autosomal dominant 1
C1842247|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT 1
C1842247|CORONARY ARTERY DISEASE/MYOCARDIAL INFARCTION
C1970440|ADCAD2
C1970440|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT 2
C1970440|CORONARY ARTERY DISEASE, AUTOSOMAL DOMINANT 2 (disorder)
C1970440|CAD autosomal dominant 2 (diagnosis)
C1970440|CAD autosomal dominant 2
C1970440|coronary artery disease autosomal dominant 2
C4039929|Coronary arteriosclerosis after percutaneous coronary angioplasty
C4039929|Coronary arteriosclerosis after percutaneous coronary angioplasty (disorder)
C4074915|Coronary arteriosclerosis following coronary artery bypass graft (disorder)
C4074915|Coronary arteriosclerosis following coronary artery bypass graft
C0340326|Accelerated coronary artery disease in transplanted heart (diagnosis)
C0340326|coronary artery disease in transplanted heart accelerated
C0340326|Accelerated coronary artery disease in transplanted heart
C0340326|Accelerated coronary artery disease in transplanted heart (disorder)
C1299432|Multi vessel coronary artery disease
C1299432|multi vessel coronary artery disease (diagnosis)
C1299432|Multi vessel coronary artery disease (disorder)
C1299433|Left main coronary artery disease (diagnosis)
C1299433|Left main coronary artery disease
C1299433|coronary artery disease left main
C1299433|Left main coronary artery disease (disorder)
C1299434|coronary artery disease of significant bypass graft
C1299434|Significant coronary bypass graft disease (diagnosis)
C1299434|Significant coronary bypass graft disease
C1299434|Significant coronary bypass graft disease (disorder)
C1384784|a.coronaria; obstruction
C1384784|obstruction; coronary artery
C1384785|a.coronaria; stricture, coronary
C0242231|Coronary Stenosis
C0242231|Stenoses, Coronary
C0242231|Stenosis, Coronary
C0242231|Coronary artery stenosis
C0242231|coronary artery stenosis (diagnosis)
C0242231|Coronary Stenosis [Disease/Finding]
C0242231|Coronary Stenoses
C0242231|Artery Stenoses, Coronary
C0242231|Artery Stenosis, Coronary
C0242231|Coronary Artery Stenoses
C0242231|Stenoses, Coronary Artery
C0242231|Stenosis, Coronary Artery
C0242231|Narrow coronary arteries
C0242231|Coronary arteries--Stenosis
C0242231|Coronary artery stenosis (disorder)
C0242231|coronary; stenosis
C0242231|a.coronaria; narrowing
C0242231|narrowing; coronary artery
C0242231|stenosis; artery, coronary
C0242231|stenosis; coronary
C0242231|artery; stenosis, coronary
C1384962|disease (or disorder); heart, arteriosclerotic or sclerotic (senile)
C1388510|cardiac; arteriosclerosis
C1388510|arteriosclerosis; cardiac
C1388511|arteriosclerosis; cardiomyopathy
C1388512|arteriosclerosis; cardiopathy
C1404464|atheroma; myocardial
C1404464|myocardium; atheroma
C1391994|cardiomyopathy; arteriosclerotic
C1392010|cardiopathy; arteriosclerotic
C1392034|cardiosclerosis
C1394006|coronary; obstruction
C1394006|obstruction; coronary
C1399178|cardiac; ossification
C1399178|coronary; ossification
C1399178|heart; ossification
C1399178|ossification; cardiac
C1399178|ossification; coronary
C1399178|ossification; heart
C1394968|degeneration; heart, atheromatous
C1394968|heart; degeneration, atheromatous
C1399129|heart; disease, artery, arterial
C1399130|heart; disease, arteriosclerotic or sclerotic (senile)
C1328505|Myocardial sclerosis
C1328505|myocardium; sclerosis
C1328505|sclerosis; myocardial
C1636672|coronary artery disease obliterative
C1636672|Obliterative coronary artery disease (diagnosis)
C1636672|Obliterative coronary artery disease
C1636672|Obliterative coronary artery disease (disorder)
C0837136|Crn ath nonatlg blg grft
C0837136|Atherosclerotic heart disease, of nonautologous bypass graft
C0837136|Coronary atherosclerosis of nonautologous biological bypass graft
C0837134|Crnry athrscl natve vssl
C0837134|Atherosclerotic heart disease of native coronary artery
C0837134|Coronary atherosclerosis of native coronary artery
C0837133|Cor ath unsp vsl ntv/gft
C0837133|Coronary atherosclerosis of unspecified type of vessel, native or graft
C0837135|Crn ath atlg vn bps grft
C0837135|Coronary atherosclerosis of autologous vein bypass graft
C0837135|Coronary atherosclerosis of autologous biological bypass graft
C1456095|Cor ath bps graft tp hrt
C1456095|Coronary atherosclerosis of bypass graft (artery) (vein) of transplanted heart
C0375264|Cor ath artry bypas grft
C0375264|Atherosclerosis of coronary artery bypass graft NOS
C0375264|atherosclerosis of coronary artery bypass graft (diagnosis)
C0375264|atherosclerosis of coronary artery bypass graft
C0375264|atherosclerosis coronary artery bypass graft
C0375264|Coronary atherosclerosis of artery bypass graft
C1135190|Cor ath natv art tp hrt
C1135190|Coronary atherosclerosis of native coronary artery of transplanted heart
C0852153|Coronary artery disorders NEC
C0852149|Ischaemic coronary artery disorders
C0852149|Ischemic coronary artery disorders
C2584623|Furcation lesion of coronary artery
C2584623|Furcation lesion of coronary artery (disorder)
C2711976|Fracture of stent of coronary artery (disorder)
C2711976|Fracture of stent of coronary artery
C1611184|Coronary artery calcification
C1611184|Calcification of coronary artery (disorder)
C1611184|Calcification of coronary artery
C2062867|rebound angina due to beta blocker withdrawal
C2062867|beta-blocker withdrawal (rebound angina)
C2062867|rebound angina due to beta blocker withdrawal (diagnosis)
C0003851|Arteriosclerosis Obliterans
C0003851|Obliterans, Arteriosclerosis
C0003851|arteriosclerosis obliterans (diagnosis)
C0003851|Arteriosclerosis Obliterans [Disease/Finding]
C0003851|Arteriosclerosis obliterans (disorder)
C0003851|Arteriosclerosis obliterans (disorder) [Ambiguous]
C0264686|Coronary artery embolism
C0264686|coronary artery embolism (diagnosis)
C0264686|coronary (artery) embolism
C0264686|Embolism;artery;coronary
C0264686|Coronary embolism
C0264686|Embolus coronary artery
C0264686|Coronary embolus
C0264686|Coronary artery embolism (disorder)
C2049072|induced CPK elevation
C2049072|induced CPK elevation (diagnosis)
C0008031|Chest Pain
C0008031|Chest Pains
C0008031|Pain, Chest
C0008031|Pains, Chest
C0008031|Chest pain, unspecified
C0008031|[D]Chest pain (context-dependent category)
C0008031|[D]Chest pain NOS (context-dependent category)
C0008031|[D]Chest pain, unspecified (context-dependent category)
C0008031|Thoracic pain
C0008031|chest pain or discomfort (symptom)
C0008031|chest pain or discomfort
C0008031|chest pain (diagnosis)
C0008031|Pain in chest
C0008031|Chest pain NOS
C0008031|Nonspecific chest pain
C0008031|Chest Pain [Disease/Finding]
C0008031|Pain;chest
C0008031|Chest pain (finding)
C0008031|[D]Chest pain NOS
C0008031|[D]Chest pain (situation)
C0008031|[D]Chest pain
C0008031|[D]Chest pain, unspecified (situation)
C0008031|[D]Chest pain, unspecified
C0008031|Chest pain NOS (finding)
C0008031|[D]Chest pain NOS (situation)
C0008031|Thorax painful
C0008031|chest pain or discomfort reported as pain
C0008031|chest pain or discomfort reported as pain (symptom)
C0008031|reported chest pain
C0008031|thoracodynia
C0008031|thoracalgia
C0008031|Unspecified chest pain
C0008031|Thorax pain
C0008031|Pain chest
C0008031|chest; pain
C0008031|pain; chest
C0008031|pain; thorax
C0008031|thorax; pain
C0008031|Chest pain, NOS
C2024793|cardiac wall motion dysfunction (diagnosis)
C2024793|cardiac wall motion dysfunction
C0010073|Artery Vasospasm, Coronary
C0010073|Artery Vasospasms, Coronary
C0010073|Coronary Artery Vasospasms
C0010073|Coronary Vasospasm
C0010073|Coronary Vasospasms
C0010073|Vasospasm, Coronary
C0010073|Vasospasm, Coronary Artery
C0010073|Vasospasms, Coronary
C0010073|Vasospasms, Coronary Artery
C0010073|coronary artery spasm
C0010073|coronary artery spasm (diagnosis)
C0010073|Arteriospasm coronary
C0010073|Coronary Vasospasm [Disease/Finding]
C0010073|Coronary Artery Vasospasm
C0010073|Spasm;artery;coronary
C0010073|Coronary spasm
C0010073|Coronary vascular spasm
C0010073|Spasm coronary artery
C0010073|Coronary artery spasm (disorder)
C0010073|coronary; spasm
C0010073|a.coronaria; spasm
C0010073|spasm; coronary artery
C0010073|spasm; coronary
C0428837|coronary collateral circulation (diagnosis)
C0428837|coronary collateral circulation
C0428837|Coronary artery collaterals
C0428837|Coronary artery collaterals (finding)
C2063730|coronary ectasia
C2063730|coronary ectasia (diagnosis)
C2063731|coronary ostial membrane
C2063731|coronary ostial membrane (diagnosis)
C0428830|coronary bypass graft stenosis (diagnosis)
C0428830|coronary bypass graft stenosis
C0428830|Coronary graft stenosis
C0428830|coronary graft; stenosis
C0428830|stenosis; coronary graft
C0428830|Coronary graft stenosis (disorder)
C0428830|Coronary graft stenosis (finding)
C0349781|hibernating myocardium (diagnosis)
C0349781|hibernating myocardium
C0349781|Hibernating myocardium (disorder)
C1299451|post-angioplasty coronary
C1299451|post coronary angioplasty (diagnosis)
C1299451|post coronary angioplasty
C1299451|post-angioplasty
C1299451|Patient post angioplasty (finding)
C1299451|Patient post angioplasty
C3665365|ASCVD (arteriosclerotic cardiovascular disease)
C3665365|arteriosclerotic CV disease
C3665365|Cardiovascular degeneration with arteriosclerosis
C3665365|Cardiovascular sclerosis with arteriosclerosis
C3665365|Cardiovascular arteriosclerosis unspecified
C3665365|ASCVD
C3665365|Cardiovascular arteriosclerosis
C3665365|Cardiovascular disease with arteriosclerosis
C3665365|Cardiovascular arteriosclerosis unspecified (disorder)
C3665365|Arteriosclerotic cardiovascular disease (disorder)
C3665365|Arteriosclerotic cardiovascular disease
C3665365|arteriosclerotic cardiovascular disease (ASCVD)
C3665365|arteriosclerotic cardiovascular disease (ASCVD) (diagnosis)
C3665365|Arteriosclerotic cardiovascular disease, NOS
C3665365|cardiovascular; arteriosclerosis
C3665365|disease (or disorder); arteriosclerotic, cardiovascular
C3665365|arteriosclerosis; cardiovascular
C2957458|native coronary artery stenosis
C2957458|native coronary artery stenosis (diagnosis)
C0340664|Coronary artery perforation
C0340664|Coronary artery perforation (disorder)
C0345134|Variant dominance of coronary circulation
C0345134|Variant dominance of coronary circulation (disorder)
C0347699|Transection of coronary artery
C0347699|Transection of coronary artery (disorder)
C0158623|congenital anomaly of coronary artery (diagnosis)
C0158623|congenital anomaly of coronary artery
C0158623|Coronary artery anomaly
C0158623|Coronary artery anomaly, congenital
C0158623|Coronary artery anomaly NOS
C0158623|Coronary artery abnormality (disorder)
C0158623|Coronary artery abnormality
C0158623|Coronary artery anomaly NOS (disorder)
C0158623|Coronary arteries--Abnormalities
C0158623|Abnormality of the coronary arteries
C0158623|Congenital coronary artery malformation NOS
C0158623|Congenital coronary artery malformation
C0158623|Congenital anomaly of coronary artery (disorder)
C0158623|coronary artery; anomaly
C0158623|coronary; artery, anomaly
C0158623|deformity; artery, coronary, congenital
C0158623|a.coronaria; anomaly
C0158623|anomaly; coronary artery
C0158623|artery; deformity, coronary, congenital
C0158623|Congenital anomaly of coronary artery, NOS
C0158623|Coronary artery abnormality [Ambiguous]
C0392158|Dissecting aneurysm of coronary artery
C0392158|Dissecting coronary artery aneurysm
C0392158|Coronary artery aneurysm and dissection
C0392158|Aneurysm dissecting coronary artery
C0392158|Dissecting aneurysm of coronary artery (disorder)
C0010051|Aneurysms, Coronary
C0010051|Coronary Aneurysm
C0010051|Coronary Aneurysms
C0010051|Coronary artery aneurysm
C0010051|aneurysm of coronary artery (diagnosis)
C0010051|aneurysm of coronary artery
C0010051|Aneurysm coronary vessel
C0010051|Coronary Aneurysm [Disease/Finding]
C0010051|Aneurysm, Coronary
C0010051|Aneurysm;artery;coronary
C0010051|Aneurysmal lesion of coronary artery
C0010051|Aneurysmal lesion of coronary artery (finding)
C0010051|Aneurysm of coronary vessels
C0010051|Aneurysm of coronary vessels (disorder)
C0010051|coronary; aneurysm
C0010051|aneurysm; coronary
C0010051|Arteriovenous aneurysm of coronary vessels
C0265899|Congenital absence of coronary artery (disorder)
C0265899|Congenital absence of coronary artery
C0265899|absence; artery, coronary
C0265899|artery; absence, coronary
C0265899|Coronary artery, absence
C0340648|Coronary artery dissection
C0340648|dissection of coronary artery
C0340648|dissection of coronary artery (diagnosis)
C0340648|Dissection cor artery
C0340648|Coronary artery dissection (disorder)
C0343692|Syphilitic coronary artery disease
C0343692|syphilis cardiovascular coronary artery
C0343692|Syphilitic coronary artery disease (diagnosis)
C0343692|Late quaternary syphilitic coronary artery disease
C0343692|Syphilitic coronary artery disease (disorder)
C2939120|Coronary artery fistula
C2939120|Congenital coronary artery fistula
C2939120|Congenital coronary artery fistula (disorder)
C0519097|aneurysm of left ventricle
C0519097|aneurysm of left ventricle (diagnosis)
C0519097|left ventricular aneurysm
C0519097|Left ventricular aneurysm (disorder)
C0519097|LV wall aneurysmal
C0519097|Left ventricular wall aneurysmal
C0519097|LVA - Left ventricular aneurysm
C0340678|Coronary steal syndrome
C0340678|Coronary steal syndrome (disorder)
C0264688|coronary (artery) rupture
C0264688|Rupture;artery;coronary
C0264688|Coronary artery rupture
C0264688|Coronary artery rupture (disorder)
C0264699|acute anteroseptal myocardial infarction (diagnosis)
C0264699|acute anteroseptal myocardial infarction
C0264699|Acute antero septal myocardial infarction
C0264699|Acute anteroseptal myocardial infarction (disorder)
C0264699|Acute myocardial infarction, anteroseptal
C0264700|acute myocardial infarction of inferior wall (diagnosis)
C0264700|acute inferior wall MI
C0264700|acute myocardial infarction of inferior wall
C0264700|Acute Inferior Myocardial Infarction
C0264700|Acute myocardial infarction of diaphragmatic wall
C0264700|Acute myocardial infarction of inferior wall (disorder)
C0264700|Acute myocardial infarction of inferior wall, NOS
C0264700|Infarction, diaphragmatic wall NOS
C0264700|Acute myocardial infarction, diaphragmatic wall NOS
C0264700|Acute myocardial infarction, inferior wall NOS
C0345117|Abnormal coronary orifice (disorder)
C0345117|Abnormal coronary orifice
C0340892|Mechanical complication of coronary bypass
C0340892|Mechanical complication of coronary bypass (disorder)
C0275847|syphilitic ostial coronary artery disease
C0275847|syphilis cardiovascular coronary artery ostial
C0275847|syphilitic ostial coronary artery disease (diagnosis)
C0275847|Syphilitic ostial coronary disease
C0275847|Syphilitic ostial coronary disease (disorder)
C0221359|Anomalous origin of coronary artery (diagnosis)
C0221359|Anomalous origin of coronary artery
C0221359|congenital anomaly of coronary artery of anomalous origin
C0221359|Anomalous coronary artery origin
C0221359|Anomalous origin of coronary artery (disorder)
C0151814|coronary occlusion
C0151814|Coronary artery occlusion
C0151814|Occlusions, Coronary
C0151814|Coronary Occlusions
C0151814|Occlusion, Coronary
C0151814|coronary (artery) occlusion
C0151814|Coronary Occlusion [Disease/Finding]
C0151814|Occlusion;coronary
C0151814|coronary artery occlusion (diagnosis)
C0151814|Occlusion coronary
C0151814|Occlusion coronary artery
C0151814|Coronary artery occluded
C0151814|Coronary occlusion (disorder)
C0151814|Coronary occlusion, NOS
C0151814|Coronary occlusion NOS
C0340297|acute myocardial infarction of septal wall (diagnosis)
C0340297|acute myocardial infarction of septal wall
C0340297|Acute myocardial infarction of septum
C0340297|Acute myocardial infarction of septum alone
C0340297|Acute septal infarction
C0340297|Acute myocardial infarction of septum (disorder)
C0340297|Infarction of septum alone
C3695002|coronary artery disease in transplanted heart (diagnosis)
C3695002|coronary artery disease in transplanted heart
C3697310|Increase in velocity of coronary artery of fetus
C3697310|Increase in velocity of coronary artery of fetus (disorder)
C1834751|CORONARY ARTERY DISEASE, DEVELOPMENT OF, IN HIV
C1859728|CORONARY SCLEROSIS, MEDIAL, OF INFANCY
C2063729|multiple coronary aneurysms
C2063729|multiple coronary aneurysms (diagnosis)
C0027051|Infarctions, Myocardial
C0027051|Myocardial Infarction
C0027051|Myocardial Infarctions
C0027051|Infarcts, Myocardial
C0027051|Myocardial Infarcts
C0027051|Infarct, Myocardial
C0027051|Infarction, Myocardial
C0027051|MI
C0027051|Myocardial infarction (MI)
C0027051|heart attack
C0027051|cardiac infarction
C0027051|Myocardial Infarction [Disease/Finding]
C0027051|Myocardial Infarct
C0027051|Infarction;heart
C0027051|Infarction;myocardial
C0027051|Attack - heart
C0027051|MI - Myocardial infarction
C0027051|Myocardial infarction (disorder)
C0027051|Cardiac infarct
C0027051|myocardial infarction (diagnosis)
C0027051|-- Heart Attack
C0027051|Cardiovascular Strokes
C0027051|Stroke, Cardiovascular
C0027051|Strokes, Cardiovascular
C0027051|Cardiovascular Stroke
C0027051|MI, Myocardial Infarction
C0027051|Myocardial Infarction, (MI)
C0027051|Infarction (MI), Myocardial
C0027051|Heart Attacks
C0027051|Attack coronary
C0027051|Attack heart (NOS)
C0027051|Infarct myocardial
C0027051|Cardio/pulm: Myocardial infarction
C0027051|Infarction of heart
C0027051|cardiac; infarction
C0027051|infarction; myocardial
C0027051|Cardiac infarction, NOS
C0027051|Heart attack, NOS
C0027051|Infarction of heart, NOS
C0027051|Myocardial infarction, NOS
C0027051|Infarctions (Myocardial)
C0027051|Myocardial infarction NOS
C0027051|heart infarction
C3165030|Systemic to pulmonary collateral from coronary artery
C3165030|Systemic to pulmonary collateral artery from coronary artery (disorder)
C3165030|Systemic to pulmonary collateral from coronary artery (disorder)
C3165030|Systemic to pulmonary collateral artery from coronary artery
C4020725|Non-occlusive coronary artery disease
C4020725|Nonocclusive coronary artery disease
C4020725|Non-occlusive coronary artery stenosis
C2676505|Post-angioplasty coronary artery restenosis
C4047786|Thrombosis of left circumflex artery
C4047786|Thrombosis of left circumflex artery (disorder)
C4075502|Abnormal ostium of coronary artery
C4075502|Abnormal ostium of coronary artery (disorder)
C1299363|Bifurcation lesion of coronary artery
C1299363|Bifurcation lesion of coronary artery (disorder)
C1299363|Bifurcation lesion of coronary artery (finding)
C0265898|Coronary artery fistula
C0265898|Coronary artery fistula (disorder)
