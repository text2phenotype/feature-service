C1953564|Hep C Virus Ab
C1953564|HCV Ab
C1953564|HCV Antibodies
C1953564|HCV Antibody Test
C1953564|Hepatitis C Virus (HCV) Antibody
C1953564|Hepatitis C virus Ab
C1953564|Hepatitis C virus Ab Signal
C1953564|Hepatitis C virus Antibody Signal
C1953564|Hepatitis C virus Antibody Test
C1953564|TEST 140659
C1953564|LOINC 48159-8
C1953564|LNC 48159-8