C0942407|T201|Laboratory studies:Cmplx:-:^Patient:Set|
C0942407|T201|Laboratory studies (set)|
C0942407|T201|Laboratory studies:Complex:-:^Patient:Set|
C0802029|T201|Collection duration of Urine|
C0802029|T201|Collect duration Time Ur|
C0802029|T201|Collection duration:Time:*:Urine:Qn|
C0802029|T201|Collection duration:Time:LIFE OF THE UNIT:Urine:Quantitative|
C1114758|T201|Dose #|
C1114758|T201|Dose number|
C1114758|T201|Dose number:Num:Pt:^Patient:Qn|
C1114758|T201|Dose number:Number:Point in time:^Patient:Quantitative|
C1317013|T201|2D echocardiogram panel:-:Pt:^Patient:-|
C1317013|T201|2D echocardiogram panel|
C1317013|T201|2D Echo Pnl|
C1317013|T201|2D echocardiogram panel:-:Point in time:^Patient:-|
C0363876|T201|Alanine aminotransferase:CCnc:Pt:Ser/Plas:Qn|
C0363876|T201|Alanine aminotransferase [Enzymatic activity/volume] in Serum or Plasma|
C0363876|T201|ALT SerPl-cCnc|
C0363876|T201|Alanine aminotransferase:Catalytic Concentration:Point in time:Serum/Plasma:Quantitative|
C1551702|T098|Alexander|
C0363885|T201|Albumin SerPl-mCnc|
C0363885|T201|Albumin:MCnc:Pt:Ser/Plas:Qn|
C0363885|T201|Albumin [Mass/volume] in Serum or Plasma|
C0363885|T201|Albumin:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1551711|T098|Chickaloon|
C0363888|T201|Albumin [Mass/volume] in Urine|
C0363888|T201|Albumin Ur-mCnc|
C0363888|T201|Albumin:MCnc:Pt:Urine:Qn|
C0363888|T201|Albumin:Mass Concentration:Point in time:Urine:Quantitative|
C1551714|T098|Circle|
C0801090|T201|Ejection time:Time:Point in time:Aortic valve:Quantitative:Ultrasound.doppler|
C0801090|T201|Ejection time:Time:Pt:Aortic valve:Qn:US.doppler|
C0801090|T201|AV Ejection time DOP|
C0801090|T201|Aortic valve Ejection time by US.doppler|
C0550189|T201|Alkaline phosphatase isoenzyme:ACnc:Pt:Ser/Plas:Qn|
C0550189|T201|Alkaline phosphatase isoenzyme [Units/volume] in Serum or Plasma|
C0550189|T201|ALP Iso SerPl-aCnc|
C0550189|T201|Alkaline phosphatase isoenzyme:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative|
C0484638|T201|Alkaline phosphatase [Enzymatic activity/volume] in Serum or Plasma|
C0484638|T201|ALP SerPl-cCnc|
C0484638|T201|Alkaline phosphatase:CCnc:Pt:Ser/Plas:Qn|
C0484638|T201|Alkaline phosphatase:Catalytic Concentration:Point in time:Serum/Plasma:Quantitative|
C0484660|T201|Anion Gap3 SerPl-sCnc|
C0484660|T201|Anion gap 3:SCnc:Pt:Ser/Plas:Qn|
C0484660|T201|Anion gap 3 in Serum or Plasma|
C0484660|T201|Anion gap 3:Substance Concentration:Point in time:Serum/Plasma:Quantitative|
C0364055|T201|Aspartate aminotransferase:CCnc:Pt:Ser/Plas:Qn|
C0364055|T201|Aspartate aminotransferase [Enzymatic activity/volume] in Serum or Plasma|
C0364055|T201|AST SerPl-cCnc|
C0364055|T201|Aspartate aminotransferase:Catalytic Concentration:Point in time:Serum/Plasma:Quantitative|
C1551869|T098|Iqurmuit (Russian Mission)|
C0801138|T201|AV Orifice Area US|
C0801138|T201|Orifice:Area:Pt:Aortic valve:Qn:US|
C0801138|T201|Aortic valve Orifice [Area] by US|
C0801138|T201|Orifice:Area:Point in time:Aortic valve:Quantitative:Ultrasound|
C0362894|T201|Basophils/100 leukocytes:NFr:Pt:Bld:Qn:Automated count|
C0362894|T201|Basophils/100 leukocytes in Blood by Automated count|
C0362894|T201|Basophils/100 leukocytes:Number Fraction:Point in time:Whole blood:Quantitative:Automated count|
C0362894|T201|Basophils/leuk NFr Bld Auto|
C0362892|T201|Basophils:NCnc:Pt:Bld:Qn:Automated count|
C0362892|T201|Basophils [#/volume] in Blood by Automated count|
C0362892|T201|Basophils # Bld Auto|
C0362892|T201|Basophils:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0881599|T201|Bas Metab 2000 Pnl SerPl|
C0881599|T201|Basic metabolic 2000 panel:-:Pt:Ser/Plas:Qn|
C0881599|T201|Basic metabolic 2000 panel:-:Point in time:Serum/Plasma:Quantitative|
C0881599|T201|Basic metabolic 2000 panel - Serum or Plasma|
C2360771|T201|Basic metabolic panel:-:Pt:Bld:Qn|
C2360771|T201|Bas Metab Pnl Bld|
C2360771|T201|Basic metabolic panel:-:Point in time:Whole blood:Quantitative|
C2360771|T201|Basic metabolic panel - Blood|
C0797802|T201|Bicarbonate:SCnc:Pt:BldV:Qn|
C0797802|T201|Bicarbonate [Moles/volume] in Venous blood|
C0797802|T201|HCO3 BldV-sCnc|
C0797802|T201|Bicarbonate:Substance Concentration:Point in time:Blood venous:Quantitative|
C0798323|T201|Bilirub Conj SerPl-mCnc|
C0798323|T201|Bilirubin.glucuronidated:MCnc:Pt:Ser/Plas:Qn|
C0798323|T201|Bilirubin.glucuronidated:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0798323|T201|Bilirubin.conjugated [Mass/volume] in Serum or Plasma|
C0364108|T201|Bilirub SerPl-mCnc|
C0364108|T201|Bilirubin:MCnc:Pt:Ser/Plas:Qn|
C0364108|T201|Bilirubin.total [Mass/volume] in Serum or Plasma|
C0364108|T201|Bilirubin:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1553276|T098|Egegik|
C0365237|T201|Urea nitrogen [Mass/volume] in Blood|
C0365237|T201|BUN Bld-mCnc|
C0365237|T201|Urea nitrogen:MCnc:Pt:Bld:Qn|
C0365237|T201|Urea nitrogen:Mass Concentration:Point in time:Whole blood:Quantitative|
C0365240|T201|Urea nitrogen:MCnc:Pt:Ser/Plas:Qn|
C0365240|T201|Urea nitrogen [Mass/volume] in Serum or Plasma|
C0365240|T201|BUN SerPl-mCnc|
C0365240|T201|Urea nitrogen:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0800968|T201|Calcium SerPl-mCnc|
C0800968|T201|Calcium [Mass/volume] in Serum or Plasma|
C0800968|T201|Calcium:MCnc:Pt:Ser/Plas:Qn|
C0800968|T201|Calcium:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0516831|T033|Breastfeeding Maintenance|
C0231528|T184|muscle aches, generalized (myalgias)|
C0231528|T184|generalized myalgia|
C0231528|T184|generalized muscle aches|
C0231528|T184|generalized muscle aches (symptom)|
C0723022|T121|Renovist|
C0723022|T130|Renovist|
C0723022|T109|Renovist|
C0995472|T007|Flexibacter roseolus Lewin 1969|
C0995472|T007|Flexibacter roseolus|
C1552038|T078|African Religions|
C0364160|T201|CO2 SerPl-sCnc|
C0364160|T201|Carbon dioxide, total [Moles/volume] in Serum or Plasma|
C0364160|T201|Carbon dioxide:SCnc:Pt:Ser/Plas:Qn|
C0364160|T201|Carbon dioxide:Substance Concentration:Point in time:Serum/Plasma:Quantitative|
C0078988|T098|Asian|
C0803374|T201|Carbon dioxide, total [Moles/volume] in Blood|
C0803374|T201|CO2 Bld-sCnc|
C0803374|T201|Carbon dioxide:SCnc:Pt:Bld:Qn|
C0803374|T201|Carbon dioxide:Substance Concentration:Point in time:Whole blood:Quantitative|
C0364201|T201|Chloride Bld-sCnc|
C0364201|T201|Chloride [Moles/volume] in Blood|
C0364201|T201|Chloride:SCnc:Pt:Bld:Qn|
C0364201|T201|Chloride:Substance Concentration:Point in time:Whole blood:Quantitative|
C1328872|T098|Dominican|
C1553338|T098|Dominican|
C0364207|T201|Chloride [Moles/volume] in Serum or Plasma|
C0364207|T201|Chloride SerPl-sCnc|
C0364207|T201|Chloride:SCnc:Pt:Ser/Plas:Qn|
C0364207|T201|Chloride:Substance Concentration:Point in time:Serum/Plasma:Quantitative|
C0425373|T098|West Indian|
C1526484|T201|Creatinine [Mass/volume] in Blood|
C1526484|T201|Creat Bld-mCnc|
C1526484|T201|Creatinine:MCnc:Pt:Bld:Qn|
C1526484|T201|Creatinine:Mass Concentration:Point in time:Whole blood:Quantitative|
C1507825|T201|Creatinine:MCnc:XXX:Urine:Qn|
C1507825|T201|Creat ?Tm Ur-mCnc|
C1507825|T201|Creatinine:Mass Concentration:time reported elsewhere:Urine:Quantitative|
C1507825|T201|Creatinine [Mass/volume] in Urine collected for unspecified duration|
C0364294|T201|Creat SerPl-mCnc|
C0364294|T201|Creatinine:MCnc:Pt:Ser/Plas:Qn|
C0364294|T201|Creatinine [Mass/volume] in Serum or Plasma|
C0364294|T201|Creatinine:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1171359|T098|Panamanian|
C1316996|T201|12 Channel EKG Pnl|
C1316996|T201|EKG 12 channel panel:-:Pt:Heart:-:EKG|
C1316996|T201|EKG 12 channel panel|
C1316996|T201|EKG 12 channel panel:-:Point in time:Heart:-:EKG|
C0801842|T201|EKG impression:Imp:Pt:Heart:Nar:EKG|
C0801842|T201|EKG impression|
C0801842|T201|EKG impression:Impression/interpretation of study:Point in time:Heart:Narrative:EKG|
C0801842|T201|EKG impression Narrative|
C0362902|T201|Eosinophils/100 leukocytes:NFr:Pt:Bld:Qn:Automated count|
C0362902|T201|Eosinophils/100 leukocytes in Blood by Automated count|
C0362902|T201|Eosinophils/100 leukocytes:Number Fraction:Point in time:Whole blood:Quantitative:Automated count|
C0362902|T201|Eosinophil/leuk NFr Bld Auto|
C0362900|T201|Eosinophils [#/volume] in Blood by Automated count|
C0362900|T201|Eosinophils:NCnc:Pt:Bld:Qn:Automated count|
C0362900|T201|Eosinophil # Bld Auto|
C0362900|T201|Eosinophils:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0362910|T201|RBC # Bld Auto|
C0362910|T201|Erythrocytes:NCnc:Pt:Bld:Qn:Automated count|
C0362910|T201|Erythrocytes [#/volume] in Blood by Automated count|
C0362910|T201|Erythrocytes:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0362908|T201|Erythrocyte mean corpuscular volume [Entitic volume] by Automated count|
C0362908|T201|MCV RBC Auto|
C0362908|T201|Erythrocyte mean corpuscular volume:EntVol:Pt:RBC:Qn:Automated count|
C0362908|T201|Erythrocyte mean corpuscular volume:Entitic Volume:Point in time:Erythrocytes:Quantitative:Automated count|
C0362906|T201|Erythrocyte mean corpuscular hemoglobin [Entitic mass] by Automated count|
C0362906|T201|MCH RBC Qn Auto|
C0362906|T201|Erythrocyte mean corpuscular hemoglobin:EntMass:Pt:RBC:Qn:Automated count|
C0362906|T201|Erythrocyte mean corpuscular hemoglobin:Entitic Mass:Point in time:Erythrocytes:Quantitative:Automated count|
C0362907|T201|MCHC RBC Auto-mCnc|
C0362907|T201|Erythrocyte mean corpuscular hemoglobin concentration [Mass/volume] by Automated count|
C0362907|T201|Erythrocyte mean corpuscular hemoglobin concentration:MCnc:Pt:RBC:Qn:Automated count|
C0362907|T201|Erythrocyte mean corpuscular hemoglobin concentration:Mass Concentration:Point in time:Erythrocytes:Quantitative:Automated count|
C0362909|T201|Erythrocyte distribution width:Ratio:Pt:RBC:Qn:Automated count|
C0362909|T201|RDW RBC Auto-Rto|
C0362909|T201|Erythrocyte distribution width [Ratio] by Automated count|
C0362909|T201|Erythrocyte distribution width:Ratio:Point in time:Erythrocytes:Quantitative:Automated count|
C1114251|T201|Erythrocytes.nucleated:NCnc:Pt:Bld:Qn|
C1114251|T201|nRBC # Bld|
C1114251|T201|Nucleated erythrocytes [#/volume] in Blood|
C1114251|T201|Erythrocytes.nucleated:Number Concentration (count/vol):Point in time:Whole blood:Quantitative|
C0945356|T201|Nucleated erythrocytes/100 erythrocytes in Blood|
C0945356|T201|Erythrocytes.nucleated/100 erythrocytes:NFr:Pt:Bld:Qn|
C0945356|T201|Erythrocytes.nucleated/100 erythrocytes:Number Fraction:Point in time:Whole blood:Quantitative|
C0945356|T201|nRBC/100 RBC NFr Bld|
C0364459|T201|GGT SerPl-cCnc|
C0364459|T201|Gamma glutamyl transferase [Enzymatic activity/volume] in Serum or Plasma|
C0364459|T201|Gamma glutamyl transferase:CCnc:Pt:Ser/Plas:Qn|
C0364459|T201|Gamma glutamyl transferase:Catalytic Concentration:Point in time:Serum/Plasma:Quantitative|
C0364479|T201|Glucose:MCnc:Pt:Bld:Qn|
C0364479|T201|Glucose [Mass/volume] in Blood|
C0364479|T201|Glucose Bld-mCnc|
C0364479|T201|Glucose:Mass Concentration:Point in time:Whole blood:Quantitative|
C0484731|T201|Glucose:MCnc:Pt:Ser/Plas:Qn|
C0484731|T201|Glucose SerPl-mCnc|
C0484731|T201|Glucose [Mass/volume] in Serum or Plasma|
C0484731|T201|Glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C2718131|T201|Deprecated Glucose [Mass/volume] in Serum or Plasma|
C2718131|T201|Deprecated Glucose SerPl-mCnc|
C2718131|T201|Glucose:MCnc:Pt:Ser/Plas:Qn|
C2718131|T201|Glucose:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0364474|T201|Globulin Ser-mCnc|
C0364474|T201|Globulin:MCnc:Pt:Ser:Qn|
C0364474|T201|Globulin [Mass/volume] in Serum|
C0364474|T201|Globulin:Mass Concentration:Point in time:Serum:Quantitative|
C1316377|T201|GFR/BSA.pred SerPl MDRD-ArVRat|
C1316377|T201|Glomerular filtration rate/1.73 sq M.predicted:ArVRat:Pt:Ser/Plas:Qn:Creatinine-based formula (MDRD)|
C1316377|T201|Glomerular filtration rate/1.73 sq M.predicted:Volume Rate/Area:Point in time:Serum/Plasma:Quantitative:Creatinine-based formula (MDRD)|
C1316377|T201|Glomerular filtration rate/1.73 sq M.predicted [Volume Rate/Area] in Serum or Plasma by Creatinine-based formula (MDRD)|
C1114184|T201|Hgb BldA-mCnc|
C1114184|T201|Hemoglobin [Mass/volume] in Arterial blood|
C1114184|T201|Hemoglobin:MCnc:Pt:BldA:Qn|
C1114184|T201|Hemoglobin:Mass Concentration:Point in time:Blood arterial:Quantitative|
C0362923|T201|Hemoglobin:MCnc:Pt:Bld:Qn|
C0362923|T201|Hemoglobin [Mass/volume] in Blood|
C0362923|T201|Hgb Bld-mCnc|
C0362923|T201|Hemoglobin:Mass Concentration:Point in time:Whole blood:Quantitative|
C0366781|T201|Hemoglobin A1c/Hemoglobin.total in Blood|
C0366781|T201|Hgb A1c MFr Bld|
C0366781|T201|Hemoglobin A1c/Hemoglobin.total:MFr:Pt:Bld:Qn|
C0366781|T201|Hemoglobin A1c/Hemoglobin.total:Mass Fraction:Point in time:Whole blood:Quantitative|
C0364473|T201|Hemoglobin.gastrointestinal [Presence] in Stool|
C0364473|T201|Hemoglobin.gastrointestinal:ACnc:Pt:Stool:Ord|
C0364473|T201|Hemoglobin.gastrointestinal:Arbitrary Concentration:Point in time:Stool = Fecal:Ordinal|
C0364473|T201|Hemoccult Stl Ql|
C0803379|T201|Hematocrit:VFr:Pt:Bld:Qn|
C0803379|T201|Hematocrit [Volume Fraction] of Blood|
C0803379|T201|Hct VFr Bld|
C0803379|T201|Hematocrit:Volume Fraction:Point in time:Whole blood:Quantitative|
C0366777|T201|Hematocrit [Volume Fraction] of Blood by Automated count|
C0366777|T201|Hematocrit:VFr:Pt:Bld:Qn:Automated count|
C0366777|T201|Hct VFr Bld Auto|
C0366777|T201|Hematocrit:Volume Fraction:Point in time:Whole blood:Quantitative:Automated count|
C0482691|T201|INR in Platelet poor plasma by Coagulation assay|
C0482691|T201|INR PPP|
C0482691|T201|Coagulation tissue factor induced.INR:RelTime:Pt:PPP:Qn:Coag|
C0482691|T201|Coagulation tissue factor induced.INR:Relative Time:Point in time:Platelet poor plasma:Quantitative:Coagulation Assay|
C0364674|T201|Lactate dehydrogenase [Enzymatic activity/volume] in Serum or Plasma|
C0364674|T201|Lactate dehydrogenase:CCnc:Pt:Ser/Plas:Qn|
C0364674|T201|LDH SerPl-cCnc|
C0364674|T201|Lactate dehydrogenase:Catalytic Concentration:Point in time:Serum/Plasma:Quantitative|
C0362952|T201|Lymphocytes/100 leukocytes:NFr:Pt:Bld:Qn:Automated count|
C0362952|T201|Lymphocytes/100 leukocytes in Blood by Automated count|
C0362952|T201|Lymphocytes/100 leukocytes:Number Fraction:Point in time:Whole blood:Quantitative:Automated count|
C0362952|T201|Lymphocytes/leuk NFr Bld Auto|
C0362947|T201|Lymphocytes # Bld Auto|
C0362947|T201|Lymphocytes:NCnc:Pt:Bld:Qn:Automated count|
C0362947|T201|Lymphocytes [#/volume] in Blood by Automated count|
C0362947|T201|Lymphocytes:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0364961|T201|Potassium:SCnc:Pt:Bld:Qn|
C0364961|T201|Potassium Bld-sCnc|
C0364961|T201|Potassium [Moles/volume] in Blood|
C0364961|T201|Potassium:Substance Concentration:Point in time:Whole blood:Quantitative|
C0882319|T201|Potassium [Mass/volume] in Serum or Plasma|
C0882319|T201|Potassium:MCnc:Pt:Ser/Plas:Qn|
C0882319|T201|Potassium SerPl-mCnc|
C0882319|T201|Potassium:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0364968|T201|Potassium:SCnc:Pt:Ser/Plas:Qn|
C0364968|T201|Potassium [Moles/volume] in Serum or Plasma|
C0364968|T201|Potassium SerPl-sCnc|
C0364968|T201|Potassium:Substance Concentration:Point in time:Serum/Plasma:Quantitative|
C0942474|T201|Platelets [#/volume] in Blood|
C0942474|T201|Platelets:NCnc:Pt:Bld:Qn|
C0942474|T201|Platelet # Bld|
C0942474|T201|Platelets:Number Concentration (count/vol):Point in time:Whole blood:Quantitative|
C1370010|T201|Phosphate [Mass/volume] in Serum or Plasma|
C1370010|T201|Phosphate:MCnc:Pt:Ser/Plas:Qn|
C1370010|T201|Phosphate SerPl-mCnc|
C1370010|T201|Phosphate:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0365029|T201|Protein [Mass/volume] in Serum or Plasma|
C0365029|T201|Prot SerPl-mCnc|
C0365029|T201|Protein:MCnc:Pt:Ser/Plas:Qn|
C0365029|T201|Protein:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0362960|T201|Monocytes/100 leukocytes:NFr:Pt:Bld:Qn:Automated count|
C0362960|T201|Monocytes/100 leukocytes in Blood by Automated count|
C0362960|T201|Monocytes/100 leukocytes:Number Fraction:Point in time:Whole blood:Quantitative:Automated count|
C0362960|T201|Monocytes/leuk NFr Bld Auto|
C0362958|T201|Monocytes:NCnc:Pt:Bld:Qn:Automated count|
C0362958|T201|Monocytes # Bld Auto|
C0362958|T201|Monocytes [#/volume] in Blood by Automated count|
C0362958|T201|Monocytes:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0798130|T201|Microalbumin [Mass/volume] in Urine|
C0798130|T201|Microalbumin Ur-mCnc|
C0798130|T201|Albumin:MCnc:Pt:Urine:Qn:Detection limit <= 20 mg/L|
C0798130|T201|Albumin:Mass Concentration:Point in time:Urine:Quantitative:Detection limit <= 20 mg/L|
C0798132|T201|Microalbumin/Creat Ur|
C0798132|T201|Microalbumin/Creatinine [Mass Ratio] in Urine|
C0798132|T201|Albumin/Creatinine:MRto:Pt:Urine:Qn:Detection limit <= 20 mg/L|
C0798132|T201|Albumin/Creatinine:Mass Ratio:Point in time:Urine:Quantitative:Detection limit <= 20 mg/L|
C0365091|T201|Sodium:SCnc:Pt:Bld:Qn|
C0365091|T201|Sodium [Moles/volume] in Blood|
C0365091|T201|Sodium Bld-sCnc|
C0365091|T201|Sodium:Substance Concentration:Point in time:Whole blood:Quantitative|
C0365095|T201|Sodium:SCnc:Pt:Ser/Plas:Qn|
C0365095|T201|Sodium [Moles/volume] in Serum or Plasma|
C0365095|T201|Sodium SerPl-sCnc|
C0365095|T201|Sodium:Substance Concentration:Point in time:Serum/Plasma:Quantitative|
C0362987|T201|Neutrophils/100 leukocytes in Blood by Automated count|
C0362987|T201|Neutrophils/100 leukocytes:NFr:Pt:Bld:Qn:Automated count|
C0362987|T201|Neutrophils/100 leukocytes:Number Fraction:Point in time:Whole blood:Quantitative:Automated count|
C0362987|T201|Neutrophils/leuk NFr Bld Auto|
C0362968|T201|Neutrophils:NCnc:Pt:Bld:Qn:Automated count|
C0362968|T201|Neutrophils [#/volume] in Blood by Automated count|
C0362968|T201|Neutrophils # Bld Auto|
C0362968|T201|Neutrophils:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0368556|T201|Bacteria identified:Prid:Pt:Sputum:Nom:Culture|
C0368556|T201|Bacteria identified in Sputum by Culture|
C0368556|T201|Bacteria Spt Cult|
C0368556|T201|Bacteria identified:Presence or Identity:Point in time:Sputum:Nominal:Culture|
C0484851|T201|Troponin T.cardiac [Mass/volume] in Serum or Plasma|
C0484851|T201|Troponin T SerPl-mCnc|
C0484851|T201|Troponin T.cardiac:MCnc:Pt:Ser/Plas:Qn|
C0484851|T201|Troponin T.cardiac:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1542867|T201|Body mass index (BMI) [Ratio]|
C1542867|T201|Body mass index:Ratio:Pt:^Patient:Qn|
C1542867|T201|BMI|
C1542867|T201|Body mass index:Ratio:Point in time:^Patient:Quantitative|
C0365284|T201|BSA Derived|
C0365284|T201|Body surface area Derived from formula|
C0365284|T201|Body surface:Area:Pt:^Patient:Qn:Derived|
C0365284|T201|Body surface:Area:Point in time:^Patient:Quantitative:Derived|
C0365286|T201|Body weight Measured|
C0365286|T201|Body weight:Mass:Pt:^Patient:Qn:Measured|
C0365286|T201|Weight Measured|
C0365286|T201|Body weight:Mass:Point in time:^Patient:Quantitative:Measured|
C0944911|T201|Body weight:Mass:Pt:^Patient:Qn|
C0944911|T201|Weight|
C0944911|T201|Body weight|
C0944911|T201|Body weight:Mass:Point in time:^Patient:Quantitative|
C1648313|T201|Body mass index:Ratio:Pt:^Patient:Qn:Calculated|
C1648313|T201|Deprecated BMI|
C1648313|T201|Deprecated Body mass index (BMI)|
C1648313|T201|Body mass index:Ratio:Point in time:^Patient:Quantitative:Calculated|
C0487995|T201|Body temperature:Temp:Pt:^Patient:Qn|
C0487995|T201|Body temperature|
C0487995|T201|Body temperature:Temperature:Point in time:^Patient:Quantitative|
C0487973|T201|Circumference.occipital-frontal:Len:Pt:Head:Qn:Tape measure|
C0487973|T201|Head Occipital-frontal circumference by Tape measure|
C0487973|T201|Circumference.occipital-frontal:Length:Point in time:Head:Quantitative:Tape measure|
C0487973|T201|Head Circumf OFC by Tape measure|
C0488794|T201|Heart rate|
C0488794|T201|Heart rate:NRat:Pt:XXX:Qn|
C0488794|T201|Heart rate:Number = Count/Time:Point in time:To be specified in another part of the message:Quantitative|
C0487985|T201|Body height|
C0487985|T201|Body height:Len:Pt:^Patient:Qn|
C0487985|T201|Body height:Length:Point in time:^Patient:Quantitative|
C0487988|T201|Body height^lying:Len:Pt:^Patient:Qn|
C0487988|T201|Body height --lying|
C0487988|T201|Body height^lying:Length:Point in time:^Patient:Quantitative|
C0487988|T201|Body height lying|
C0489258|T201|Breaths:NRat:Pt:Respiratory system:Qn|
C0489258|T201|Respiratory rate|
C0489258|T201|Breaths:Number = Count/Time:Point in time:Respiratory system:Quantitative|
C0489258|T201|Resp rate|
C0797821|T201|Cholesterol.in HDL:SCnc:Pt:Ser/Plas:Qn|
C0797821|T201|Cholesterol in HDL [Moles/volume] in Serum or Plasma|
C0797821|T201|HDLc SerPl-sCnc|
C0797821|T201|Cholesterol.in HDL:Substance Concentration:Point in time:Serum/Plasma:Quantitative|
C0364225|T201|Cholesterol in LDL [Mass/volume] in Serum or Plasma|
C0364225|T201|Cholesterol.in LDL:MCnc:Pt:Ser/Plas:Qn|
C0364225|T201|LDLc SerPl-mCnc|
C0364225|T201|Cholesterol.in LDL:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1553344|T098|Mariana Islander|
C0364708|T201|Cholesterol:MCnc:Pt:Ser/Plas:Qn|
C0364708|T201|Cholest SerPl-mCnc|
C0364708|T201|Cholesterol [Mass/volume] in Serum or Plasma|
C0364708|T201|Cholesterol:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1553346|T098|Kosraean|
C0364221|T201|Cholesterol.in HDL:MCnc:Pt:Ser/Plas:Qn|
C0364221|T201|Cholesterol in HDL [Mass/volume] in Serum or Plasma|
C0364221|T201|HDLc SerPl-mCnc|
C0364221|T201|Cholesterol.in HDL:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1556099|T098|Micronesian|
C0550534|T201|Triglyceride:MCnc:Pt:Ser/Plas:Qn:Calculated|
C0550534|T201|Triglyceride [Mass/volume] in Serum or Plasma by calculation|
C0550534|T201|Trigl SerPl Calc-mCnc|
C0550534|T201|Triglyceride:Mass Concentration:Point in time:Serum/Plasma:Quantitative:Calculated|
C0364714|T201|Trigl SerPl-mCnc|
C0364714|T201|Triglyceride:MCnc:Pt:Ser/Plas:Qn|
C0364714|T201|Triglyceride [Mass/volume] in Serum or Plasma|
C0364714|T201|Triglyceride:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C1316229|T201|WBC # Pheresis BPU Auto|
C1316229|T201|Leukocytes:NCnc:Pt:^BPU.platelet pheresis:Qn:Automated count|
C1316229|T201|Leukocytes [#/volume] in Blood Product unit.platelet pheresis by Automated count|
C1316229|T201|Leukocytes:Number Concentration (count/vol):Point in time:^Blood product unit (Pack).platelet pheresis:Quantitative:Automated count|
C0945357|T201|Leukocytes:NCnc:Pt:Bld:Qn|
C0945357|T201|Leukocytes [#/volume] in Blood|
C0945357|T201|WBC # Bld|
C0945357|T201|Leukocytes:Number Concentration (count/vol):Point in time:Whole blood:Quantitative|
C0484430|T201|Leukocytes [#/volume] in Blood by Automated count|
C0484430|T201|Leukocytes:NCnc:Pt:Bld:Qn:Automated count|
C0484430|T201|WBC # Bld Auto|
C0484430|T201|Leukocytes:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0488052|T201|Intravascular diastolic:Pres:Pt:Arterial system:Qn|
C0488052|T201|Diastolic blood pressure|
C0488052|T201|BP dias|
C0488052|T201|Intravascular diastolic:Pressure:Point in time:Arterial system:Quantitative|
C0488055|T201|Intravascular systolic:Pres:Pt:Arterial system:Qn|
C0488055|T201|Systolic blood pressure|
C0488055|T201|BP sys|
C0488055|T201|Intravascular systolic:Pressure:Point in time:Arterial system:Quantitative|
C1114363|T201|C reactive protein [Mass/volume] in Serum or Plasma by High sensitivity method|
C1114363|T201|C reactive protein:MCnc:Pt:Ser/Plas:Qn:High sensitivity|
C1114363|T201|CRP SerPl HS-mCnc|
C1114363|T201|C reactive protein:Mass Concentration:Point in time:Serum/Plasma:Quantitative:High sensitivity|
C0484872|T201|Microscopic observation:Prid:Pt:Cvx:Nom:Cyto stain|
C0484872|T201|Microscopic observation [Identifier] in Cervix by Cyto stain|
C0484872|T201|Cyto Cervix|
C0484872|T201|Microscopic observation:Presence or Identity:Point in time:Cervix:Nominal:Cytology Stain|
C1147461|T201|C trach Ag XXX Ql|
C1147461|T201|Chlamydia trachomatis Ag:ACnc:Pt:XXX:Ord|
C1147461|T201|Chlamydia trachomatis Ag [Presence] in Unspecified specimen|
C1147461|T201|Chlamydia trachomatis Antigen:Arbitrary Concentration:Point in time:To be specified in another part of the message:Ordinal|
C1978488|T201|Protein [Mass/volume] in Urine by Automated test strip|
C1978488|T201|Prot Ur Strip.auto-mCnc|
C1978488|T201|Protein:MCnc:Pt:Urine:Qn:Test strip.automated|
C1978488|T201|Protein:Mass Concentration:Point in time:Urine:Quantitative:Test strip.automated|
C0364239|T201|HCG SerPl-sCnc|
C0364239|T201|Choriogonadotropin [Moles/volume] in Serum or Plasma|
C0364239|T201|Choriogonadotropin:SCnc:Pt:Ser/Plas:Qn|
C0364239|T201|Choriogonadotropin:Substance Concentration:Point in time:Serum/Plasma:Quantitative|
C1553354|T098|Assyrian|
C3654136|T201|HIV1+2 IgG Bld Ql EIA.rapid|
C3654136|T201|HIV 1+2 Ab.IgG:Threshold:Pt:Bld:Ord:EIA.rapid|
C3654136|T201|human immunodeficiency virus 1+2 Antibody.immunoglobulin G:Threshold:Point in time:Whole blood:Ordinal:Enzyme Immunoassay.rapid|
C3654136|T201|HIV 1+2 IgG Ab [Presence] in Blood by Rapid immunoassay|
C0482428|T201|Rh immune globulin screen:Imp:Pt:Bld:Nom|
C0482428|T201|Rh immune globulin screen [interpretation]|
C0482428|T201|Rh Ig Scn Bld-Imp|
C0482428|T201|Rh immune globulin screen:Impression/interpretation of study:Point in time:Whole blood:Nominal|
C1555254|T098|Lower Elwha|
C1370055|T201|Gleason Score Spec Ql|
C1370055|T201|Gleason score in Specimen Qualitative|
C1370055|T201|Gleason score:Score:Pt:Specimen:Ord|
C1370055|T201|Gleason score:Score:Point in time:Specimen:Ordinal|
C0362994|T201|Platelet # Bld Auto|
C0362994|T201|Platelets:NCnc:Pt:Bld:Qn:Automated count|
C0362994|T201|Platelets [#/volume] in Blood by Automated count|
C0362994|T201|Platelets:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count|
C0364719|T201|VLDL SerPl-mCnc|
C0364719|T201|Lipoprotein.pre-beta:MCnc:Pt:Ser/Plas:Qn|
C0364719|T201|Lipoprotein.pre-beta [Mass/volume] in Serum or Plasma|
C0364719|T201|Lipoprotein.pre-beta:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0802113|T201|Prostate specific Ag:ACnc:Pt:Ser/Plas:Qn|
C0802113|T201|Prostate specific Ag [Units/volume] in Serum or Plasma|
C0802113|T201|PSA SerPl-aCnc|
C0802113|T201|Prostate specific Antigen:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative|
C1147655|T201|Streptococcus pyogenes Ag [Presence] in Unspecified specimen|
C1147655|T201|Streptococcus pyogenes Ag:ACnc:Pt:XXX:Ord|
C1147655|T201|Streptococcus pyogenes Antigen:Arbitrary Concentration:Point in time:To be specified in another part of the message:Ordinal|
C1147655|T201|S pyo Ag XXX Ql|
C0367888|T201|Reagin Ab:ACnc:Pt:Ser:Ord:VDRL|
C0367888|T201|Reagin Ab [Presence] in Serum by VDRL|
C0367888|T201|VDRL Ser Ql|
C0367888|T201|Reagin Antibody:Arbitrary Concentration:Point in time:Serum:Ordinal:Venereal Disease Research Laboratory|
C0365194|T201|T3RU NFr SerPl|
C0365194|T201|Triiodothyronine resin uptake (T3RU):Number Fraction:Point in time:Serum/Plasma:Quantitative|
C0365194|T201|Triiodothyronine resin uptake (T3RU):NFr:Pt:Ser/Plas:Qn|
C0365194|T201|Triiodothyronine resin uptake (T3RU) in Serum or Plasma|
C0365170|T201|Thyroxine:MCnc:Pt:Ser/Plas:Qn|
C0365170|T201|T4 SerPl-mCnc|
C0365170|T201|Thyroxine:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0365170|T201|Thyroxine (T4) [Mass/volume] in Serum or Plasma|
C0365166|T201|Thyroxine free index:MCnc:Pt:Ser/Plas:Qn|
C0365166|T201|Deprecated Thyroxine free index in Serum or Plasma|
C0365166|T201|Deprecated FTI SerPl-mCnc|
C0365166|T201|Thyroxine free index:Mass Concentration:Point in time:Serum/Plasma:Quantitative|
C0550529|T201|Thyrotropin:ACnc:Pt:Ser/Plas:Qn:Detection limit <= 0.05 mIU/L|
C0550529|T201|TSH SerPl DL<=0.05 mIU/L-aCnc|
C0550529|T201|Thyrotropin [Units/volume] in Serum or Plasma by Detection limit <= 0.05 mIU/L|
C0550529|T201|Thyrotropin:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative:Detection limit <= 0.05 mIU/L|
C0365160|T201|Thyrotropin:ACnc:Pt:Ser/Plas:Qn|
C0365160|T201|Thyrotropin [Units/volume] in Serum or Plasma|
C0365160|T201|TSH SerPl-aCnc|
C0365160|T201|Thyrotropin:Arbitrary Concentration:Point in time:Serum/Plasma:Quantitative|
C1954396|T201|Annotation comment Imp|
C1954396|T201|Annotation comment:Imp:Pt:{system}:Nar|
C1954396|T201|Annotation comment:Impression/interpretation of study:Point in time:{system}:Narrative|
C1954396|T201|Annotation comment [Interpretation] Narrative|
C0801360|T201|Morphology Bld-Imp|
C0801360|T201|Morphology:Imp:Pt:Bld:Nar|
C0801360|T201|Morphology:Impression/interpretation of study:Point in time:Whole blood:Narrative|
C0801360|T201|Morphology [Interpretation] in Blood Narrative|
C0945731|T201|Diagnosis|
C0945731|T201|Dx|
C0945731|T201|Diagnosis:Imp:Pt:^Patient:Nom|
C0945731|T201|Diagnosis:Impression/interpretation of study:Point in time:^Patient:Nominal|
C0551568|T201|General health Reported|
C0551568|T201|General health:Find:Pt:^Patient:Nom:Reported|
C0551568|T201|General health - Reported|
C0551568|T201|General health:Finding:Point in time:^Patient:Nominal:Reported|
C1954395|T201|Information source|
C1954395|T201|Source of info|
C1954395|T201|Information source:Type:Pt:{system}:Nom|
C1954395|T201|Information source:Type:Point in time:{system}:Nominal|
C1316462|T201|Status {Dx}|
C1316462|T201|Status:Class:Pt:{Diagnosis}:Nom|
C1316462|T201|Status [Class] {Diagnosis}|
C1316462|T201|Status:Class:Point in time:{Diagnosis}:Nominal|