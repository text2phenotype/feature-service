C0412621|Computed Tomography (CT) of Liver
C0882012|Multisection:Finding:Point in time:Liver:Narrative:Computerized Tomography
C0807679|Radiology studies
C0411971|Diagnostic radiography of soft tissues
C1962945|Radiographic imaging procedure
C1860232|X-RAY SENSITIVITY
C0202565|GENERAL RADIOLOGY PROCEDURES, TECHNIQUES AND SERVICES
C0043299|Diagnostic radiologic examination
C0918141|Magnetic resonance angiography, head; without contrast material(s)
C0918143|Magnetic resonance angiography, head; without contrast material(s), followed by contrast material(s) and further sequences
C0039985|Plain chest X-ray
C0438647|Radiology/physics in medicine 	
C3668860|Radiologic examination of the Lower Extremities
C3668861|Radiologic examination of the Head and Neck
C3668859|Radiologic examination of the Gastrointestinal Tract
C3668858|Radiologic examination of the Upper Extremities
C2729424|Positron emission tomography (pet) or pet/computed tomography (ct) to inform the initial treatment strategy of tumors that are biopsy proven or strongly suspected of being cancerous based on other diagnostic testing
C2711860|Imaging of liver
C0203765|Liver and spleen imaging
C2711446|Imaging of liver abnormal
C0495790|Abnormal findings diagnostic imaging of liver+biliary tract
C0203758|Radioisotope function study of liver
C0203759|Isotope static scan liver	
C0011923|Diagnostic Imaging
C0203761|Liver imaging with vascular flow
C0203767|Liver and spleen imaging with vascular flow
C0361417|Liver and spleen imaging agents and kits
C0412694|Magnetic Resonance Imaging (MRI) of Liver
C1644183|Radionuclide liver and spleen study
C2314954|MRI of liver with contrast
C2317182|MRI of liver and spleen
C0589338|Dynamic non-imaging isotope study: liver
C2315791|MRI of liver and biliary tract with contrast
C2318037|MRI of liver without contrast
C2584955|MRI guided ablation of liver
C4039879|Imaging guided percutaneous fine needle aspiration biopsy of liver
C2584862|MRI guided focused ultrasound ablation of liver
C2711639|MRI of heart and liver for assessment of cardiac and hepatic iron load
C3880151|Diagnostic imaging table, multi-purpose
C3881113|Diagnostic imaging chair, multi-purpose	
C0043299|Diagnostic radiologic examination
C2317166|Computed tomography of liver with contrast (procedure)
C2317166|Computed tomography (CT) of liver with contrast
C2317166|CT scan of liver with contrast
C2317166|computed tomography of liver with contrast
C2317166|CT of liver with contrast
C2317407|Ablation of lesion of liver using computed tomography (CT) guidance
C2317407|Ablation of lesion of liver using computed tomography guidance (procedure)
C2317407|Ablation of lesion of liver using computed tomography guidance
C2317407|CT guided ablation of lesion of liver
C2315699|Computed tomography of liver and portal vein (procedure)
C2315699|Computed tomography (CT) of liver and portal vein
C2315699|CT of liver and portal vein
C2315699|Computed tomography of liver and portal vein
C2585273|Computed tomography dual phase study of liver (procedure)
C2585273|Computed tomography dual phase study of liver
C2585273|CT dual phase study of liver
C2585560|Computed tomography triple phase study of liver (procedure)
C2585560|Computed tomography triple phase study of liver
C2585560|CT triple phase study of liver
C2321544|computed tomography of liver first without, then with contrast
C2321544|CT scan of liver first without, then with contrast
C2321544|computed tomography of liver first without, then with contrast (procedure)
C0412621|CT of liver (procedure)
C0412621|Computed tomography of liver (procedure)
C0412621|Computed tomography of liver
C0412621|abdominal computed tomography liver
C0412621|Computed Tomography (CT) of Liver
C0412621|CT scan of liver
C0412621|CT of liver
C0412621|CT scan of liver (procedure)
C0412621|Computerised tomogram liver
C0412621|CT scan liver
C0412621|Computerized tomogram liver
C0412621|CT scan;liver
C0412621|CT scan of the liver
C2733010|Single photon emission computed tomography with computed tomography of haemangioma of liver
C2733010|Single photon emission computed tomography with computed tomography of hemangioma of liver (procedure)
C2733010|Single photon emission computed tomography with computed tomography of hemangioma of liver
C2733442|Single photon emission computed tomography with computed tomography of liver and spleen
C2733442|Single photon emission computed tomography with computed tomography of liver and spleen (procedure)
C2123630|abdominal CT liver nonspecific abnormality
C2123630|CT of abdomen nonspecific abnormality of liver
C2123630|computed tomography of abdomen: appearance of nonspecific abnormality of liver
C2123630|computed tomography of abdomen: appearance of nonspecific abnormality of liver (procedure)
C2220596|abdominal computed tomography liver mass lesion
C2220596|CT scan of liver: mass lesion
C2220596|abdominal CT liver mass lesion
C2220596|CT scan of liver mass lesion
C2220596|CT scan of liver: mass lesion (procedure)
C2220584|CT of abdomen liver cyst
C2220584|abdominal CT liver cyst
C2220584|computed tomography of abdomen: liver cyst
C2220584|computed tomography of abdomen: liver cyst (procedure)
C2220588|CT of abdomen diffuse enlargement of liver
C2220588|computed tomography of abdomen: diffuse enlargement of liver
C2220588|computed tomography of abdomen: diffuse enlargement of liver (procedure)
C2220590|CT of abdomen focal enlargement of liver
C2220590|computed tomography of abdomen: focal enlargement of liver (procedure)
C2220590|computed tomography of abdomen: focal enlargement of liver
C2220583|CT of abdomen calcification of liver
C2220583|computed tomography of abdomen: calcification of liver (procedure)
C2220583|computed tomography of abdomen: calcification of liver
C2220587|liver density
C2220587|abdominal CT liver density (HU)
C2220587|CT of abdomen liver density (HU)
C2220587|computed tomography of abdomen: liver density (HU) (procedure)
C2220587|computed tomography of abdomen: liver density (HU)
C2021976|abdominal computed tomography scan liver fibrotic changes
C2021976|abdominal CT fibrotic changes in liver
C2021976|CT of abdomen fibrotic changes in liver
C2021976|computed tomography of abdomen: fibrotic changes in liver (procedure)
C2021976|computed tomography of abdomen: fibrotic changes in liver
C2021977|abdominal CT liver regenerating nodules
C2021977|CT of abdomen regenerating nodules of liver
C2021977|computed tomography of abdomen: regenerating nodules of liver
C2021977|computed tomography of abdomen: regenerating nodules of liver (procedure)
C2021978|CT of abdomen shrunken liver
C2021978|abdominal CT shrunken liver
C2021978|computed tomography of abdomen: shrunken liver
C2021978|computed tomography of abdomen: shrunken liver (procedure)
C2321546|computed tomography of liver without contrast
C2321546|CT scan of liver without contrast
C2321546|computed tomography of liver without contrast (procedure)
C3697202|Positron emission tomography with computed tomography of liver using yttrium 90 microspheres
C3697202|Positron emission tomography with computed tomography of liver using yttrium 90 microspheres (procedure)
C0412627|CT arterioportography (procedure)
C0412627|Computed tomography arterioportography (procedure)
C0412627|Computed tomography arterioportography
C0412627|CT arterioportography
C1636186|CT and drainage of liver
C1636186|Computed tomography and drainage of liver (procedure)
C1636186|Computed tomography and drainage of liver
C1640379|CT and aspiration of liver
C1640379|Computed tomography and aspiration of liver (procedure)
C1640379|Computed tomography and aspiration of liver
C1628488|CT and biopsy of liver
C1628488|Computed tomography and biopsy of liver (procedure)
C1628488|Computed tomography and biopsy of liver
C0882012|Liver CT
C0882012|Multisection:Finding:Point in time:Liver:Narrative:Computerized Tomography
C0882012|Multisection:Find:Pt:Abdomen>Liver:Doc:CT
C0882012|Multisection:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C0807679|RAD
C0807679|Radiology
C0807679|Radiology studies
C0807679|Radiology Procedures
C0942215|TO-Bl MRI
C0942215|Thoracic outlet - bilateral MRI
C0942215|Multisection:Finding:Point in time:Thoracic outlet.bilateral:Document:MRI
C0942215|Multisection:Find:Pt:Thoracic outlet.bilateral:Doc:MRI
C0942230|Lower extremity joint - right MRI
C0942230|LE.joint-R MRI
C0942230|Multisection:Finding:Point in time:Lower extremity.joint.right:Document:MRI
C0942230|Multisection:Find:Pt:Lower extremity.joint.right:Doc:MRI
C0945328|Hand-Bl MRI
C0945328|Hand - bilateral MRI
C0945328|Multisection:Finding:Point in time:Hand.bilateral:Document:MRI
C0945328|Multisection:Find:Pt:Hand.bilateral:Doc:MRI
C0942245|Hand - left MRI
C0942245|Hand-L MRI
C0942245|Multisection:Find:Pt:Hand.left:Doc:MRI
C0942245|Multisection:Finding:Point in time:Hand.left:Document:MRI
C2709261|Deprecated Multisection:Finding:Point in time:Thigh.left:Narrative:MRI
C2709261|Multisection:Find:Pt:Thigh.left:Nar:MRI
C2709261|Deprecated Thigh Left MRI Multisection
C2709261|Deprecated Thigh-L MRI
C2709261|Multisection:Finding:Point in time:Thigh.left:Narrative:MRI
C0942274|Wrist - left US
C0942274|Wrist-L US
C0942274|Multisection:Find:Pt:Wrist.left:Doc:US
C0942274|Multisection:Finding:Point in time:Wrist.left:Document:Ultrasound
C0942282|Breast - left Mammogram limited
C0942282|Brst-L Mam Ltd
C0942282|Views limited:Finding:Point in time:Breast.left:Document:Mam
C0942282|Views limited:Find:Pt:Breast.left:Doc:Mam
C0942284|Breast - right Mammogram limited
C0942284|Brst-R Mam Ltd
C0942284|Views limited:Find:Pt:Breast.right:Doc:Mam
C0942284|Views limited:Finding:Point in time:Breast.right:Document:Mam
C0945334|Vein-Bl XRA Atherect guid W contr IV
C0945334|Fluoroscopic angiogram Guidance for atherectomy of Vein - bilateral-- W contrast IV
C0945334|Guidance for atherectomy^W contrast IV:Find:Pt:Vein.bilateral:Doc:XR.fluor.angio
C0945334|Guidance for atherectomy^W contrast Intravenous:Finding:Point in time:Vein.bilateral:Document:XR.fluor.angio
C0942293|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - left
C0942293|Cent v-L XRA LT per cath plac guid
C0942293|Guidance for placement of longterm peripheral catheter:Find:Pt:Central vein.left:Doc:XR.fluor.angio
C0942293|Guidance for placement of longterm peripheral catheter:Finding:Point in time:Central vein.left:Document:XR.fluor.angio
C0942355|Tibl a-R XRA Angpsty W contr IA
C0942355|Tibial artery - right Fluoroscopic angiogram Angioplasty W contrast IA
C0942355|Angioplasty^W contrast IA:Find:Pt:Tibial artery.right:Doc:XR.fluor.angio
C0942355|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibial artery.right:Document:XR.fluor.angio
C0882073|US Guidance for repair of Pseudoaneurysm/AV fistula
C0882073|PA/AV fistula US Repair guid
C0882073|Guidance for repair:Find:Pt:Pseudoaneurysm/AV fistula:Doc:US
C0882073|Guidance for repair:Finding:Point in time:Pseudoaneurysm/AV fistula:Document:Ultrasound
C0882156|Fluoroscopy Guidance for replacement of percutaneous gastrostomy in Stomach
C0882156|Stom Flr Replac of PEG guid
C0882156|Guidance for replacement of percutaneous gastrostomy:Find:Pt:Stomach:Doc:XR.fluor
C0882156|Guidance for replacement of percutaneous gastrostomy:Finding:Point in time:Stomach:Document:XR.fluor
C0882201|Multisection:Finding:Point in time:To be specified in another part of the message:Narrative:COMPUTERIZED TOMOGRAPHY
C0882201|XXX CT
C0882201|Unspecified body region CT
C0882201|Multisection:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882201|Multisection:Find:Pt:XXX:Doc:CT
C0942114|Foot - bilateral X-ray standing
C0942114|Ft-Bl XR stand
C0942114|Views^standing:Finding:Point in time:Foot.bilateral:Document:XR
C0942114|Views^standing:Find:Pt:Foot.bilateral:Doc:XR
C0945310|Upper extremity - bilateral X-ray
C0945310|UE-Bl XR
C0945310|Views:Find:Pt:Upper extremity.bilateral:Doc:XR
C0945310|Views:Finding:Point in time:Upper extremity.bilateral:Document:XR
C0942139|Deprecated Views:Finding:Point in time:Femur.right:Narrative:XR.DEXA
C0942139|Views:Find:Pt:Femur.right:Nar:XR.DEXA
C0942139|Deprecated Femur-R DEXA
C0942139|Views:Finding:Point in time:Femur.right:Narrative:XR.DEXA
C0942139|Deprecated Femur- right DEXA Bone density
C0882519|Thoracic outlet MRI WO and W contrast IV
C0882519|Multisection^WO & W contrast IV:Find:Pt:Thoracic outlet:Doc:MRI
C0882519|TO MRI WO+W contr IV
C0882519|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thoracic outlet:Document:MRI
C0881829|Deprecated Brain RI
C0881829|Views^W 99m Tc DISIDA or MIBIDA:Find:Pt:Brain:Nar:Radnuc
C0881829|Deprecated Views^W 99m Tc DISIDA or MIBIDA
C0881829|Views^W 99m Tc DISIDA or MIBIDA:Finding:Point in time:Brain:Narrative:Radnuc
C0881840|Brst Mam Dx
C0881840|Breast Mammogram diagnostic
C0881840|Views diagnostic:Find:Pt:Breast:Doc:Mam
C0881840|Views diagnostic:Finding:Point in time:Breast:Document:Mam
C0881903|Esophagus Fluoroscopy W contrast PO
C0881903|Esoph Flr W contr PO
C0881903|Views^W contrast PO:Find:Pt:Esophagus:Doc:XR.fluor
C0881903|Views^W contrast Oral:Finding:Point in time:Esophagus:Document:XR.fluor
C0881928|Foot MRI
C0881928|Ft MRI
C0881928|Multisection:Find:Pt:Foot:Doc:MRI
C0881928|Multisection:Finding:Point in time:Foot:Document:MRI
C0881929|Ft XR stand
C0881929|Foot X-ray standing
C0881929|Views^standing:Find:Pt:Foot:Doc:XR
C0881929|Views^standing:Finding:Point in time:Foot:Document:XR
C0882534|Fluoroscopic angiogram Guidance for placement of stent in Vein
C0882534|Vein XRA Stent plac guid
C0882534|Guidance for placement of stent:Finding:Point in time:Vein:Document:XR.fluor.angio
C0882534|Guidance for placement of stent:Find:Pt:Vein:Doc:XR.fluor.angio
C0881977|Deprecated
C0881977|Multisection:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:Ultrasound
C0881977|Multisection:Find:Pt:Kidney.bilateral+Collecting system:Nar:US
C0881977|Deprecated Kidney - bilateral and Collecting system US
C0881981|Guidance for exchange of percutaneous nephrostomy tube^W contrast:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C0881981|Kdny-Bl Flr PNT exchange guid W contr
C0881981|Fluoroscopy Guidance for exchange of percutaneous nephrostomy tube of Kidney - bilateral-- W contrast
C0881981|Guidance for exchange of percutaneous nephrostomy tube^W contrast:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C1114528|T+L-spine XR Scoli AP 1V
C1114528|View scoliosis AP:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1114528|View scoliosis AP:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1114528|Spine Thoracic and Lumbar X-ray scoliosis AP
C1114541|C-spine XR AP V1 port
C1114541|View AP portable:Find:Pt:Spine.cervical:Doc:XR
C1114541|View AP portable:Finding:Point in time:Spine.cervical:Document:XR
C1114541|Cervical spine X-ray AP portable single view
C1114558|Views portable:Finding:Point in time:Chest:Narrative:XR
C1114558|Chest X-ray portable
C1114558|Chest XR port
C1114558|Views portable:Find:Pt:Chest:Doc:XR
C1114558|Views portable:Finding:Point in time:Chest:Document:XR
C1114596|Views:Finding:Point in time:Patella:Narrative:XR
C1114596|Patella XR
C1114596|Patella X-ray
C1114596|Views:Find:Pt:Patella:Doc:XR
C1114596|Views:Finding:Point in time:Patella:Document:XR
C1114622|Head+Neck a-Bl XRA W contr IA
C1114622|Head artery - bilateral and Neck artery - bilateral Fluoroscopic angiogram W contrast IA
C1114622|Views^W contrast Intra-arterial:Finding:Point in time:Head artery.bilateral+Neck artery.bilateral:Document:XR.fluor.angio
C1114622|Views^W contrast IA:Find:Pt:Head artery.bilateral+Neck artery.bilateral:Doc:XR.fluor.angio
C1114687|BD+PDs Flr Cath guid W contr retro
C1114687|Fluoroscopy Guidance for catheterization of Biliary ducts and Pancreatic duct-- W contrast retrograde
C1114687|Guidance for catheterization^W contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1114687|Guidance for catheterization^W contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1543862|Bone Scan W Sm-153 IV
C1543862|Bone RI W Sm-153 IV
C1543862|Views^W Sm-153 Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543862|Views^W Sm-153 IV:Find:Pt:Bone:Doc:Radnuc
C1543881|Kidney - bilateral SPECT W Tc-99m Mertiatide IV
C1543881|Multisection^W Tc-99m Mertiatide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc.SPECT
C1543881|Multisection^W Tc-99m Mertiatide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc.SPECT
C1543881|Kdny-Bl SPECT W Tc99mMAG3 IV
C1543897|RI Delayed W Ga-67 IV
C1543897|Views delayed^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543897|Views delayed^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543897|Scan delayed W Ga-67 IV
C1543961|Lung RI V+EQ+WO W RNC IH SB
C1543961|Views ventilation & equilibrium & washout^W radionuclide IH single breath:Find:Pt:Lung:Doc:Radnuc
C1543961|Views ventilation & equilibrium & washout^W radionuclide Inhalation single breath:Finding:Point in time:Lung:Document:Radnuc
C1543961|Lung Scan ventilation and equilibrium and washout W radionuclide IH single breath
C1543498|Lower extremity vessels - bilateral US.doppler
C1543498|Multisection:Find:Pt:Lower extremity vessels.bilateral:Doc:US.doppler
C1543498|Multisection:Finding:Point in time:Lower extremity vessels.bilateral:Document:Ultrasound.doppler
C1543498|LE ves-Bl DOP
C1543571|Extr ves-Bl DOP
C1543571|Extremity vessels - bilateral US.doppler
C1543571|Multisection:Find:Pt:Extremity vessels.bilateral:Doc:US.doppler
C1543571|Multisection:Finding:Point in time:Extremity vessels.bilateral:Document:Ultrasound.doppler
C1526357|Skeletal system DXA Bone density
C1526357|Skeletal DXA BDM
C1526357|Bone density:Find:Pt:Skeletal system:Doc:XR.DXA
C1526357|Bone density:Finding:Point in time:Skeletal system:Document:XR.DXA
C1543185|Ribs XR Ant+Lat
C1543185|Ribs X-ray anterior and lateral
C1543185|Views anterior & lateral:Find:Pt:Ribs:Doc:XR
C1543185|Views anterior & lateral:Finding:Point in time:Ribs:Document:XR
C1543264|Deprecated Gastrointestine upper Fluoroscopy W contrast retrograde PR
C1543264|View^W contrast retrograde Rectal:Finding:Point in time:Gastrointestine.upper:Narrative:XR.fluor
C1543264|Deprecated UGI Flr W contr retro PR
C1543264|View^W contrast retrograde PR:Find:Pt:Gastrointestine.upper:Nar:XR.fluor
C1543687|Artery Scan W Tc-99m DTPA IA
C1543687|Artery RI W Tc99mDTPA IA
C1543687|Views^W Tc-99m DTPA Intra-arterial:Finding:Point in time:To be specified in another part of the message artery:Document:Radnuc
C1543687|Views^W Tc-99m DTPA IA:Find:Pt:XXX artery:Doc:Radnuc
C1543695|Brain Scan static
C1543695|Brain RI Static W RNC IV
C1543695|Views static^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc
C1543695|Views static^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1524267|Ft-R XR Tarsal
C1524267|Foot - right X-ray tarsal
C1524267|Views tarsal:Find:Pt:Foot.right:Doc:XR
C1524267|Views tarsal:Finding:Point in time:Foot.right:Document:XR
C1526755|Aorta+Fem a-R XRA Runoff W contr IA
C1526755|Aorta and Femoral artery - right Fluoroscopic angiogram runoff W contrast IA
C1526755|Views runoff^W contrast IA:Find:Pt:Aorta+Femoral artery.right:Doc:XR.fluor.angio
C1526755|Views runoff^W contrast Intra-arterial:Finding:Point in time:Aorta+Femoral artery.right:Document:XR.fluor.angio
C1526769|Lymph-R Flr W contr IL
C1526769|Lymphatics - right Fluoroscopy W contrast intra lymphatic
C1526769|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.right:Doc:XR.fluor
C1526769|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.right:Document:XR.fluor
C1526776|Brst implant-R Mam
C1526776|Breast implant - right Mammogram
C1526776|Views:Finding:Point in time:Breast implant.right:Document:Mam
C1526776|Views:Find:Pt:Breast implant.right:Doc:Mam
C1543415|Ankle-Bl XR AP+Lat stand
C1543415|Ankle - bilateral X-ray AP and lateral standing
C1543415|Views AP & lateral^standing:Finding:Point in time:Ankle.bilateral:Document:XR
C1543415|Views AP & lateral^standing:Find:Pt:Ankle.bilateral:Doc:XR
C1524431|Larynx X-ray tomograph
C1524431|Larynx XRTomo
C1524431|Multisection:Find:Pt:Larynx:Doc:XR.tomo
C1524431|Multisection:Finding:Point in time:Larynx:Document:XR.tomo
C1524182|L-spine XRTomo
C1524182|Multisection:Finding:Point in time:Spine.lumbar:Document:XR.tomo
C1524182|Multisection:Find:Pt:Spine.lumbar:Doc:XR.tomo
C1524182|Lumbar spine X-ray tomograph
C1524192|Upper extremity veins MRI angiogram
C1524192|UE vv MRI.Angio
C1524192|Multisection:Finding:Point in time:Upper extremity veins:Document:MRI.angio
C1524192|Multisection:Find:Pt:Upper extremity veins:Doc:MRI.angio
C1524823|Brst-L MRI WO contr
C1524823|Breast - left MRI WO contrast
C1524823|Multisection^WO contrast:Find:Pt:Breast.left:Doc:MRI
C1524823|Multisection^WO contrast:Finding:Point in time:Breast.left:Document:MRI
C1524843|Upper extremity - right CT WO contrast
C1524843|UE-R CT WO contr
C1524843|Multisection^WO contrast:Find:Pt:Upper extremity.right:Doc:CT
C1524843|Multisection^WO contrast:Finding:Point in time:Upper extremity.right:Document:Computerized Tomography
C1525104|Mastoid X-ray tomograph
C1525104|Mastoid XRTomo
C1525104|Multisection:Find:Pt:Mastoid:Doc:XR.tomo
C1525104|Multisection:Finding:Point in time:Mastoid:Document:XR.tomo
C1524445|Extr CT Ltd
C1524445|Extremity CT limited
C1524445|Multisection limited:Find:Pt:Extremity:Doc:CT
C1524445|Multisection limited:Finding:Point in time:Extremity:Document:Computerized Tomography
C1524448|Lower Extremity Joint MRI limited
C1524448|LE.joint MRI Ltd
C1524448|Multisection limited:Finding:Point in time:Lower extremity.joint:Document:MRI
C1524448|Multisection limited:Find:Pt:Lower extremity.joint:Doc:MRI
C1525220|Multisection^WO & W contrast IV:Find:Pt:Abdominal veins:Doc:MRI.angio
C1525220|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdominal veins:Document:MRI.angio
C1525220|Abdominal veins MRI angiogram WO and W contrast IV
C1525220|Abd vv MRI.Angio WO+W contr IV
C1525222|Multisection^WO & W contrast IV:Find:Pt:Chest veins:Doc:MRI.angio
C1525222|Chest veins MRI angiogram WO and W contrast IV
C1525222|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest veins:Document:MRI.angio
C1525222|Chest vv MRI.Angio WO+W contr IV
C1525224|Multisection^WO & W contrast IV:Find:Pt:Lower extremity veins.right:Doc:MRI.angio
C1525224|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity veins.right:Document:MRI.angio
C1525224|Lower extremity veins - right MRI angiogram WO and W contrast IV
C1525224|LE vv-R MRI.Angio WO+W contr IV
C1525231|Multisection^WO & W contrast IV:Find:Pt:Head vessels:Doc:MRI.angio
C1525231|Head vessels MRI angiogram WO and W contrast IV
C1525231|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head vessels:Document:MRI.angio
C1525231|Head ves MRI.Angio WO+W contr IV
C1525328|Abd XR R-Lat
C1525328|Abdomen X-ray right lateral
C1525328|View R-lateral:Find:Pt:Abdomen:Doc:XR
C1525328|View R-lateral:Finding:Point in time:Abdomen:Document:XR
C1524684|Breast - bilateral Mammogram roll
C1524684|Brst-Bl Mam Roll
C1524684|Views roll:Finding:Point in time:Breast.bilateral:Document:Mam
C1524684|Views roll:Find:Pt:Breast.bilateral:Doc:Mam
C1525461|Should-L XR Transthoracic
C1525461|Shoulder - left X-ray transthoracic
C1525461|View transthoracic:Find:Pt:Shoulder.left:Doc:XR
C1525461|View transthoracic:Finding:Point in time:Shoulder.left:Document:XR
C1525463|Breast Mammogram true lateral
C1525463|Brst Mam True Lat
C1525463|View true lateral:Find:Pt:Breast:Doc:Mam
C1525463|View true lateral:Finding:Point in time:Breast:Document:Mam
C1524220|Wrist - bilateral X-ray ulnar variance
C1524220|Wrist-Bl XR Ulnar Variance
C1524220|View ulnar variance:Find:Pt:Wrist.bilateral:Doc:XR
C1524220|View ulnar variance:Finding:Point in time:Wrist.bilateral:Document:XR
C1525498|Hip-L XR AP+Lat Xtable
C1525498|Hip - left X-ray AP and lateral crosstable
C1525498|Views AP & lateral crosstable:Finding:Point in time:Hip.left:Document:XR
C1525498|Views AP & lateral crosstable:Find:Pt:Hip.left:Doc:XR
C1524246|C-spine XR AP+Obl+Lat W FE
C1524246|Views AP & oblique & lateral^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C1524246|Views AP & oblique & lateral^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C1524246|Cervical spine X-ray AP and oblique and lateral W flexion and W extension
C1525550|Unspecified body region Fluoroscopy portable
C1525550|XXX Flr port
C1525550|Views portable:Find:Pt:XXX:Doc:XR.fluor
C1525550|Views portable:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1525554|Knee XR Obl+Sunrise+Tunnel
C1525554|Knee X-ray oblique and Sunrise and tunnel
C1525554|Views oblique & Sunrise & tunnel:Finding:Point in time:Knee:Document:XR
C1525554|Views oblique & Sunrise & tunnel:Find:Pt:Knee:Doc:XR
C1525586|Views^W contrast Intrasynovial:Finding:Point in time:Sacroiliac joint.bilateral:Document:XR.fluor
C1525586|Views^W contrast IS:Find:Pt:Sacroiliac joint.bilateral:Doc:XR.fluor
C1525586|Sacroiliac joint - bilateral Fluoroscopy W contrast IS
C1525586|SIJ-Bl Flr W contr IS
C1525587|Views^W contrast IS:Find:Pt:Sacroiliac joint.left:Doc:XR.fluor
C1525587|Views^W contrast Intrasynovial:Finding:Point in time:Sacroiliac joint.left:Document:XR.fluor
C1525587|Sacroiliac joint - left Fluoroscopy W contrast IS
C1525587|SIJ-L Flr W contr IS
C1525599|Ankle - left X-ray standing
C1525599|Ankle-L XR stand
C1525599|Views^standing:Finding:Point in time:Ankle.left:Document:XR
C1525599|Views^standing:Find:Pt:Ankle.left:Doc:XR
C1525640|TMJ-L CT W contr IV
C1525640|Temporomandibular joint - left CT W contrast IV
C1525640|Multisection^W contrast Intravenous:Finding:Point in time:Temporomandibular joint.left:Document:Computerized Tomography
C1525640|Multisection^W contrast IV:Find:Pt:Temporomandibular joint.left:Doc:CT
C1525659|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spinal vein:Document:MRI.angio
C1525659|Multisection^WO & W contrast IV:Find:Pt:Spinal vein:Doc:MRI.angio
C1525659|Spinal vein MRI angiogram WO and W contrast IV
C1525659|Spinal v MRI.Angio WO+W contr IV
C1525702|Aorta+Fem a-L XRA Runoff W contr IA
C1525702|Aorta and Femoral artery - left Fluoroscopic angiogram runoff W contrast IA
C1525702|Views runoff^W contrast IA:Find:Pt:Aorta+Femoral artery.left:Doc:XR.fluor.angio
C1525702|Views runoff^W contrast Intra-arterial:Finding:Point in time:Aorta+Femoral artery.left:Document:XR.fluor.angio
C1525727|SMA+IMA XRA W contr IA
C1525727|Superior mesenteric artery and Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C1525727|Views^W contrast Intra-arterial:Finding:Point in time:Superior mesenteric artery+Inferior mesenteric artery:Document:XR.fluor.angio
C1525727|Views^W contrast IA:Find:Pt:Superior mesenteric artery+Inferior mesenteric artery:Doc:XR.fluor.angio
C1525747|Fluoroscopy Guidance for injection of Spine
C1525747|Spine Flr Inj guid
C1525747|Guidance for injection:Finding:Point in time:Spine:Document:XR.fluor
C1525747|Guidance for injection:Find:Pt:Spine:Doc:XR.fluor
C1524699|Wrist-R MRI W contr IV
C1524699|Wrist - right MRI W contrast IV
C1524699|Multisection^W contrast IV:Find:Pt:Wrist.right:Doc:MRI
C1524699|Multisection^W contrast Intravenous:Finding:Point in time:Wrist.right:Document:MRI
C1525785|C+T-spine XR
C1525785|Spine Cervical and Spine Thoracic X-ray
C1525785|Views:Find:Pt:Spine.cervical+Spine.thoracic:Doc:XR
C1525785|Views:Finding:Point in time:Spine.cervical+Spine.thoracic:Document:XR
C1525796|Guidance for biopsy:Find:Pt:Chest>Pleura:Doc:CT
C1525796|Guidance for biopsy:Finding:Point in time:Chest>Pleura:Document:Computerized Tomography
C1525796|CT Guidance for biopsy of Chest Pleura
C1525796|Chest Pleura CT Bx guid
C1525846|Wrist-L XR PA+Lat+Obl
C1525846|Wrist - left X-ray PA and lateral and oblique
C1525846|Views PA & lateral & oblique:Finding:Point in time:Wrist.left:Document:XR
C1525846|Views PA & lateral & oblique:Find:Pt:Wrist.left:Doc:XR
C1525854|Ankle - left X-ray W manual stress
C1525854|Ankle-L XR W Stress
C1525854|Views^W manual stress:Find:Pt:Ankle.left:Doc:XR
C1525854|Views^W manual stress:Finding:Point in time:Ankle.left:Document:XR
C1525869|Deprecated Upper extremity arteries - left Fluoroscopic angiogram W contrast
C1525869|Views^W contrast Intravenous:Finding:Point in time:Upper extremity arteries.left:Narrative:XR.fluor.angio
C1525869|Deprecated UE aa-L XRA W contr IV
C1525869|Views^W contrast IV:Find:Pt:Upper extremity arteries.left:Nar:XR.fluor.angio
C1525806|L-spine ves MRI.Angio W contr IV
C1525806|Lumbar Spine vessels MRI angiogram W contrast IV
C1525806|Multisection^W contrast IV:Find:Pt:Spine.lumbar vessels:Doc:MRI.angio
C1525806|Multisection^W contrast Intravenous:Finding:Point in time:Spine.lumbar vessels:Document:MRI.angio
C1525833|Toe 3rd-L XR
C1525833|Toe third - left X-ray
C1525833|Views:Finding:Point in time:Toe.third.left:Document:XR
C1525833|Views:Find:Pt:Toe.third.left:Doc:XR
C1525962|Wrist - right X-ray ulnar deviation
C1525962|Wrist-R XR Ulnar Deviation
C1525962|View ulnar deviation:Finding:Point in time:Wrist.right:Document:XR
C1525962|View ulnar deviation:Find:Pt:Wrist.right:Doc:XR
C1525900|Wrist-R XR 6V
C1525900|Wrist - right X-ray 6 views
C1525900|Views 6:Finding:Point in time:Wrist.right:Document:XR
C1525900|Views 6:Find:Pt:Wrist.right:Doc:XR
C1526031|Hand-R XR PA+Lat+Obl
C1526031|Hand - right X-ray PA and lateral and oblique
C1526031|Views PA & lateral & oblique:Find:Pt:Hand.right:Doc:XR
C1526031|Views PA & lateral & oblique:Finding:Point in time:Hand.right:Document:XR
C1526034|Views 2:Finding:Point in time:Calcaneus.right:Document:XR
C1526034|Deprecated Calcaneus - right X-ray 2 views
C1526034|Deprecated Heel-R XR 2V
C1526034|Views 2:Find:Pt:Calcaneus.right:Doc:XR
C1526062|Knee - right X-ray AP W manual stress
C1526062|Knee-R XR AP W Stress
C1526062|Views AP^W manual stress:Finding:Point in time:Knee.right:Document:XR
C1526062|Views AP^W manual stress:Find:Pt:Knee.right:Doc:XR
C1524272|Sternum XR 2V
C1524272|Sternum X-ray 2 views
C1524272|Views 2:Find:Pt:Sternum:Doc:XR
C1524272|Views 2:Finding:Point in time:Sternum:Document:XR
C1526211|Ankle aa-R XRA W contr IA
C1526211|Ankle arteries - right Fluoroscopic angiogram W contrast IA
C1526211|Views^W contrast IA:Find:Pt:Ankle arteries.right:Doc:XR.fluor.angio
C1526211|Views^W contrast Intra-arterial:Finding:Point in time:Ankle arteries.right:Document:XR.fluor.angio
C1526219|Extr vv-R XRA W contr IV
C1526219|Extremity veins - right Fluoroscopic angiogram W contrast IV
C1526219|Views^W contrast Intravenous:Finding:Point in time:Extremity veins.right:Document:XR.fluor.angio
C1526219|Views^W contrast IV:Find:Pt:Extremity veins.right:Doc:XR.fluor.angio
C1526221|Carot a+Cerebral a Int-R XRA W contr IA
C1526221|Carotid artery and Cerebral artery internal - right Fluoroscopic angiogram W contrast IA
C1526221|Views^W contrast IA:Find:Pt:Carotid artery+Cerebral artery internal.right:Doc:XR.fluor.angio
C1526221|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Cerebral artery internal.right:Document:XR.fluor.angio
C1526252|Elbow-L XR Radial Head Capitellar
C1526252|Elbow - left X-ray radial head capitellar
C1526252|View radial head capitellar:Find:Pt:Elbow.left:Doc:XR
C1526252|View radial head capitellar:Finding:Point in time:Elbow.left:Document:XR
C1525915|Lower extremity artery - bilateral US
C1525915|LE a-Bl US
C1525915|Multisection:Finding:Point in time:Lower extremity artery.bilateral:Document:Ultrasound
C1525915|Multisection:Find:Pt:Lower extremity artery.bilateral:Doc:US
C1526347|Guidance for superficial biopsy:Find:Pt:Bone:Doc:XR.fluor
C1526347|Fluoroscopy Guidance for superficial biopsy of Bone
C1526347|Guidance for superficial biopsy:Finding:Point in time:Bone:Document:XR.fluor
C1526347|Bone Flr Bx super guid
C1526309|Bones X-ray survey limited for metastasis
C1526309|Bones XR Survey Ltd for Metastasis
C1526309|Views survey limited for metastasis:Find:Pt:Bones:Doc:XR
C1526309|Views survey limited for metastasis:Finding:Point in time:Bones:Document:XR
C1526326|Kidney - right Fluoroscopy W contrast via nephrostomy tube
C1526326|Kidney-R Flr W contr via NT
C1526326|Views^W contrast via nephrostomy tube:Find:Pt:Kidney.right:Doc:XR.fluor
C1526326|Views^W contrast via nephrostomy tube:Finding:Point in time:Kidney.right:Document:XR.fluor
C1524500|Chest MRI W contr IV
C1524500|Chest MRI W contrast IV
C1524500|Multisection^W contrast IV:Find:Pt:Chest:Doc:MRI
C1524500|Multisection^W contrast Intravenous:Finding:Point in time:Chest:Document:MRI
C1524878|Upper arm - left MRI WO contrast
C1524878|Upper arm-L MRI WO contr
C1524878|Multisection^WO contrast:Find:Pt:Upper arm.left:Doc:MRI
C1524878|Multisection^WO contrast:Finding:Point in time:Upper arm.left:Document:MRI
C1524886|SIJ CT WO contr
C1524886|Sacroiliac Joint CT WO contrast
C1524886|Multisection^WO contrast:Find:Pt:Sacroiliac joint:Doc:CT
C1524886|Multisection^WO contrast:Finding:Point in time:Sacroiliac joint:Document:Computerized Tomography
C1524525|Ft-L CT W contr IV
C1524525|Foot - left CT W contrast IV
C1524525|Multisection^W contrast Intravenous:Finding:Point in time:Foot.left:Document:Computerized Tomography
C1524525|Multisection^W contrast IV:Find:Pt:Foot.left:Doc:CT
C1524545|Upper arm-R CT W contr IV
C1524545|Upper arm - right CT W contrast IV
C1524545|Multisection^W contrast IV:Find:Pt:Upper arm.right:Doc:CT
C1524545|Multisection^W contrast Intravenous:Finding:Point in time:Upper arm.right:Document:Computerized Tomography
C1524309|Guidance for biopsy^WO & W contrast Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C1524309|Chest CT Bx guid WO+W contr IV
C1524309|Guidance for biopsy^WO & W contrast IV:Find:Pt:Chest:Doc:CT
C1524309|CT Guidance for biopsy of Chest-- WO and W contrast IV
C1524310|CT Guidance for biopsy of Chest-- WO contrast
C1524310|Chest CT Bx guid WO contr
C1524310|Guidance for biopsy^WO contrast:Finding:Point in time:Chest:Document:Computerized Tomography
C1524310|Guidance for biopsy^WO contrast:Find:Pt:Chest:Doc:CT
C1524131|Chest MRI WO+W contr IV
C1524131|Multisection^WO & W contrast IV:Find:Pt:Chest:Doc:MRI
C1524131|Chest MRI WO and W contrast IV
C1524131|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest:Document:MRI
C1524975|Breast - left Mammogram
C1524975|Brst-L Mam
C1524975|Views:Find:Pt:Breast.left:Doc:Mam
C1524975|Views:Finding:Point in time:Breast.left:Document:Mam
C1525017|Knee - bilateral X-ray 6 views
C1525017|Knee-Bl XR 6V
C1525017|Views 6:Find:Pt:Knee.bilateral:Doc:XR
C1525017|Views 6:Finding:Point in time:Knee.bilateral:Document:XR
C1524752|Upper arm CT WO and W contrast IV
C1524752|Upper arm CT WO+W contr IV
C1524752|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper arm:Document:Computerized Tomography
C1524752|Multisection^WO & W contrast IV:Find:Pt:Upper arm:Doc:CT
C1525044|Pelvis+Hip XR AP+Lat
C1525044|Pelvis and Hip X-ray AP and lateral
C1525044|Views AP & lateral:Find:Pt:Pelvis+Hip:Doc:XR
C1525044|Views AP & lateral:Finding:Point in time:Pelvis+Hip:Document:XR
C1525055|Should-Bl XR AP+Lat
C1525055|Shoulder - bilateral X-ray AP and lateral
C1525055|Views AP & lateral:Find:Pt:Shoulder.bilateral:Doc:XR
C1525055|Views AP & lateral:Finding:Point in time:Shoulder.bilateral:Document:XR
C1524414|Upper arm MRI
C1524414|Multisection:Finding:Point in time:Upper arm:Document:MRI
C1524414|Multisection:Find:Pt:Upper arm:Doc:MRI
C1524783|Sinuses CT WO and W contrast IV
C1524783|Sinuses CT WO+W contr IV
C1524783|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head>Sinuses:Document:Computerized Tomography
C1524783|Multisection^WO & W contrast IV:Find:Pt:Head>Sinuses:Doc:CT
C1525076|C-spine XR Obl
C1525076|Views oblique:Find:Pt:Spine.cervical:Doc:XR
C1525076|Views oblique:Finding:Point in time:Spine.cervical:Document:XR
C1525076|Cervical spine X-ray oblique
C1525081|Hand-L XR PA+Lat
C1525081|Hand - left X-ray PA and lateral
C1525081|Views PA & lateral:Find:Pt:Hand.left:Doc:XR
C1525081|Views PA & lateral:Finding:Point in time:Hand.left:Document:XR
C1830196|Brst-L Mam Bx CN Str Guid
C1830196|Guidance for stereotactic biopsy.core needle:Find:Pt:Breast.left:Doc:Mam
C1830196|Guidance for stereotactic biopsy.core needle:Finding:Point in time:Breast.left:Document:Mam
C1830196|Mammogram Guidance for stereotactic core needle biopsy of Breast - left
C1830215|Multisection^WO & W reduced contrast volume Intravenous:Finding:Point in time:Internal auditory canal:Document:Computerized Tomography
C1830215|IAC CT WO+W red contr vol IV
C1830215|Internal auditory canal CT WO and W reduced contrast volume IV
C1830215|Multisection^WO & W reduced contrast volume IV:Find:Pt:Internal auditory canal:Doc:CT
C1830247|Wrist-L XR GE 3V
C1830247|Wrist - left X-ray GE 3 views
C1830247|Views GE 3:Finding:Point in time:Wrist.left:Document:XR
C1830247|Views GE 3:Find:Pt:Wrist.left:Doc:XR
C1830091|Skull XR GE 3V
C1830091|Skull X-ray GE 3 views
C1830091|Views GE 3:Find:Pt:Skull:Doc:XR
C1830091|Views GE 3:Finding:Point in time:Skull:Document:XR
C1830281|Fluoroscopy Guidance for injection of Sinuses
C1830281|Sinuses Flr Inj guid
C1830281|Guidance for injection:Find:Pt:Sinuses:Doc:XR.fluor
C1830281|Guidance for injection:Finding:Point in time:Sinuses:Document:XR.fluor
C1831070|Hip X-ray during surgery
C1831070|Hip XR in Surg
C1831070|Views^during surgery:Finding:Point in time:Hip:Document:XR
C1831070|Views^during surgery:Find:Pt:Hip:Doc:XR
C1715414|BM RI W Tc99mSC IV
C1715414|Bone marrow Scan W Tc-99m SC IV
C1715414|Views^W Tc-99m SC IV:Find:Pt:Bone marrow:Doc:Radnuc
C1715414|Views^W Tc-99m Subcutaneous Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc
C1715463|Views 1 or 2 limited:Finding:Point in time:Sinuses:Narrative:XR
C1715463|Deprecated Sinuses XR 1V or 2V Ltd
C1715463|Views 1 or 2 limited:Find:Pt:Sinuses:Nar:XR
C1715463|Deprecated Sinuses X-ray 1 or 2 views limited
C1715498|Periph aa-Bl XRA W contr IA
C1715498|Peripheral arteries - bilateral Fluoroscopic angiogram W contrast IA
C1715498|Views^W contrast IA:Find:Pt:Peripheral arteries.bilateral:Doc:XR.fluor.angio
C1715498|Views^W contrast Intra-arterial:Finding:Point in time:Peripheral arteries.bilateral:Document:XR.fluor.angio
C1645315|US Guidance for drainage of Abdomen retroperitoneum
C1645315|Abd.reper US Drain guid
C1645315|Guidance for drainage:Finding:Point in time:Abdomen.retroperitoneum:Document:Ultrasound
C1645315|Guidance for drainage:Find:Pt:Abdomen.retroperitoneum:Doc:US
C1649412|Extremity veins - right US
C1649412|Extr vv-R US
C1649412|Multisection:Find:Pt:Extremity veins.right:Doc:US
C1649412|Multisection:Finding:Point in time:Extremity veins.right:Document:Ultrasound
C1635068|Ankle-L XR AP+Lat stand
C1635068|Ankle - left X-ray AP and lateral standing
C1635068|Views AP & lateral^standing:Find:Pt:Ankle.left:Doc:XR
C1635068|Views AP & lateral^standing:Finding:Point in time:Ankle.left:Document:XR
C1636066|Spine Lumbar X-ray (AP W R-bending and W L-bending and WO bending) and Lateral
C1636066|L-spine XR (AP W+WO R+L-bending)+Lat
C1636066|Views (AP^W R-bending & W L-bending & WO bending) & lateral:Finding:Point in time:Spine.lumbar:Document:XR
C1636066|Views (AP^W R-bending & W L-bending & WO bending) & lateral:Find:Pt:Spine.lumbar:Doc:XR
C1714900|Foot - left X-ray 3 or 4 views
C1714900|Ft-L XR 3V or 4V
C1714900|Views 3 or 4:Find:Pt:Foot.left:Doc:XR
C1714900|Views 3 or 4:Finding:Point in time:Foot.left:Document:XR
C1714959|Abdominal vessels US.doppler limited
C1714959|Abd ves DOP Ltd
C1714959|Multisection limited:Finding:Point in time:Abdominal vessels:Document:Ultrasound.doppler
C1714959|Multisection limited:Find:Pt:Abdominal vessels:Doc:US.doppler
C1714498|Renal ves RI Flow W Tc99mDTPA IV
C1714498|Renal vessels Scan flow W Tc-99m DTPA IV
C1714498|Views flow^W Tc-99m DTPA IV:Find:Pt:Renal vessels:Doc:Radnuc
C1714498|Views flow^W Tc-99m DTPA Intravenous:Finding:Point in time:Renal vessels:Document:Radnuc
C1715094|Kidney - bilateral CT W contrast IV
C1715094|Multisection^W contrast IV:Find:Pt:Kidney.bilateral:Doc:CT
C1715094|Multisection^W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:Computerized Tomography
C1715094|Kdny-Bl CT W contr IV
C1717275|Extremity vessels US.doppler
C1717275|Extr ves DOP
C1717275|Multisection:Find:Pt:Extremity vessels:Doc:US.doppler
C1717275|Multisection:Finding:Point in time:Extremity vessels:Document:Ultrasound.doppler
C1715108|Iliac a XRA W contr IA
C1715108|Iliac artery Fluoroscopic angiogram W contrast IA
C1715108|Views^W contrast Intra-arterial:Finding:Point in time:Iliac artery:Document:XR.fluor.angio
C1715108|Views^W contrast IA:Find:Pt:Iliac artery:Doc:XR.fluor.angio
C1715123|US Guidance for biopsy of Superficial lymph node
C1715123|Superf LN US Bx guid
C1715123|Guidance for biopsy:Finding:Point in time:Superficial lymph node:Document:Ultrasound
C1715123|Guidance for biopsy:Find:Pt:Superficial lymph node:Doc:US
C1625792|Fluoroscopy Guidance for percutaneous drainage of abscess of Chest
C1625792|Chest Flr PC Abscess Drain guid
C1625792|Guidance for percutaneous drainage of abscess:Find:Pt:Chest:Doc:XR.fluor
C1625792|Guidance for percutaneous drainage of abscess:Finding:Point in time:Chest:Document:XR.fluor
C1637283|Neck X-ray magnification
C1637283|Neck XR Mag
C1637283|View magnification:Finding:Point in time:Neck:Document:XR
C1637283|View magnification:Find:Pt:Neck:Doc:XR
C1644147|UGI+SB Flr W Air contr PO
C1644147|Upper Gastrointestine and Small bowel Fluoroscopy W air contrast PO
C1644147|View^W air contrast Oral:Finding:Point in time:Gastrointestine.upper+Small bowel:Document:XR.fluor
C1644147|View^W air contrast PO:Find:Pt:Gastrointestine.upper+Small bowel:Doc:XR.fluor
C1624130|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower leg.bilateral:Document:MRI
C1624130|Lower leg-Bl MRI WO+W contr IV
C1624130|Multisection^WO & W contrast IV:Find:Pt:Lower leg.bilateral:Doc:MRI
C1624130|Lower leg - bilateral MRI WO and W contrast IV
C1977327|Ankle - bilateral X-ray GE 6 views
C1977327|Ankle-Bl XR GE 6V
C1977327|Views GE 6:Find:Pt:Ankle.bilateral:Doc:XR
C1977327|Views GE 6:Finding:Point in time:Ankle.bilateral:Document:XR
C1953966|Unspecified body region MRI limited
C1953966|XXX MRI Ltd
C1953966|Multisection limited:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1953966|Multisection limited:Find:Pt:XXX:Doc:MRI
C1953976|L-spine XR 2V or 3V
C1953976|Views 2 or 3:Finding:Point in time:Spine.lumbar:Document:XR
C1953976|Views 2 or 3:Find:Pt:Spine.lumbar:Doc:XR
C1953976|Lumbar spine X-ray 2 or 3 views
C1953987|Face XR GE 3V
C1953987|Facial bones X-ray GE 3 views
C1953987|Views GE 3:Find:Pt:Facial bones:Doc:XR
C1953987|Views GE 3:Finding:Point in time:Facial bones:Document:XR
C3175182|FR-R Flr Cath guid transcervical
C3175182|Fluoroscopy Guidance for catheterization of Fallopian tube -right-- transcervical
C3175182|Guidance for catheterization^transcervical:Find:Pt:Fallopian tube.right:Doc:XR.fluor
C3175182|Guidance for catheterization^transcervical:Finding:Point in time:Fallopian tube.right:Document:XR.fluor
C3169524|Renal a-R XRA W contr IA
C3169524|Renal artery - right Fluoroscopic angiogram W contrast IA
C3169524|Views^W contrast IA:Find:Pt:Renal artery.right:Doc:XR.fluor.angio
C3169524|Views^W contrast Intra-arterial:Finding:Point in time:Renal artery.right:Document:XR.fluor.angio
C3169580|Fluoroscopic angiogram Guidance for placement of ilio-iliac tube endoprosthesis in Iliac artery - right-- W contrast IA
C3169580|Iliac a-R XRA Ilio tube guid W contr IA
C3169580|Guidance for placement of ilio-iliac tube endoprosthesis^W contrast IA:Find:Pt:Iliac artery.right:Doc:XR.fluor.angio
C3169580|Guidance for placement of ilio-iliac tube endoprosthesis^W contrast Intra-arterial:Finding:Point in time:Iliac artery.right:Document:XR.fluor.angio
C3533564|Fluoroscopic angiogram Guidance for removal of longterm peripheral catheter from Central vein
C3533564|Centl v XRA LT per cath removal guid
C3533564|Guidance for removal of longterm peripheral catheter:Find:Pt:Central vein:Doc:XR.fluor.angio
C3533564|Guidance for removal of longterm peripheral catheter:Finding:Point in time:Central vein:Document:XR.fluor.angio
C3533559|Guidance for intercostal nerve devervation:Finding:Point in time:Spine.thoracic:Document:XR.fluor
C3533559|T-spine Flr ICN DN guid
C3533559|Guidance for intercostal nerve devervation:Find:Pt:Spine.thoracic:Doc:XR.fluor
C3533559|Fluoroscopy Guidance for intercostal nerve devervation of Thoracic spine
C3533479|Extr v-R US Sclerosing agent inj guid
C3533479|Guidance for injection of sclerosing agent:Find:Pt:Extremity vein.right:Doc:US
C3533479|Guidance for injection of sclerosing agent:Finding:Point in time:Extremity vein.right:Document:Ultrasound
C3533479|US Guidance for injection of sclerosing agent of Extremity vein - right
C3262954|Hip XR Danelius Miller
C3262954|Hip XR +Danelius Miller
C3262954|Hip X-ray and Danelius Miller
C3262954|Hip X-ray Danelius Miller
C3262954|Views & Danelius Miller:Finding:Point in time:Hip:Document:XR
C3262954|Views & Danelius Miller:Find:Pt:Hip:Doc:XR
C3262954|View Danelius Miller:Finding:Point in time:Hip:Document:XR
C3262954|View Danelius Miller:Find:Pt:Hip:Doc:XR
C3263010|Breast implant MRI W contrast IV
C3263010|Brst implant MRI W contr IV
C3263010|Multisection^W contrast Intravenous:Finding:Point in time:Breast implant:Document:MRI
C3263010|Multisection^W contrast IV:Find:Pt:Breast implant:Doc:MRI
C3263031|Should-R MRI WO+W contr IS
C3263031|Multisection^WO & W contrast IS:Find:Pt:Shoulder.right:Doc:MRI
C3263031|Shoulder - right MRI WO and W contrast IS
C3263031|Multisection^WO & W contrast Intrasynovial:Finding:Point in time:Shoulder.right:Document:MRI
C3263034|Scrotum and Testicle MRI W contrast IV
C3263034|Scrotum+Test MRI W contr IV
C3263034|Multisection^W contrast Intravenous:Finding:Point in time:Scrotum+Testicle:Document:MRI
C3263034|Multisection^W contrast IV:Find:Pt:Scrotum+Testicle:Doc:MRI
C3263066|Renal ves XRA Atherect W contr
C3263066|Renal vessels Fluoroscopic angiogram Atherectomy W contrast
C3263066|Atherectomy^W contrast:Finding:Point in time:Renal vessels:Document:XR.fluor.angio
C3263066|Atherectomy^W contrast:Find:Pt:Renal vessels:Doc:XR.fluor.angio
C3261477|View 1:Find:Pt:Calcaneus.right:Doc:XR
C3261477|View 1:Finding:Point in time:Calcaneus.right:Document:XR
C3261477|Deprecated Heel-R XR 1V
C3261477|Deprecated Calcaneus - right X-ray Single view
C3261477|Deprecated View 1:Find:Pt:Calcaneus.right:Doc:XR
C3263218|US Guidance for chorionic villus sampling
C3263218|US CVS Guid
C3263218|Guidance for chorionic villus sampling:Finding:Point in time:Placenta:Document:Ultrasound
C3263218|Guidance for chorionic villus sampling:Find:Pt:Placenta:Doc:US
C3262907|Chest vessels CT angiogram WO contrast
C3262907|Multisection^WO contrast:Finding:Point in time:Chest>Vessels:Document:Computerized Tomography.angio
C3262907|Multisection^WO contrast:Find:Pt:Chest>Vessels:Doc:CT.angio
C3262907|Chest Ves CT.Angio WO contr
C3262910|Ankle-Bl CT WO contr
C3262910|Ankle - bilateral CT WO contrast
C3262910|Multisection^WO contrast:Finding:Point in time:Ankle.bilateral:Document:Computerized Tomography
C3262910|Multisection^WO contrast:Find:Pt:Ankle.bilateral:Doc:CT
C3262925|Multisection^W contrast IS:Find:Pt:Ankle.left:Doc:CT
C3262925|Ankle-L CT W contr IS
C3262925|Multisection^W contrast Intrasynovial:Finding:Point in time:Ankle.left:Document:Computerized Tomography
C3262925|Ankle - left CT W contrast IS
C0942184|Breast - bilateral Mammogram screening
C0942184|Brst-Bl Mam Screening
C0942184|Views screening:Find:Pt:Breast.bilateral:Doc:Mam
C0942184|Views screening:Finding:Point in time:Breast.bilateral:Document:Mam
C0942229|LE.joint-L MRI
C0942229|Lower extremity joint - left MRI
C0942229|Multisection:Find:Pt:Lower extremity.joint.left:Doc:MRI
C0942229|Multisection:Finding:Point in time:Lower extremity.joint.left:Document:MRI
C0942248|Internal auditory canal - bilateral X-ray tomograph
C0942248|IAC-Bl XRTomo
C0942248|Multisection:Finding:Point in time:Internal auditory canal.bilateral:Document:XR.tomo
C0942248|Multisection:Find:Pt:Internal auditory canal.bilateral:Doc:XR.tomo
C0942255|Pelvis+Hip-L MRI
C0942255|Pelvis and Hip - left MRI
C0942255|Multisection:Finding:Point in time:Pelvis+Hip.left:Document:MRI
C0942255|Multisection:Find:Pt:Pelvis+Hip.left:Doc:MRI
C0945333|Cent v-R XRA Cath repos W contr IV
C0945333|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - right-- W contrast IV
C0945333|Guidance for reposition of catheter^W contrast IV:Find:Pt:Central vein.right:Doc:XR.fluor.angio
C0945333|Guidance for reposition of catheter^W contrast Intravenous:Finding:Point in time:Central vein.right:Document:XR.fluor.angio
C0942299|Cent v-R XRA Cath plac guid W contr IV
C0942299|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - right-- W contrast IV
C0942299|Guidance for placement of catheter^W contrast Intravenous:Finding:Point in time:Central vein.right:Document:XR.fluor.angio
C0942299|Guidance for placement of catheter^W contrast IV:Find:Pt:Central vein.right:Doc:XR.fluor.angio
C0942340|Knee - right X-ray AP single view standing
C0942340|Knee-R XR AP 1V stand
C0942340|View AP^standing:Finding:Point in time:Knee.right:Document:XR
C0942340|View AP^standing:Find:Pt:Knee.right:Doc:XR
C0942364|Ankle - bilateral X-ray 2 views
C0942364|Ankle-Bl XR 2V
C0942364|Views 2:Find:Pt:Ankle.bilateral:Doc:XR
C0942364|Views 2:Finding:Point in time:Ankle.bilateral:Document:XR
C0882044|Orbit-Bl MRI WO+W contr IV
C0882044|Multisection^WO & W contrast Intravenous:Finding:Point in time:Orbit.bilateral:Document:MRI
C0882044|Multisection^WO & W contrast IV:Find:Pt:Orbit.bilateral:Doc:MRI
C0882044|Orbit - bilateral MRI WO and W contrast IV
C0882145|T-spine Flr W contr IT
C0882145|Views^W contrast Intrathecal:Finding:Point in time:Spine.thoracic:Document:XR.fluor
C0882145|Views^W contrast IT:Find:Pt:Spine.thoracic:Doc:XR.fluor
C0882145|Thoracic spine Fluoroscopy W contrast IT
C0882152|Splenic artery Fluoroscopic angiogram W contrast IA
C0882152|Splenic a XRA W contr IA
C0882152|Views^W contrast IA:Find:Pt:Splenic artery:Doc:XR.fluor.angio
C0882152|Views^W contrast Intra-arterial:Finding:Point in time:Splenic artery:Document:XR.fluor.angio
C0882196|Deprecated Unspecified body region CT 3D
C0882196|Multisection:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography.3D
C0882196|Deprecated XXX CT.3D
C0882196|Multisection:Find:Pt:XXX:Doc:CT.3D
C0882198|XXX CT Asp or Bx guid
C0882198|CT Guidance for aspiration or biopsy of Unspecified body region
C0882198|Guidance for aspiration or biopsy:Find:Pt:XXX:Doc:CT
C0882198|Guidance for aspiration or biopsy:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882223|Zygomatic arch X-ray
C0882223|Zygomatic arch XR
C0882223|Views:Find:Pt:Zygomatic arch:Doc:XR
C0882223|Views:Finding:Point in time:Zygomatic arch:Document:XR
C0942089|Vein-L XRA W contr IV
C0942089|Vein - left Fluoroscopic angiogram W contrast IV
C0942089|Views^W contrast Intravenous:Finding:Point in time:Vein.left:Document:XR.fluor.angio
C0942089|Views^W contrast IV:Find:Pt:Vein.left:Doc:XR.fluor.angio
C0881804|Views AP (KUB & upright) & upright chest:Finding:Point in time:Chest+Abdomen:Narrative:XR
C0881804|Deprecated Chest+Abd XR
C0881804|Views AP (KUB & upright) & upright chest:Find:Pt:Chest+Abdomen:Nar:XR
C0881804|Deprecated Chest and Abdomen Narrative X-ray
C0881808|AV shunt XRA W contr IV
C0881808|AV shunt Fluoroscopic angiogram W contrast IV
C0881808|Views^W contrast IV:Find:Pt:AV shunt:Doc:XR.fluor.angio
C0881808|Views^W contrast Intravenous:Finding:Point in time:AV shunt:Document:XR.fluor.angio
C0881898|Duodenum Flr W contr PO+Hypo Agent NG
C0881898|Duodenum Fluoroscopy W contrast PO and hypotonic agent per ng
C0881898|Views^W contrast PO & hypotonic agent per ng:Find:Pt:Duodenum:Doc:XR.fluor
C0881898|Views^W contrast Oral & hypotonic agent per ng:Finding:Point in time:Duodenum:Document:XR.fluor
C0881910|Periph vv XRA W contr IV
C0881910|Peripheral veins Fluoroscopic angiogram W contrast IV
C0881910|Views^W contrast Intravenous:Finding:Point in time:Peripheral veins.To be specified in another part of the message:Document:XR.fluor.angio
C0881910|Views^W contrast IV:Find:Pt:Peripheral veins.XXX:Doc:XR.fluor.angio
C0881946|Multisection:Find:Pt:Head:Doc:CT.perfusion
C0881946|Multisection:Finding:Point in time:Head:Document:Computerized Tomography.perfusion
C0881946|Head CT perfusion
C0881946|Head CT.perfusion
C0881972|Fluoroscopy Guidance for aspiration of Joint space
C0881972|Guidance for aspiration:Find:Pt:Joint space:Doc:XR.fluor
C0881972|Guidance for aspiration:Finding:Point in time:Joint space:Document:XR.fluor
C0881972|Joint space Flr Asp guid
C0881983|Kidney - bilateral Fluoroscopy Urodynamics
C0881983|Urodynamics:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C0881983|Urodynamics:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C0881983|Kdny-Bl Flr Urodynamics
C0882015|Liver+Diaphragm US
C0882015|Liver and Diaphragm US
C0882015|Multisection:Find:Pt:Liver+Diaphragm:Doc:US
C0882015|Multisection:Finding:Point in time:Liver+Diaphragm:Document:Ultrasound
C1114606|Maxillofacial region CT WO and W contrast IV
C1114606|Maxillofacial CT WO+W contr IV
C1114606|Multisection^WO & W contrast IV:Find:Pt:Head>Maxillofacial region:Doc:CT
C1114606|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1114645|Renal v-Bl XRA W contr IV
C1114645|Renal vein - bilateral Fluoroscopic angiogram W contrast IV
C1114645|Views^W contrast IV:Find:Pt:Renal vein.bilateral:Doc:XR.fluor.angio
C1114645|Views^W contrast Intravenous:Finding:Point in time:Renal vein.bilateral:Document:XR.fluor.angio
C1114427|Chest CT WO+W contr IV
C1114427|Chest CT WO and W contrast IV
C1114427|Multisection^WO & W contrast IV:Find:Pt:Chest:Doc:CT
C1114427|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C1114442|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Pancreas:Doc:CT
C1114442|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C1114442|Pancreas CT WO+W contr IV
C1114442|Pancreas CT WO and W contrast IV
C1114930|US Guidance for placement of catheter in Central vein
C1114930|Centl v US Cath plac guid
C1114930|Guidance for placement of catheter:Find:Pt:Central vein:Doc:US
C1114930|Guidance for placement of catheter:Finding:Point in time:Central vein:Document:Ultrasound
C1543433|Should-L XR AP(w IR+ER)+Y
C1543433|Shoulder - left X-ray AP (W internal rotation and W external rotation) and Y
C1543433|Views AP (W internal rotation & W external rotation) & Y:Finding:Point in time:Shoulder.left:Document:XR
C1543433|Views AP (W internal rotation & W external rotation) & Y:Find:Pt:Shoulder.left:Doc:XR
C1543752|Hrt SPECT PF W ADE+RNC IV
C1543752|Heart SPECT perfusion W adenosine and W radionuclide IV
C1543752|Multisection perfusion^W adenosine & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543752|Multisection perfusion^W adenosine & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543765|Hrt RI PF W Tl-201 IV+Tc99mTF IV
C1543765|Heart Scan perfusion W Tl-201 IV and Tc-99m Tetrofosmin IV
C1543765|Views perfusion^W Tl-201 Intravenous & Tc-99m Tetrofosmin Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543765|Views perfusion^W Tl-201 IV & Tc-99m Tetrofosmin IV:Find:Pt:Heart:Doc:Radnuc
C1543771|Hrt RI PF Rest+W ADE+RNC IV
C1543771|Heart Scan perfusion at rest and W adenosine and W radionuclide IV
C1543771|Views perfusion^at rest & W adenosine & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543771|Views perfusion^at rest & W adenosine & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543774|Hrt RI PF Rest+W DPY+RNC IV
C1543774|Heart Scan perfusion at rest and W dipyridamole and W radionuclide IV
C1543774|Views perfusion^at rest & W dipyridamole & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543774|Views perfusion^at rest & W dipyridamole & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543789|Neck Scan
C1543789|Neck RI W RNC IV
C1543789|Views^W radionuclide Intravenous:Finding:Point in time:Neck:Document:Radnuc
C1543789|Views^W radionuclide IV:Find:Pt:Neck:Doc:Radnuc
C1543864|Bone marrow Scan limited
C1543864|BM RI Ltd W RNC IV
C1543864|Views limited^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc
C1543864|Views limited^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc
C1543868|Bone marrow Scan whole body
C1543868|BM RI WB W RNC IV
C1543868|Views whole body^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc
C1543868|Views whole body^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc
C1543885|Scrotum+Test RI Static W RNC IV
C1543885|Scrotum and Testicle Scan static
C1543885|Views static^W radionuclide IV:Find:Pt:Scrotum+Testicle:Doc:Radnuc
C1543885|Views static^W radionuclide Intravenous:Finding:Point in time:Scrotum+Testicle:Document:Radnuc
C1543891|Heart Scan blood pool
C1543891|Hrt RI BP W RNC IV
C1543891|Views blood pool^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543891|Views blood pool^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543906|Bone RI BP W RNC IV
C1543906|Bone Scan blood pool
C1543906|Views blood pool^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543906|Views blood pool^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543962|RI Mul Areas W In-111 Satmb IV
C1543962|Scan multiple areas W In-111 Satumomab IV
C1543962|Views multiple areas^W In-111 Satumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543962|Views multiple areas^W In-111 Satumomab IV:Find:Pt:^Patient:Doc:Radnuc
C1543152|Extr a-Bl DOP
C1543152|Extremity artery - bilateral US.doppler
C1543152|Multisection:Finding:Point in time:Extremity artery.bilateral:Document:Ultrasound.doppler
C1543152|Multisection:Find:Pt:Extremity artery.bilateral:Doc:US.doppler
C1543567|Ribs upper ant+post-R XR
C1543567|Ribs upper anterior and posterior - right X-ray
C1543567|Views:Find:Pt:Ribs.upper.anterior+posterior.right:Doc:XR
C1543567|Views:Finding:Point in time:Ribs.upper.anterior+posterior.right:Document:XR
C1526352|Bone density:T Score:Point in time:Femur:Quantitative:XR.DXA
C1526352|Femur DXA [T-score] Bone density
C1526352|Femur DXA T-score BDM
C1526352|Bone density:Tscore:Pt:Femur:Qn:XR.DXA
C1543187|Chest Flr AP+Lat
C1543187|Chest Fluoroscopy AP and lateral
C1543187|Views AP & lateral:Finding:Point in time:Chest:Document:XR.fluor
C1543187|Views AP & lateral:Find:Pt:Chest:Doc:XR.fluor
C1542861|Breast FFD mammogram Post Localization
C1542861|Views^post localization:Find:Pt:Breast:Doc:Mam.FFD
C1542861|Brst FFDM p local
C1542861|Views^post localization:Finding:Point in time:Breast:Document:Mam.FFD
C1543698|Brain Scan flow
C1543698|Brain RI Flow W RNC IV
C1543698|Views flow^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1543698|Views flow^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc
C1526760|Hand-R XR Bora
C1526760|Hand - right X-ray Bora
C1526760|View Bora:Find:Pt:Hand.right:Doc:XR
C1526760|View Bora:Finding:Point in time:Hand.right:Document:XR
C1526761|Shoulder - right X-ray Grashey
C1526761|Should-R XR Grashey
C1526761|View Grashey:Find:Pt:Shoulder.right:Doc:XR
C1526761|View Grashey:Finding:Point in time:Shoulder.right:Document:XR
C1526766|Great toe-R XR stand
C1526766|Great toe - right X-ray standing
C1526766|Views^standing:Finding:Point in time:Great toe.right:Document:XR
C1526766|Views^standing:Find:Pt:Great toe.right:Doc:XR
C1542970|SPECT for Inf W Ga-67 IV
C1542970|Multisection for infection^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1542970|Multisection for infection^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1542970|SPECT for infection W Ga-67 IV
C1542972|RI for Inf W Ga-67 IV
C1542972|Views for infection^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1542972|Views for infection^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542972|Scan for infection W Ga-67 IV
C1526784|Multisection^W contrast IS:Find:Pt:Shoulder.left:Doc:CT
C1526784|Shoulder - left CT W contrast IS
C1526784|Multisection^W contrast Intrasynovial:Finding:Point in time:Shoulder.left:Document:Computerized Tomography
C1526784|Should-L CT W contr IS
C1526792|Orbit-L MRI
C1526792|Orbit - left MRI
C1526792|Multisection:Find:Pt:Orbit.left:Doc:MRI
C1526792|Multisection:Finding:Point in time:Orbit.left:Document:MRI
C1526800|Elbow-L XR 2V Obl
C1526800|Elbow - left X-ray 2 views Oblique
C1526800|Views 2 oblique:Find:Pt:Elbow.left:Doc:XR
C1526800|Views 2 oblique:Finding:Point in time:Elbow.left:Document:XR
C1527066|Pancreas MRI
C1527066|Multisection:Find:Pt:Pancreas:Doc:MRI
C1527066|Multisection:Finding:Point in time:Pancreas:Document:MRI
C1524437|Multisection:Finding:Point in time:Posterior fossa:Narrative:COMPUTERIZED TOMOGRAPHY
C1524437|Posterior fossa CT
C1524437|Post fossa CT
C1524437|Multisection:Finding:Point in time:Posterior fossa:Document:Computerized Tomography
C1524437|Multisection:Find:Pt:Posterior fossa:Doc:CT
C1524839|Lower extremity - right CT WO contrast
C1524839|LE-R CT WO contr
C1524839|Multisection^WO contrast:Find:Pt:Lower extremity.right:Doc:CT
C1524839|Multisection^WO contrast:Finding:Point in time:Lower extremity.right:Document:Computerized Tomography
C1525102|Upper extremity joint - left MRI
C1525102|UE joint-L MRI
C1525102|Multisection:Find:Pt:Upper extremity.joint.left:Doc:MRI
C1525102|Multisection:Finding:Point in time:Upper extremity.joint.left:Document:MRI
C1525103|UE joint-R MRI
C1525103|Upper extremity joint - right MRI
C1525103|Multisection:Find:Pt:Upper extremity.joint.right:Doc:MRI
C1525103|Multisection:Finding:Point in time:Upper extremity.joint.right:Document:MRI
C1524451|Brain MRI Ltd W contr IV
C1524451|Brain MRI limited W contrast IV
C1524451|Multisection limited^W contrast IV:Find:Pt:Brain:Doc:MRI
C1524451|Multisection limited^W contrast Intravenous:Finding:Point in time:Brain:Document:MRI
C1524460|Multisection^W contrast IS:Find:Pt:Ankle.left:Doc:MRI
C1524460|Ankle - left MRI W contrast IS
C1524460|Multisection^W contrast Intrasynovial:Finding:Point in time:Ankle.left:Document:MRI
C1524460|Ankle-L MRI W contr IS
C1525225|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity veins.left:Document:MRI.angio
C1525225|UE vv-L MRI.Angio WO+W contr IV
C1525225|Multisection^WO & W contrast IV:Find:Pt:Upper extremity veins.left:Doc:MRI.angio
C1525225|Upper extremity veins - left MRI angiogram WO and W contrast IV
C1525271|Deprecated Spine CT stereotactic
C1525271|Deprecated Spine CT Stereo
C1525271|Multisection stereotactic:Find:Pt:Spine:Doc:CT
C1525271|Multisection stereotactic:Finding:Point in time:Spine:Document:Computerized Tomography
C1525344|Views ski jump:Find:Pt:Calcaneus:Doc:XR
C1525344|Views ski jump:Finding:Point in time:Calcaneus:Document:XR
C1525344|Deprecated Heel XR Ski Jump
C1525344|Deprecated Calcaneus X-ray ski jump
C1525476|Acetabulum-L XR 2V
C1525476|Acetabulum - left X-ray 2 views
C1525476|Views 2:Finding:Point in time:Acetabulum.left:Document:XR
C1525476|Views 2:Find:Pt:Acetabulum.left:Doc:XR
C1525495|Should-L XR AP+Ax+Y
C1525495|Shoulder - left X-ray AP and axillary and Y
C1525495|Views AP & axillary & Y:Finding:Point in time:Shoulder.left:Document:XR
C1525495|Views AP & axillary & Y:Find:Pt:Shoulder.left:Doc:XR
C1525495|VIEWS AP & AXILLARY & Y:FINDING:POINT IN TIME:SHOULDER.LEFT:NARRATIVE:XR
C1525513|Knee-Bl XR AP+Lat+Tunnel
C1525513|Knee - bilateral X-ray AP and lateral and tunnel
C1525513|Views AP & lateral & tunnel:Finding:Point in time:Knee.bilateral:Document:XR
C1525513|Views AP & lateral & tunnel:Find:Pt:Knee.bilateral:Doc:XR
C1525543|Chest XR PA+Lat+AP l-Lat-Decub
C1525543|Chest X-ray PA and lateral and AP left lateral-decubitus
C1525543|Views PA & lateral & AP L-lateral-decubitus:Find:Pt:Chest:Doc:XR
C1525543|Views PA & lateral & AP L-lateral-decubitus:Finding:Point in time:Chest:Document:XR
C1525548|Patella-L XR PA+Lat+Sunrise
C1525548|Patella - left X-ray PA and lateral and Sunrise
C1525548|Views PA & lateral & Sunrise:Find:Pt:Patella.left:Doc:XR
C1525548|Views PA & lateral & Sunrise:Finding:Point in time:Patella.left:Document:XR
C1525559|Should-L XR Grashey+Ax
C1525559|Shoulder - left X-ray Grashey and axillary
C1525559|Views Grashey & axillary:Find:Pt:Shoulder.left:Doc:XR
C1525559|Views Grashey & axillary:Finding:Point in time:Shoulder.left:Document:XR
C1525637|TMJ CT W contr IV
C1525637|Temporomandibular joint CT W contrast IV
C1525637|Multisection^W contrast IV:Find:Pt:Temporomandibular joint:Doc:CT
C1525637|Multisection^W contrast Intravenous:Finding:Point in time:Temporomandibular joint:Document:Computerized Tomography
C1525657|TMJ-R MRI WO+W contr IV
C1525657|Multisection^WO & W contrast IV:Find:Pt:Temporomandibular joint.right:Doc:MRI
C1525657|Multisection^WO & W contrast Intravenous:Finding:Point in time:Temporomandibular joint.right:Document:MRI
C1525657|Temporomandibular joint - right MRI WO and W contrast IV
C1525686|TMJ-Bl XR
C1525686|Temporomandibular joint - bilateral X-ray
C1525686|Views:Find:Pt:Temporomandibular joint.bilateral:Doc:XR
C1525686|Views:Finding:Point in time:Temporomandibular joint.bilateral:Document:XR
C1525695|L-spine+SIJ XR 5V
C1525695|Spine Lumbar and Sacroiliac Joint X-ray 5 views
C1525695|Views 5:Find:Pt:Spine.lumbar+Sacroiliac joint:Doc:XR
C1525695|Views 5:Finding:Point in time:Spine.lumbar+Sacroiliac joint:Document:XR
C1525704|Aorta+Abd aa XRA W contr IA
C1525704|Abdominal Aorta and Arteries Fluoroscopic angiogram W contrast IA
C1525704|Views^W contrast IA:Find:Pt:Aorta+Abdominal arteries:Doc:XR.fluor.angio
C1525704|Views^W contrast Intra-arterial:Finding:Point in time:Aorta+Abdominal arteries:Document:XR.fluor.angio
C1525721|Extremity arteries - left Fluoroscopic angiogram W contrast IA
C1525721|Extr aa-L XRA W contr IA
C1525721|Views^W contrast Intra-arterial:Finding:Point in time:Extremity arteries.left:Document:XR.fluor.angio
C1525721|Views^W contrast IA:Find:Pt:Extremity arteries.left:Doc:XR.fluor.angio
C1525733|Views^W contrast Intrasynovial:Finding:Point in time:Temporomandibular joint.bilateral:Document:XR.fluor
C1525733|TMJ-Bl Flr W contr IS
C1525733|Views^W contrast IS:Find:Pt:Temporomandibular joint.bilateral:Doc:XR.fluor
C1525733|Temporomandibular joint - bilateral Fluoroscopy W contrast IS
C1525760|Multisection^WO contrast:Find:Pt:Chest>Lung parenchyma:Doc:CT
C1525760|Multisection^WO contrast:Finding:Point in time:Chest>Lung parenchyma:Document:Computerized Tomography
C1525760|Lung parenchyma CT WO contr
C1525760|Lung parenchyma CT WO contrast
C1525768|Wrist - bilateral CT WO contrast
C1525768|Wrist-Bl CT WO contr
C1525768|Multisection^WO contrast:Find:Pt:Wrist.bilateral:Doc:CT
C1525768|Multisection^WO contrast:Finding:Point in time:Wrist.bilateral:Document:Computerized Tomography
C1525861|XXX Flr W Ba via Fistula
C1525861|Unspecified body region Fluoroscopy W barium contrast via fistula
C1525861|Views^W barium contrast via fistula:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1525861|Views^W barium contrast via fistula:Find:Pt:XXX:Doc:XR.fluor
C1525866|Wrist-Bl Flr W contr IS
C1525866|Views^W contrast IS:Find:Pt:Wrist.bilateral:Doc:XR.fluor
C1525866|Views^W contrast Intrasynovial:Finding:Point in time:Wrist.bilateral:Document:XR.fluor
C1525866|Wrist - bilateral Fluoroscopy W contrast IS
C1525875|Views^WO & W weight:Finding:Point in time:Acromioclavicular joint:Document:XR
C1525875|Views^WO & W weight:Find:Pt:Acromioclavicular joint:Doc:XR
C1525875|AC joint XR WO+W Wt
C1525875|Acromioclavicular Joint X-ray WO and W weight
C1525811|Thoracic Spine vessels MRI angiogram WO and W contrast IV
C1525811|T-spine ves MRI.Angio WO+W contr IV
C1525811|Multisection^WO & W contrast IV:Find:Pt:Spine.thoracic vessels:Doc:MRI.angio
C1525811|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.thoracic vessels:Document:MRI.angio
C1525832|Toe 2nd-L XR
C1525832|Toe second - left X-ray
C1525832|Views:Find:Pt:Toe.second.left:Doc:XR
C1525832|Views:Finding:Point in time:Toe.second.left:Document:XR
C1525979|AC joint-R XR WO+W Wt
C1525979|Acromioclavicular joint - right X-ray WO and W weight
C1525979|Views^WO & W weight:Find:Pt:Acromioclavicular joint.right:Doc:XR
C1525979|Views^WO & W weight:Finding:Point in time:Acromioclavicular joint.right:Document:XR
C1525989|Ankle - right X-ray W manual stress
C1525989|Ankle-R XR W Stress
C1525989|Views^W manual stress:Find:Pt:Ankle.right:Doc:XR
C1525989|Views^W manual stress:Finding:Point in time:Ankle.right:Document:XR
C1526133|Should XR AP+Lat
C1526133|Shoulder X-ray AP and lateral
C1526133|Views AP & lateral:Finding:Point in time:Shoulder:Document:XR
C1526133|Views AP & lateral:Find:Pt:Shoulder:Doc:XR
C1526039|Hip-R XR AP+Lat Xtable
C1526039|Hip - right X-ray AP and lateral crosstable
C1526039|Views AP & lateral crosstable:Find:Pt:Hip.right:Doc:XR
C1526039|Views AP & lateral crosstable:Finding:Point in time:Hip.right:Document:XR
C1526145|Sinuses X-ray 2 views
C1526145|Sinuses XR 2V
C1526145|Views 2:Finding:Point in time:Sinuses:Document:XR
C1526145|Views 2:Find:Pt:Sinuses:Doc:XR
C1526155|Sinuses XR Waters
C1526155|Sinuses X-ray Waters
C1526155|View Waters:Finding:Point in time:Sinuses:Document:XR
C1526155|View Waters:Find:Pt:Sinuses:Doc:XR
C1526186|T-spine XR 3V
C1526186|Views 3:Find:Pt:Spine.thoracic:Doc:XR
C1526186|Views 3:Finding:Point in time:Spine.thoracic:Document:XR
C1526186|Thoracic spine X-ray 3 views
C1526216|Elbow - right Fluoroscopy W contrast IS
C1526216|Views^W contrast Intrasynovial:Finding:Point in time:Elbow.right:Document:XR.fluor
C1526216|Elbow-R Flr W contr IS
C1526216|Views^W contrast IS:Find:Pt:Elbow.right:Doc:XR.fluor
C1526236|Subclavian v XRA W contr IV
C1526236|Subclavian vein Fluoroscopic angiogram W contrast IV
C1526236|Views^W contrast Intravenous:Finding:Point in time:Subclavian vein:Document:XR.fluor.angio
C1526236|Views^W contrast IV:Find:Pt:Subclavian vein:Doc:XR.fluor.angio
C1525136|T-spine XR Lat W FE
C1525136|Views lateral^W flexion & W extension:Finding:Point in time:Spine.thoracic:Document:XR
C1525136|Views lateral^W flexion & W extension:Find:Pt:Spine.thoracic:Doc:XR
C1525136|Thoracic spine X-ray lateral W flexion and W extension
C1526268|US Guidance for needle biopsy of Kidney - bilateral
C1526268|Guidance for biopsy.needle:Find:Pt:Kidney.bilateral:Doc:US
C1526268|Guidance for biopsy.needle:Finding:Point in time:Kidney.bilateral:Document:Ultrasound
C1526268|Kdny-Bl US Bx needle guid
C1524501|Elbow CT W contr IV
C1524501|Elbow CT W contrast IV
C1524501|Multisection^W contrast IV:Find:Pt:Elbow:Doc:CT
C1524501|Multisection^W contrast Intravenous:Finding:Point in time:Elbow:Document:Computerized Tomography
C1524854|Foot - left MRI WO contrast
C1524854|Ft-L MRI WO contr
C1524854|Multisection^WO contrast:Finding:Point in time:Foot.left:Document:MRI
C1524854|Multisection^WO contrast:Find:Pt:Foot.left:Doc:MRI
C1524859|Forearm - left MRI WO contrast
C1524859|Forearm-L MRI WO contr
C1524859|Multisection^WO contrast:Finding:Point in time:Forearm.left:Document:MRI
C1524859|Multisection^WO contrast:Find:Pt:Forearm.left:Doc:MRI
C1524864|Hand-L MRI WO contr
C1524864|Hand - left MRI WO contrast
C1524864|Multisection^WO contrast:Finding:Point in time:Hand.left:Document:MRI
C1524864|Multisection^WO contrast:Find:Pt:Hand.left:Doc:MRI
C1524514|UE-R CT W contr IV
C1524514|Upper extremity - right CT W contrast IV
C1524514|Multisection^W contrast IV:Find:Pt:Upper extremity.right:Doc:CT
C1524514|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.right:Document:Computerized Tomography
C1524529|Forearm CT W contr IV
C1524529|Forearm CT W contrast IV
C1524529|Multisection^W contrast IV:Find:Pt:Forearm:Doc:CT
C1524529|Multisection^W contrast Intravenous:Finding:Point in time:Forearm:Document:Computerized Tomography
C1524897|Mandible CT WO contr
C1524897|Mandible CT WO contrast
C1524897|Multisection^WO contrast:Finding:Point in time:Mandible:Document:Computerized Tomography
C1524897|Multisection^WO contrast:Find:Pt:Mandible:Doc:CT
C1524924|UE ves MRI.Angio WO contr
C1524924|Upper extremity vessels MRI angiogram WO contrast
C1524924|Multisection^WO contrast:Find:Pt:Upper extremity vessels:Doc:MRI.angio
C1524924|Multisection^WO contrast:Finding:Point in time:Upper extremity vessels:Document:MRI.angio
C1524558|Knee-Bl MRI W contr IV
C1524558|Knee - bilateral MRI W contrast IV
C1524558|Multisection^W contrast IV:Find:Pt:Knee.bilateral:Doc:MRI
C1524558|Multisection^W contrast Intravenous:Finding:Point in time:Knee.bilateral:Document:MRI
C1524563|Larynx CT W contr IV
C1524563|Larynx CT W contrast IV
C1524563|Multisection^W contrast Intravenous:Finding:Point in time:Neck>Larynx:Document:Computerized Tomography
C1524563|Multisection^W contrast IV:Find:Pt:Neck>Larynx:Doc:CT
C1524581|Sacrum+Coccyx MRI W contr IV
C1524581|Sacrum and Coccyx MRI W contrast IV
C1524581|Multisection^W contrast IV:Find:Pt:Sacrum+Coccyx:Doc:MRI
C1524581|Multisection^W contrast Intravenous:Finding:Point in time:Sacrum+Coccyx:Document:MRI
C1524206|Finger fifth X-ray AP single view
C1524206|Finger.5th XR AP 1V
C1524206|View AP:Find:Pt:Finger.fifth:Doc:XR
C1524206|View AP:Finding:Point in time:Finger.fifth:Document:XR
C1524219|Knee-Bl XR AP+Lat
C1524219|Knee - bilateral X-ray AP and lateral
C1524219|Views AP & lateral:Finding:Point in time:Knee.bilateral:Document:XR
C1524219|Views AP & lateral:Find:Pt:Knee.bilateral:Doc:XR
C1524600|Chest vessels CT angiogram W contrast IV
C1524600|Multisection^W contrast IV:Find:Pt:Chest>Vessels:Doc:CT.angio
C1524600|Multisection^W contrast Intravenous:Finding:Point in time:Chest>Vessels:Document:Computerized Tomography.angio
C1524600|Chest Ves CT.Angio W contr IV
C1524622|Ankle - left X-ray 3 views
C1524622|Ankle-L XR 3V
C1524622|Views 3:Finding:Point in time:Ankle.left:Document:XR
C1524622|Views 3:Find:Pt:Ankle.left:Doc:XR
C1524977|Hand - bilateral X-ray
C1524977|Hand-Bl XR
C1524977|Views:Finding:Point in time:Hand.bilateral:Document:XR
C1524977|Views:Find:Pt:Hand.bilateral:Doc:XR
C1524311|Fluoroscopy Guidance for placement of catheter in Unspecified body region
C1524311|XXX Flr Cath plac guid
C1524311|Guidance for placement of catheter:Find:Pt:XXX:Doc:XR.fluor
C1524311|Guidance for placement of catheter:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1524327|Brst-L CT Localization guid
C1524327|CT Guidance for localization of Breast - left
C1524327|Guidance for localization:Finding:Point in time:Breast.left:Document:Computerized Tomography
C1524327|Guidance for localization:Find:Pt:Breast.left:Doc:CT
C1524335|Spine Flr PC Vertebroplasty guid
C1524335|Fluoroscopy Guidance for percutaneous vertebroplasty of Spine
C1524335|Guidance for percutaneous vertebroplasty:Finding:Point in time:Spine:Document:XR.fluor
C1524335|Guidance for percutaneous vertebroplasty:Find:Pt:Spine:Doc:XR.fluor
C1526996|Multisection:Find:Pt:Chest+Abdomen>Aorta:Doc:CT
C1526996|Multisection:Finding:Point in time:Chest+Abdomen>Aorta:Document:Computerized Tomography
C1526996|Chest and Abdomen Aorta CT
C1526996|Chest+Abd Aorta CT
C1524344|Multisection:Find:Pt:Abdomen>Aorta.abdominal:Doc:CT
C1524344|Multisection:Finding:Point in time:Abdomen>Aorta.abdominal:Document:Computerized Tomography
C1524344|Abd Aorta CT
C1524344|Abdominal Aorta CT
C1524345|Ab Ao MRI
C1524345|Aorta abdominal MRI
C1524345|Multisection:Find:Pt:Aorta.abdominal:Doc:MRI
C1524345|Multisection:Finding:Point in time:Aorta.abdominal:Document:MRI
C1524350|Brst-R MRI
C1524350|Breast - right MRI
C1524350|Multisection:Finding:Point in time:Breast.right:Document:MRI
C1524350|Multisection:Find:Pt:Breast.right:Doc:MRI
C1524637|Knee - left X-ray 3 views
C1524637|Knee-L XR 3V
C1524637|Views 3:Find:Pt:Knee.left:Doc:XR
C1524637|Views 3:Finding:Point in time:Knee.left:Document:XR
C1524657|C-spine XR 4V
C1524657|Views 4:Find:Pt:Spine.cervical:Doc:XR
C1524657|Views 4:Finding:Point in time:Spine.cervical:Document:XR
C1524657|Cervical spine X-ray 4 views
C1524749|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip.left:Document:MRI
C1524749|Multisection^WO & W contrast IV:Find:Pt:Hip.left:Doc:MRI
C1524749|Hip-L MRI WO+W contr IV
C1524749|Hip - left MRI WO and W contrast IV
C1524761|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sacroiliac joint:Document:Computerized Tomography
C1524761|Sacroiliac Joint CT WO and W contrast IV
C1524761|Multisection^WO & W contrast IV:Find:Pt:Sacroiliac joint:Doc:CT
C1524761|SIJ CT WO+W contr IV
C1524762|SIJ MRI WO+W contr IV
C1524762|Multisection^WO & W contrast IV:Find:Pt:Sacroiliac joint:Doc:MRI
C1524762|Sacroiliac Joint MRI WO and W contrast IV
C1524762|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sacroiliac joint:Document:MRI
C1524801|LE vv MRI.Angio WO+W contr IV
C1524801|Multisection^WO & W contrast IV:Find:Pt:Lower extremity veins:Doc:MRI.angio
C1524801|Lower extremity veins MRI angiogram WO and W contrast IV
C1524801|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity veins:Document:MRI.angio
C1524808|Multisection^WO & W contrast IV:Find:Pt:Neck vessels:Doc:MRI.angio
C1524808|Neck vessels MRI angiogram WO and W contrast IV
C1524808|Neck ves MRI.Angio WO+W contr IV
C1524808|Multisection^WO & W contrast Intravenous:Finding:Point in time:Neck vessels:Document:MRI.angio
C1830220|Multisection^W contrast Intrasynovial:Finding:Point in time:Elbow:Document:MRI
C1830220|Elbow MRI W contrast IS
C1830220|Elbow MRI W contr IS
C1830220|Multisection^W contrast IS:Find:Pt:Elbow:Doc:MRI
C1715393|Guidance.stereotactic for localization^WO & W contrast IV:Find:Pt:Brain:Doc:MRI
C1715393|MRI Guidance.stereotactic for localization in Brain-- WO and W contrast IV
C1715393|Guidance.stereotactic for localization^WO & W contrast Intravenous:Finding:Point in time:Brain:Document:MRI
C1715393|Brain MRI Local Str Guid WO+W contr IV
C1715407|Hrt PET
C1715407|Heart PET
C1715407|Multisection:Finding:Point in time:Heart:Document:Radnuc.PET
C1715407|Multisection:Find:Pt:Heart:Doc:Radnuc.PET
C1715485|Liver Flr Bx needle guid W contr IV
C1715485|Fluoroscopy Guidance for needle biopsy of Liver-- W contrast IV
C1715485|Guidance for biopsy.needle^W contrast IV:Find:Pt:Liver:Doc:XR.fluor
C1715485|Guidance for biopsy.needle^W contrast Intravenous:Finding:Point in time:Liver:Document:XR.fluor
C1715493|Views^W Tc-99m glucoheptonate IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1715493|Kidney - bilateral Scan W Tc-99m glucoheptonate IV
C1715493|Views^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1715493|Kdny-Bl RI W Tc99mGHA IV
C1633404|Portal v XRA Cath plac guid W contr IV
C1633404|Fluoroscopic angiogram Guidance for placement of catheter in Portal vein-- W contrast IV
C1633404|Guidance for placement of catheter^W contrast IV:Find:Pt:Portal vein:Doc:XR.fluor.angio
C1633404|Guidance for placement of catheter^W contrast Intravenous:Finding:Point in time:Portal vein:Document:XR.fluor.angio
C1645313|Multisection & 3D reconstruction:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1645313|Deprecated XXX CT +3DR
C1645313|Multisection & 3D reconstruction:Find:Pt:XXX:Doc:CT
C1645313|Deprecated Unspecified body region CT and 3D reconstruction
C1635070|Multisection^W endorectal coil:Find:Pt:Pelvis:Doc:MRI
C1635070|Pelvis MRI W endorectal coil
C1635070|Multisection^W endorectal coil:Finding:Point in time:Pelvis:Document:MRI
C1714497|Renal ves RI Flow W Tc99mGHA IV
C1714497|Renal vessels Scan flow W Tc-99m glucoheptonate IV
C1714497|Views flow^W Tc-99m glucoheptonate IV:Find:Pt:Renal vessels:Doc:Radnuc
C1714497|Views flow^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Renal vessels:Document:Radnuc
C1637794|Chest US Tube plac guid
C1637794|US Guidance for placement of tube in Chest
C1637794|Guidance for placement of tube:Find:Pt:Chest:Doc:US
C1637794|Guidance for placement of tube:Finding:Point in time:Chest:Document:Ultrasound
C1644658|Hrt RI 2V Rest+W Tl201 IV
C1644658|Heart Scan 2 views at rest and W Tl-201 IV
C1644658|Views 2^at rest & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1644658|Views 2^at rest & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1652991|Chest and Abdomen CT W contrast IV
C1652991|Chest+Abd CT W contr IV
C1652991|Multisection^W contrast Intravenous:Finding:Point in time:Chest+Abdomen:Document:Computerized Tomography
C1652991|Multisection^W contrast IV:Find:Pt:Chest+Abdomen:Doc:CT
C1631787|Guidance for drainage of abscess:Find:Pt:Kidney:Doc:CT
C1631787|CT Guidance for drainage of abscess of Kidney
C1631787|Guidance for drainage of abscess:Finding:Point in time:Kidney:Document:Computerized Tomography
C1631787|Kidney CT Abscess drain guid
C1644663|EU ves CT.Angio W contr IV
C1644663|Multisection^W contrast IV:Find:Pt:Upper extremity>Vessels:Doc:CT.angio
C1644663|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity>Vessels:Document:Computerized Tomography.angio
C1644663|Upper extremity Vessels CT angiogram W contrast IV
C1978440|Deprecated Views AP & lateral:Finding:Point in time:Abdomen:Narrative:XR
C1978440|Deprecated Abd XR AP+Lat
C1978440|Deprecated Abdomen X-ray AP & lateral
C1978440|Views AP & lateral:Find:Pt:Abdomen:Nar:XR
C1978440|Views AP & lateral:Finding:Point in time:Abdomen:Narrative:XR
C1978759|LE-Bl CT W contr IV
C1978759|Lower extremity - bilateral CT W contrast IV
C1978759|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.bilateral:Document:Computerized Tomography
C1978759|Multisection^W contrast IV:Find:Pt:Lower extremity.bilateral:Doc:CT
C1954305|LE v-R US
C1954305|Lower extremity vein - right US
C1954305|Multisection:Find:Pt:Lower extremity vein.right:Doc:US
C1954305|Multisection:Finding:Point in time:Lower extremity vein.right:Document:Ultrasound
C2923659|Deprecated Cht>Ht.LA+Pul v CT.Angio +3DR
C2923659|Multisection & 3D reconstruction^W contrast IV:Find:Pt:Chest>Heart.atrium.left+Pulmonary veins:Doc:CT.angio
C2923659|Deprecated Chest>Heart.atrium.left+Pulmonary veins CT angiogram and 3D reconstruction W contrast IV
C2923659|Multisection & 3D reconstruction^W contrast Intravenous:Finding:Point in time:Chest>Heart.atrium.left+Pulmonary veins:Document:Computerized Tomography.angio
C3175181|Fluoroscopy Guidance for catheterization of Fallopian tube - left-- transcervical
C3175181|FT-L Flr Cath guid transcervical
C3175181|Guidance for catheterization^transcervical:Finding:Point in time:Fallopian tube.left:Document:XR.fluor
C3175181|Guidance for catheterization^transcervical:Find:Pt:Fallopian tube.left:Doc:XR.fluor
C3174367|Kidney - left Fluoroscopy View for cyst examination
C3174367|Kidney-L Flr View for cyst exam
C3174367|View for cyst examination:Finding:Point in time:Kidney.left:Document:XR.fluor
C3174367|View for cyst examination:Find:Pt:Kidney.left:Doc:XR.fluor
C3173625|Renal vessels - right Fluoroscopic angiogram W contrast
C3173625|Renal ves-R XRA W contr
C3173625|Views^W contrast:Finding:Point in time:Renal vessels.right:Document:XR.fluor.angio
C3173625|Views^W contrast:Find:Pt:Renal vessels.right:Doc:XR.fluor.angio
C3169578|Fluoroscopic angiogram Guidance for placement of ilio-iliac tube endoprosthesis in Iliac artery - left-- W contrast IA
C3169578|Iliac a-L XRA Ilio tube guid W contr IA
C3169578|Guidance for placement of ilio-iliac tube endoprosthesis^W contrast IA:Find:Pt:Iliac artery.left:Doc:XR.fluor.angio
C3169578|Guidance for placement of ilio-iliac tube endoprosthesis^W contrast Intra-arterial:Finding:Point in time:Iliac artery.left:Document:XR.fluor.angio
C3533360|Abdomen and Pelvis MRI W contrast PO and WO and W contrast IV
C3533360|Abd+Pelvis MRI W contr PO+WO+W IV
C3533360|Multisection^W contrast Oral+WO & W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis:Document:MRI
C3533360|Multisection^W contrast PO+WO & W contrast IV:Find:Pt:Abdomen+Pelvis:Doc:MRI
C1525319|Hip - left X-ray lateral crosstable
C1525319|Hip-L XR Lat Xtable
C1525319|Hip - left X-ray and lateral crosstable
C1525319|Hip-L XR +Lat Xtable
C1525319|View lateral crosstable:Finding:Point in time:Hip.left:Document:XR
C1525319|Views & lateral crosstable:Find:Pt:Hip.left:Doc:XR
C1525319|View lateral crosstable:Find:Pt:Hip.left:Doc:XR
C1525319|Views & lateral crosstable:Finding:Point in time:Hip.left:Document:XR
C3262970|Wrist - left X-ray 3 views scaphoid
C3262970|Wrist-L XR 3V scaphoid
C3262970|Views 3 scaphoid:Finding:Point in time:Wrist.left:Document:XR
C3262970|Views 3 scaphoid:Find:Pt:Wrist.left:Doc:XR
C3263005|Lower leg-Bl MRI WO contr
C3263005|Lower leg - bilateral MRI WO contrast
C3263005|Multisection^WO contrast:Find:Pt:Lower leg.bilateral:Doc:MRI
C3263005|Multisection^WO contrast:Finding:Point in time:Lower leg.bilateral:Document:MRI
C3483139|C-spine CT Nerve Block guid
C3483139|Guidance for nerve block:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C3483139|Guidance for nerve block:Find:Pt:Spine.cervical:Doc:CT
C3483139|CT Guidance for nerve block of Cervical spine
C3263024|Nasal bones MRI
C3263024|Multisection:Finding:Point in time:Nasal bones:Document:MRI
C3263024|Multisection:Find:Pt:Nasal bones:Doc:MRI
C3263027|Multisection^WO & W contrast Intravenous:Finding:Point in time:Finger.right:Document:MRI
C3263027|Finger-R MRI WO+W contr IV
C3263027|Multisection^WO & W contrast IV:Find:Pt:Finger.right:Doc:MRI
C3263027|Finger - right MRI WO and W contrast IV
C3263060|Fluoroscopy Guidance for percutaneous needle biopsy of Salivary gland
C3263060|Salivary gland Flr PC Bx needle guid
C3263060|Guidance for percutaneous biopsy.needle:Find:Pt:Salivary gland:Doc:XR.fluor
C3263060|Guidance for percutaneous biopsy.needle:Finding:Point in time:Salivary gland:Document:XR.fluor
C3263064|Breast Mammogram Post Wire Placement
C3263064|Brst Mam p wire plac
C3263064|Views^post wire placement:Finding:Point in time:Breast:Document:Mam
C3263064|Views^post wire placement:Find:Pt:Breast:Doc:Mam
C3262915|CT Guidance for biopsy of Liver-- WO contrast
C3262915|Liver CT Bx guid WO contr
C3262915|Guidance for biopsy^WO contrast:Find:Pt:Abdomen>Liver:Doc:CT
C3262915|Guidance for biopsy^WO contrast:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C0942166|Scapula-R XR
C0942166|Scapula - right X-ray
C0942166|Views:Find:Pt:Scapula.right:Doc:XR
C0942166|Views:Finding:Point in time:Scapula.right:Document:XR
C0942176|Toes - bilateral X-ray
C0942176|Toes-Bl XR
C0942176|Views:Finding:Point in time:Toes.bilateral:Document:XR
C0942176|Views:Find:Pt:Toes.bilateral:Doc:XR
C0945319|Femoral artery - left Fluoroscopic angiogram runoff W contrast IA
C0945319|Fem a-L XRA Runoff W contr IA
C0945319|View runoff^W contrast IA:Find:Pt:Femoral artery.left:Doc:XR.fluor.angio
C0945319|View runoff^W contrast Intra-arterial:Finding:Point in time:Femoral artery.left:Document:XR.fluor.angio
C0942187|Fem a-R XRA Runoff W contr IA
C0942187|Femoral artery - right Fluoroscopic angiogram runoff W contrast IA
C0942187|View runoff^W contrast Intra-arterial:Finding:Point in time:Femoral artery.right:Document:XR.fluor.angio
C0942187|View runoff^W contrast IA:Find:Pt:Femoral artery.right:Doc:XR.fluor.angio
C0942204|Knee-L MRI WO+W contr IV
C0942204|Multisection^WO & W contrast IV:Find:Pt:Knee.left:Doc:MRI
C0942204|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee.left:Document:MRI
C0942204|Knee - left MRI WO and W contrast IV
C0945323|Elbow-Bl MRI
C0945323|Elbow - bilateral MRI
C0945323|Multisection:Find:Pt:Elbow.bilateral:Doc:MRI
C0945323|Multisection:Finding:Point in time:Elbow.bilateral:Document:MRI
C0942224|Elbow - right MRI
C0942224|Elbow-R MRI
C0942224|Multisection:Finding:Point in time:Elbow.right:Document:MRI
C0942224|Multisection:Find:Pt:Elbow.right:Doc:MRI
C0942272|Wrist - bilateral US
C0942272|Wrist-Bl US
C0942272|Multisection:Find:Pt:Wrist.bilateral:Doc:US
C0942272|Multisection:Finding:Point in time:Wrist.bilateral:Document:Ultrasound
C0942283|Breast - right US limited
C0942283|Brst-R US Ltd
C0942283|Multisection limited:Find:Pt:Breast.right:Doc:US
C0942283|Multisection limited:Finding:Point in time:Breast.right:Document:Ultrasound
C0942332|Brst-R Mam Dx
C0942332|Breast - right Mammogram diagnostic
C0942332|Views diagnostic:Finding:Point in time:Breast.right:Document:Mam
C0942332|Views diagnostic:Find:Pt:Breast.right:Doc:Mam
C0882027|Mesenteric artery Fluoroscopic angiogram W contrast IA
C0882027|Mesenteric a XRA W contr IA
C0882027|Views^W contrast Intra-arterial:Finding:Point in time:Mesenteric artery:Document:XR.fluor.angio
C0882027|Views^W contrast IA:Find:Pt:Mesenteric artery:Doc:XR.fluor.angio
C0882543|Patella X-ray 2 views
C0882543|Patella XR 2V
C0882543|Views 2:Find:Pt:Patella:Doc:XR
C0882543|Views 2:Finding:Point in time:Patella:Document:XR
C0882099|Views:Finding:Point in time:Sinuses:Narrative:XR
C0882099|Sinuses X-ray
C0882099|Sinuses XR
C0882099|Views:Find:Pt:Sinuses:Doc:XR
C0882099|Views:Finding:Point in time:Sinuses:Document:XR
C0882136|L-spine Flr W contr IT
C0882136|Views^W contrast IT:Find:Pt:Spine.lumbar:Doc:XR.fluor
C0882136|Views^W contrast Intrathecal:Finding:Point in time:Spine.lumbar:Document:XR.fluor
C0882136|Lumbar spine Fluoroscopy W contrast IT
C0882557|Multisection:Finding:Point in time:Spine.thoracic:Narrative:MRI
C0882557|T-spine MRI
C0882557|Multisection:Find:Pt:Spine.thoracic:Doc:MRI
C0882557|Multisection:Finding:Point in time:Spine.thoracic:Document:MRI
C0882557|Thoracic spine MRI
C0882162|Scrotum+Test US
C0882162|Scrotum and Testicle US
C0882162|Multisection:Find:Pt:Scrotum+Testicle:Doc:US
C0882162|Multisection:Finding:Point in time:Scrotum+Testicle:Document:Ultrasound
C0882210|XXX MRI W conscious sedation
C0882210|Unspecified body region MRI W conscious sedation
C0882210|Multisection^W conscious sedation:Find:Pt:XXX:Doc:MRI
C0882210|Multisection^W conscious sedation:Finding:Point in time:To be specified in another part of the message:Document:MRI
C0942111|Scrotum+Test-Bl RI W Tc99mP IV
C0942111|Scrotum and Testicle - bilateral Scan W Tc-99m pertechnetate IV
C0942111|Views^W Tc-99m pertechnetate Intravenous:Finding:Point in time:Scrotum+Testicle.bilateral:Document:Radnuc
C0942111|Views^W Tc-99m pertechnetate IV:Find:Pt:Scrotum+Testicle.bilateral:Doc:Radnuc
C0945313|Foot - right X-ray
C0945313|Ft-R XR
C0945313|Views:Find:Pt:Foot.right:Doc:XR
C0945313|Views:Finding:Point in time:Foot.right:Document:XR
C0882516|Ankle X-ray 2 views
C0882516|Ankle XR 2V
C0882516|Views 2:Finding:Point in time:Ankle:Document:XR
C0882516|Views 2:Find:Pt:Ankle:Doc:XR
C0881796|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen:Document:MRI
C0881796|Multisection^WO & W contrast IV:Find:Pt:Abdomen:Doc:MRI
C0881796|Abdomen MRI WO and W contrast IV
C0881796|Abd MRI WO+W contr IV
C0881831|Mammogram Guidance for needle localization of mass of Breast
C0881831|Brst Mam Needle local mass guid
C0881831|Guidance for needle localization of mass:Finding:Point in time:Breast:Document:Mam
C0881831|Guidance for needle localization of mass:Find:Pt:Breast:Doc:Mam
C0882525|Chest XR PA+R-Lat+R-Obl+L-Obl Upr Port
C0882525|Chest X-ray PA and right lateral and right oblique and left oblique upright portable
C0882525|Views PA & R-lateral & R-oblique & L-oblique upright portable:Find:Pt:Chest:Doc:XR
C0882525|Views PA & R-lateral & R-oblique & L-oblique upright portable:Finding:Point in time:Chest:Document:XR
C0881881|Chest Flr Image intensifier in Surg
C0881881|Chest Fluoroscopy Image intensifier during surgery
C0881881|Image intensifier^during surgery:Finding:Point in time:Chest:Document:XR.fluor
C0881881|Image intensifier^during surgery:Find:Pt:Chest:Doc:XR.fluor
C0881906|Esoph+HP XRVideo W contr PO Swlw
C0881906|Esophagus and Hypopharynx Fluoroscopy video W contrast PO during swallowing
C0881906|Views^W contrast Oral during swallowing:Finding:Point in time:Esophagus+Hypopharynx:Document:XR.fluor.video
C0881906|Views^W contrast PO during swallowing:Find:Pt:Esophagus+Hypopharynx:Doc:XR.fluor.video
C0881907|Esoph+HP XRVideo W Liq+Paste contr Swlw
C0881907|Esophagus and Hypopharynx Fluoroscopy video W liquid and paste contrast PO during swallowing
C0881907|Views^W liquid & paste contrast PO during swallowing:Find:Pt:Esophagus+Hypopharynx:Doc:XR.fluor.video
C0881907|Views^W liquid & paste contrast Oral during swallowing:Finding:Point in time:Esophagus+Hypopharynx:Document:XR.fluor.video
C0881931|Gallbladder US
C0881931|GB US
C0881931|Multisection:Find:Pt:Gallbladder:Doc:US
C0881931|Multisection:Finding:Point in time:Gallbladder:Document:Ultrasound
C0882533|Views 2:Finding:Point in time:Hand:Narrative:XR
C0882533|Hand XR 2V
C0882533|Hand X-ray 2 views
C0882533|Views 2:Find:Pt:Hand:Doc:XR
C0882533|Views 2:Finding:Point in time:Hand:Document:XR
C0881953|IAC+Post fossa MRI
C0881953|Internal auditory canal and Posterior fossa MRI
C0881953|Multisection:Find:Pt:Internal auditory canal+Posterior fossa:Doc:MRI
C0881953|Multisection:Finding:Point in time:Internal auditory canal+Posterior fossa:Document:MRI
C0881958|Heart MRI
C0881958|Hrt MRI
C0881958|Multisection:Finding:Point in time:Heart:Narrative:MRI
C0881958|Multisection:Finding:Point in time:Heart:Document:MRI
C0881958|Multisection:Find:Pt:Heart:Doc:MRI
C0881961|Hrt XRVideo
C0881961|Heart Fluoroscopy video
C0881961|Views:Find:Pt:Heart:Doc:XR.fluor.video
C0881961|Views:Finding:Point in time:Heart:Document:XR.fluor.video
C0881975|Deprecated Kidney - bilateral and Collecting system CT
C0881975|Multisection:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:Computerized Tomography
C0881975|Multisection:Find:Pt:Kidney.bilateral+Collecting system:Nar:CT
C0881975|Deprecated KD-Bl+CS CT
C1114483|Orbit - bilateral MRI WO contrast
C1114483|Orbit-Bl MRI WO contr
C1114483|Multisection^WO contrast:Find:Pt:Orbit.bilateral:Doc:MRI
C1114483|Multisection^WO contrast:Finding:Point in time:Orbit.bilateral:Document:MRI
C1114511|Lower extremity MRI
C1114511|LE MRI
C1114511|Multisection:Find:Pt:Lower extremity:Doc:MRI
C1114511|Multisection:Finding:Point in time:Lower extremity:Document:MRI
C1114539|C-spine XR AP 1V
C1114539|View AP:Find:Pt:Spine.cervical:Doc:XR
C1114539|View AP:Finding:Point in time:Spine.cervical:Document:XR
C1114539|Cervical spine X-ray AP single view
C1114552|Chest X-ray right or-left oblique portable
C1114552|Chest XR R-or-L-Obl port
C1114552|Views R-or-L-oblique portable:Finding:Point in time:Chest:Document:XR
C1114552|Views R-or-L-oblique portable:Find:Pt:Chest:Doc:XR
C1114940|Shoulder X-ray Single view portable
C1114940|Should XR 1V port
C1114940|View 1 portable:Finding:Point in time:Shoulder:Document:XR
C1114940|View 1 portable:Find:Pt:Shoulder:Doc:XR
C1114566|T-spine XR Lat
C1114566|View lateral:Find:Pt:Spine.thoracic:Doc:XR
C1114566|View lateral:Finding:Point in time:Spine.thoracic:Document:XR
C1114566|Thoracic spine X-ray lateral
C1114944|Pelvis XR 3V
C1114944|Pelvis X-ray 3 views
C1114944|Views 3:Find:Pt:Pelvis:Doc:XR
C1114944|Views 3:Finding:Point in time:Pelvis:Document:XR
C1114604|MRI Guidance.stereotactic for localization in Brain-- WO contrast
C1114604|Brain MRI Local Str Guid WO contr
C1114604|Guidance.stereotactic for localization^WO contrast:Finding:Point in time:Brain:Document:MRI
C1114604|Guidance.stereotactic for localization^WO contrast:Find:Pt:Brain:Doc:MRI
C1114625|Orbit Vv XRA W contr IV
C1114625|Orbit veins Fluoroscopic angiogram W contrast IV
C1114625|Views^W contrast IV:Find:Pt:Orbit veins:Doc:XR.fluor.angio
C1114625|Views^W contrast Intravenous:Finding:Point in time:Orbit veins:Document:XR.fluor.angio
C1114633|Renal a-Bl XRA W contr IA
C1114633|Renal artery - bilateral Fluoroscopic angiogram W contrast IA
C1114633|Views^W contrast IA:Find:Pt:Renal artery.bilateral:Doc:XR.fluor.angio
C1114633|Views^W contrast Intra-arterial:Finding:Point in time:Renal artery.bilateral:Document:XR.fluor.angio
C1114953|Head veins MRI angiogram
C1114953|Head vv MRI.Angio
C1114953|Multisection:Find:Pt:Head veins:Doc:MRI.angio
C1114953|Multisection:Finding:Point in time:Head veins:Document:MRI.angio
C1114678|Views:Finding:Point in time:Coccyx:Narrative:XR
C1114678|Coccyx XR
C1114678|Coccyx X-ray
C1114678|Views:Finding:Point in time:Coccyx:Document:XR
C1114678|Views:Find:Pt:Coccyx:Doc:XR
C2718103|Deprecated Upper extremity vessels MRI angio Multisection W contrast IV
C2718103|Deprecated MRI.Angio
C2718103|Multisection^W contrast.XXX IV:Find:Pt:Vessel.upper extremity:Nar:MRI.angio
C2718103|Multisection^W contrast.XXX Intravenous:Finding:Point in time:Vessel.upper extremity:Narrative:MRI.angio
C1114924|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head>Vessels:Document:Computerized Tomography.angio
C1114924|Multisection^WO & W contrast IV:Find:Pt:Head>Vessels:Doc:CT.angio
C1114924|Head vess CT.Angio WO+W contr IV
C1114924|Head vessels CT angiogram WO and W contrast IV
C1114432|Pancreas CT Bx guid
C1114432|CT Guidance for biopsy of Pancreas
C1114432|Guidance for biopsy:Find:Pt:Abdomen>Pancreas:Doc:CT
C1114432|Guidance for biopsy:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C1114454|UE CT W contr IV
C1114454|Upper extremity CT W contrast IV
C1114454|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity:Document:Computerized Tomography
C1114454|Multisection^W contrast IV:Find:Pt:Upper extremity:Doc:CT
C1114475|US Guidance for aspiration of cyst of Breast
C1114475|Brst US Cyst Asp guid
C1114475|Guidance for aspiration of cyst:Find:Pt:Breast:Doc:US
C1114475|Guidance for aspiration of cyst:Finding:Point in time:Breast:Document:Ultrasound
C1543449|Wrist-R XR 3V+Ulnar Deviation
C1543449|Wrist - right X-ray 3 views and ulnar deviation
C1543449|Views 3 & ulnar deviation:Find:Pt:Wrist.right:Doc:XR
C1543449|Views 3 & ulnar deviation:Finding:Point in time:Wrist.right:Document:XR
C1543803|RI Tum local guid Ltd W Tc99mMIBI IV
C1543803|Scan Guidance for localization of tumor limited-- W Tc-99m Sestamibi IV
C1543803|Guidance for localization of tumor limited^W Tc-99m Sestamibi IV:Find:Pt:^Patient:Doc:Radnuc
C1543803|Guidance for localization of tumor limited^W Tc-99m Sestamibi Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542925|Hrt RI Flow W Tc99mP IV
C1542925|Heart Scan flow W Tc-99m pertechnetate IV
C1542925|Views flow^W Tc-99m pertechnetate Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542925|Views flow^W Tc-99m pertechnetate IV:Find:Pt:Heart:Doc:Radnuc
C1543917|GB RI EF W Tc99mDISIDA IV
C1543917|Gallbladder Scan ejection fraction W Tc-99m DISIDA IV
C1543917|Views ejection fraction^W Tc-99m DISIDA IV:Find:Pt:Gallbladder:Doc:Radnuc
C1543917|Views ejection fraction^W Tc-99m DISIDA Intravenous:Finding:Point in time:Gallbladder:Document:Radnuc
C1543575|Lower extremity artery - left US.doppler
C1543575|LE a-L DOP
C1543575|Multisection:Finding:Point in time:Lower extremity artery.left:Document:Ultrasound.doppler
C1543575|Multisection:Find:Pt:Lower extremity artery.left:Doc:US.doppler
C1543215|Carot a.cervical XRA W contr IA
C1543215|Carotid artery.cervical Fluoroscopic angiogram W contrast IA
C1543215|Views^W contrast IA:Find:Pt:Carotid artery.cervical:Doc:XR.fluor.angio
C1543215|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.cervical:Document:XR.fluor.angio
C1526774|Hip-R XR in Surg
C1526774|Hip - right X-ray during surgery
C1526774|View^during surgery:Finding:Point in time:Hip.right:Document:XR
C1526774|View^during surgery:Find:Pt:Hip.right:Doc:XR
C1526793|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee vessels.left:Document:MRI.angio
C1526793|Knee ves-L MRI.Angio WO+W contr IV
C1526793|Multisection^WO & W contrast IV:Find:Pt:Knee vessels.left:Doc:MRI.angio
C1526793|Knee vessels - left MRI angiogram WO and W contrast IV
C1526814|Shoulder - left X-ray Y
C1526814|Should-L XR Y
C1526814|View Y:Finding:Point in time:Shoulder.left:Document:XR
C1526814|View Y:Find:Pt:Shoulder.left:Doc:XR
C2713073|Abd+Fetus XR FTA
C2713073|Abdomen and Fetus X-ray for fetal age
C2713073|Views for fetal age:Find:Pt:Abdomen+Fetus:Doc:XR
C2713073|Views for fetal age:Finding:Point in time:Abdomen+Fetus:Document:XR
C1527063|Neck CT
C1527063|Multisection:Finding:Point in time:Neck:Narrative:Computerized Tomography
C1527063|Multisection:Find:Pt:Neck:Doc:CT
C1527063|Multisection:Finding:Point in time:Neck:Document:Computerized Tomography
C1524190|Renal vein MRI angiogram
C1524190|Renal v MRI.Angio
C1524190|Multisection:Find:Pt:Renal vein:Doc:MRI.angio
C1524190|Multisection:Finding:Point in time:Renal vein:Document:MRI.angio
C1524832|Elbow - right CT WO contrast
C1524832|Elbow-R CT WO contr
C1524832|Multisection^WO contrast:Find:Pt:Elbow.right:Doc:CT
C1524832|Multisection^WO contrast:Finding:Point in time:Elbow.right:Document:Computerized Tomography
C1524834|Lower extremity - bilateral CT WO contrast
C1524834|LE-Bl CT WO contr
C1524834|Multisection^WO contrast:Finding:Point in time:Lower extremity.bilateral:Document:Computerized Tomography
C1524834|Multisection^WO contrast:Find:Pt:Lower extremity.bilateral:Doc:CT
C1525099|Fluoroscopy Guidance for injection of Joint
C1525099|Joint Flr Inj guid
C1525099|Guidance for injection:Finding:Point in time:Joint:Document:XR.fluor
C1525099|Guidance for injection:Find:Pt:Joint:Doc:XR.fluor
C1525185|Hepatic artery CT angiogram W contrast IA
C1525185|Multisection^W contrast IA:Find:Pt:Abdomen>Hepatic artery:Doc:CT.angio
C1525185|Multisection^W contrast Intra-arterial:Finding:Point in time:Abdomen>Hepatic artery:Document:Computerized Tomography.angio
C1525185|Abd>Hep a CT.Angio W contr IA
C1524452|UE CT Ltd W contr IV
C1524452|Upper extremity CT limited W contrast IV
C1524452|Multisection limited^W contrast IV:Find:Pt:Upper extremity:Doc:CT
C1524452|Multisection limited^W contrast Intravenous:Finding:Point in time:Upper extremity:Document:Computerized Tomography
C1524243|Brst-Bl MRI Dyn W contr IV
C1524243|Breast - bilateral MRI dynamic W contrast IV
C1524243|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Breast.bilateral:Document:MRI
C1524243|Multisection dynamic^W contrast IV:Find:Pt:Breast.bilateral:Doc:MRI
C1525320|Knee X-ray lateral crosstable
C1525320|Knee XR Lat Xtable
C1525320|View lateral crosstable:Find:Pt:Knee:Doc:XR
C1525320|View lateral crosstable:Finding:Point in time:Knee:Document:XR
C1525238|Shoulder vessels - left MRI angiogram WO and W contrast IV
C1525238|Should ves-L MRI.Angio WO+W contr IV
C1525238|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder vessels.left:Document:MRI.angio
C1525238|Multisection^WO & W contrast IV:Find:Pt:Shoulder vessels.left:Doc:MRI.angio
C1525248|Ovary MRI WO contrast
C1525248|Ovary MRI WO contr
C1525248|Multisection^WO contrast:Finding:Point in time:Ovary:Document:MRI
C1525248|Multisection^WO contrast:Find:Pt:Ovary:Doc:MRI
C1525478|Chest X-ray 2 views W nipple markers
C1525478|Chest XR 2V W nipple markers
C1525478|Views 2^W nipple markers:Finding:Point in time:Chest:Document:XR
C1525478|Views 2^W nipple markers:Find:Pt:Chest:Doc:XR
C1525566|Should-L XR Grashey+West Point
C1525566|Shoulder - left X-ray Grashey and West Point
C1525566|Views Grashey & West Point:Finding:Point in time:Shoulder.left:Document:XR
C1525566|Views Grashey & West Point:Find:Pt:Shoulder.left:Doc:XR
C1525572|Femoral artery Fluoroscopic angiogram W contrast IA
C1525572|Fem a XRA W contr IA
C1525572|Views^W contrast IA:Find:Pt:Femoral artery:Doc:XR.fluor.angio
C1525572|Views^W contrast Intra-arterial:Finding:Point in time:Femoral artery:Document:XR.fluor.angio
C1525574|Iliac artery - bilateral Fluoroscopic angiogram W contrast IA
C1525574|Iliac a-Bl XRA W contr IA
C1525574|Views^W contrast Intra-arterial:Finding:Point in time:Iliac artery.bilateral:Document:XR.fluor.angio
C1525574|Views^W contrast IA:Find:Pt:Iliac artery.bilateral:Doc:XR.fluor.angio
C1525582|Views^W contrast IS:Find:Pt:Ankle.left:Doc:XR.fluor
C1525582|Ankle-L Flr W contr IS
C1525582|Ankle - left Fluoroscopy W contrast IS
C1525582|Views^W contrast Intrasynovial:Finding:Point in time:Ankle.left:Document:XR.fluor
C1527061|Mediastinum MRI
C1527061|Multisection:Finding:Point in time:Mediastinum:Document:MRI
C1527061|Multisection:Find:Pt:Mediastinum:Doc:MRI
C1525693|Temporomandibular joint - bilateral X-ray 5 views
C1525693|TMJ-Bl XR 5V
C1525693|Views 5:Finding:Point in time:Temporomandibular joint.bilateral:Document:XR
C1525693|Views 5:Find:Pt:Temporomandibular joint.bilateral:Doc:XR
C1525707|Ac arch+Carot a XRA W contr IA
C1525707|Aortic arch and Carotid artery Fluoroscopic angiogram W contrast IA
C1525707|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery:Document:XR.fluor.angio
C1525707|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery:Doc:XR.fluor.angio
C1524693|Wrist CT W contr IV
C1524693|Wrist CT W contrast IV
C1524693|Multisection^W contrast IV:Find:Pt:Wrist:Doc:CT
C1524693|Multisection^W contrast Intravenous:Finding:Point in time:Wrist:Document:Computerized Tomography
C1525763|Wrist - left X-ray 3 views
C1525763|Wrist-L XR 3V
C1525763|Views 3:Find:Pt:Wrist.left:Doc:XR
C1525763|Views 3:Finding:Point in time:Wrist.left:Document:XR
C1525841|Hip - left X-ray oblique crosstable
C1525841|Hip-L XR Obl Xtable
C1525841|View oblique crosstable:Find:Pt:Hip.left:Doc:XR
C1525841|View oblique crosstable:Finding:Point in time:Hip.left:Document:XR
C1525960|Wrist - right X-ray oblique
C1525960|Wrist-R XR Obl
C1525960|Views oblique:Find:Pt:Wrist.right:Doc:XR
C1525960|Views oblique:Finding:Point in time:Wrist.right:Document:XR
C1525990|Ankle - right X-ray tomograph
C1525990|Ankle-R XRTomo
C1525990|Multisection:Finding:Point in time:Ankle.right:Document:XR.tomo
C1525990|Multisection:Find:Pt:Ankle.right:Doc:XR.tomo
C1526027|Hand-R XR AP+Lat+Obl
C1526027|Hand - right X-ray AP and lateral and oblique
C1526027|Views AP & lateral & oblique:Find:Pt:Hand.right:Doc:XR
C1526027|Views AP & lateral & oblique:Finding:Point in time:Hand.right:Document:XR
C1526110|Should-R XR Y
C1526110|Shoulder - right X-ray Y
C1526110|View Y:Find:Pt:Shoulder.right:Doc:XR
C1526110|View Y:Finding:Point in time:Shoulder.right:Document:XR
C1526111|Should-R XR Grashey+Ax+Outlet
C1526111|Shoulder - right X-ray Grashey and axillary and outlet
C1526111|Views Grashey & axillary & outlet:Finding:Point in time:Shoulder.right:Document:XR
C1526111|Views Grashey & axillary & outlet:Find:Pt:Shoulder.right:Doc:XR
C1526114|Should-R XR West Point
C1526114|Shoulder - right X-ray West Point
C1526114|View West Point:Finding:Point in time:Shoulder.right:Document:XR
C1526114|View West Point:Find:Pt:Shoulder.right:Doc:XR
C1526118|Thumb-R XR AP+Lat+Obl
C1526118|Thumb - right X-ray AP and lateral and oblique
C1526118|Views AP & lateral & oblique:Finding:Point in time:Thumb.right:Document:XR
C1526118|Views AP & lateral & oblique:Find:Pt:Thumb.right:Doc:XR
C1526142|Shoulder X-ray tomograph
C1526142|Should XRTomo
C1526142|Multisection:Find:Pt:Shoulder:Doc:XR.tomo
C1526142|Multisection:Finding:Point in time:Shoulder:Document:XR.tomo
C1526151|Sinuses XR PA+Lat+Waters
C1526151|Sinuses X-ray PA and lateral and Waters
C1526151|Views PA & lateral & Waters:Find:Pt:Sinuses:Doc:XR
C1526151|Views PA & lateral & Waters:Finding:Point in time:Sinuses:Document:XR
C1526207|Ribs Ant XR
C1526207|Ribs anterior X-ray
C1526207|Views:Finding:Point in time:Ribs.anterior:Document:XR
C1526207|Views:Find:Pt:Ribs.anterior:Doc:XR
C1526239|Spine thoracolumbar junction XR AP+Lat
C1526239|Spine Thoracolumbar Junction X-ray AP and lateral
C1526239|Views AP & lateral:Finding:Point in time:Spine.thoracolumbar junction:Document:XR
C1526239|Views AP & lateral:Find:Pt:Spine.thoracolumbar junction:Doc:XR
C1526241|Upper extremity vessels Fluoroscopic angiogram W contrast
C1526241|UE ves XRA W contr
C1526241|Views^W contrast:Find:Pt:Upper extremity vessels:Doc:XR.fluor.angio
C1526241|Views^W contrast:Finding:Point in time:Upper extremity vessels:Document:XR.fluor.angio
C1525137|Aorta US Ltd
C1525137|Aorta US limited
C1525137|Multisection limited:Finding:Point in time:Aorta:Document:Ultrasound
C1525137|Multisection limited:Find:Pt:Aorta:Doc:US
C1526264|Brst-L US PC Bx CN guid
C1526264|US Guidance for core needle percutaneous biopsy of Breast - left
C1526264|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast.left:Document:Ultrasound
C1526264|Guidance for percutaneous biopsy.core needle:Find:Pt:Breast.left:Doc:US
C1526331|Sinuses X-ray Waters upright
C1526331|Sinuses XR Waters Upr
C1526331|View Waters upright:Find:Pt:Sinuses:Doc:XR
C1526331|View Waters upright:Finding:Point in time:Sinuses:Document:XR
C1526300|Brst implant-L Mam
C1526300|Breast implant - left Mammogram
C1526300|Views:Find:Pt:Breast implant.left:Doc:Mam
C1526300|Views:Finding:Point in time:Breast implant.left:Document:Mam
C1524472|Multisection^W contrast Intrasynovial:Finding:Point in time:Shoulder:Document:Computerized Tomography
C1524472|Shoulder CT W contrast IS
C1524472|Should CT W contr IS
C1524472|Multisection^W contrast IS:Find:Pt:Shoulder:Doc:CT
C1524855|Foot - right CT WO contrast
C1524855|Ft-R CT WO contr
C1524855|Multisection^WO contrast:Find:Pt:Foot.right:Doc:CT
C1524855|Multisection^WO contrast:Finding:Point in time:Foot.right:Document:Computerized Tomography
C1524541|Upper arm CT W contr IV
C1524541|Upper arm CT W contrast IV
C1524541|Multisection^W contrast IV:Find:Pt:Upper arm:Doc:CT
C1524541|Multisection^W contrast Intravenous:Finding:Point in time:Upper arm:Document:Computerized Tomography
C1524898|Nasopharynx MRI WO contrast
C1524898|Nasoph MRI WO contr
C1524898|Multisection^WO contrast:Find:Pt:Nasopharynx:Doc:MRI
C1524898|Multisection^WO contrast:Finding:Point in time:Nasopharynx:Document:MRI
C1524212|Hip - left X-ray AP single view
C1524212|Hip-L XR AP 1V
C1524212|View AP:Finding:Point in time:Hip.left:Document:XR
C1524212|View AP:Find:Pt:Hip.left:Doc:XR
C1524285|Brst CT Asp guid
C1524285|CT Guidance for aspiration of Breast
C1524285|Guidance for aspiration:Finding:Point in time:Breast:Document:Computerized Tomography
C1524285|Guidance for aspiration:Find:Pt:Breast:Doc:CT
C1524125|Brst-Bl MRI WO+W contr IV
C1524125|Breast - bilateral MRI WO and W contrast IV
C1524125|Multisection^WO & W contrast IV:Find:Pt:Breast.bilateral:Doc:MRI
C1524125|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast.bilateral:Document:MRI
C1524623|Face XR 3V
C1524623|Facial bones X-ray 3 views
C1524623|Views 3:Finding:Point in time:Facial bones:Document:XR
C1524623|Views 3:Find:Pt:Facial bones:Doc:XR
C1524155|Ft-Bl XR 2V
C1524155|Foot - bilateral X-ray 2 views
C1524155|Views 2:Find:Pt:Foot.bilateral:Doc:XR
C1524155|Views 2:Finding:Point in time:Foot.bilateral:Document:XR
C1524364|Extr XRTomo
C1524364|Extremity X-ray tomograph
C1524364|Multisection:Find:Pt:Extremity:Doc:XR.tomo
C1524364|Multisection:Finding:Point in time:Extremity:Document:XR.tomo
C1524379|Femur X-ray tomograph
C1524379|Femur XRTomo
C1524379|Multisection:Find:Pt:Femur:Doc:XR.tomo
C1524379|Multisection:Finding:Point in time:Femur:Document:XR.tomo
C1524742|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hand.right:Document:MRI
C1524742|Hand - right MRI WO and W contrast IV
C1524742|Multisection^WO & W contrast IV:Find:Pt:Hand.right:Doc:MRI
C1524742|Hand-R MRI WO+W contr IV
C1525024|Ankle-L XR AP+Lat
C1525024|Ankle - left X-ray AP and lateral
C1525024|Views AP & lateral:Find:Pt:Ankle.left:Doc:XR
C1525024|Views AP & lateral:Finding:Point in time:Ankle.left:Document:XR
C1525036|Ft-L XR AP+Lat
C1525036|Foot - left X-ray AP and lateral
C1525036|Views AP & lateral:Find:Pt:Foot.left:Doc:XR
C1525036|Views AP & lateral:Finding:Point in time:Foot.left:Document:XR
C1525040|Deprecated Calcaneus - left X-ray AP and lateral
C1525040|Views AP & lateral:Finding:Point in time:Calcaneus.left:Document:XR
C1525040|Views AP & lateral:Find:Pt:Calcaneus.left:Doc:XR
C1525040|Deprecated Heel-L XR AP+Lat
C1524406|Hip-Bl MRI
C1524406|Hip - bilateral MRI
C1524406|Multisection:Finding:Point in time:Hip.bilateral:Document:MRI
C1524406|Multisection:Find:Pt:Hip.bilateral:Doc:MRI
C1524407|Hip-L CT
C1524407|Hip - left CT
C1524407|Multisection:Find:Pt:Hip.left:Doc:CT
C1524407|Multisection:Finding:Point in time:Hip.left:Document:Computerized Tomography
C1524419|Upper arm - right MRI
C1524419|Upper arm-R MRI
C1524419|Multisection:Find:Pt:Upper arm.right:Doc:MRI
C1524419|Multisection:Finding:Point in time:Upper arm.right:Document:MRI
C1524798|Uterus MRI WO+W contr IV
C1524798|Uterus MRI WO and W contrast IV
C1524798|Multisection^WO & W contrast IV:Find:Pt:Uterus:Doc:MRI
C1524798|Multisection^WO & W contrast Intravenous:Finding:Point in time:Uterus:Document:MRI
C1524805|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest vessels:Document:MRI.angio
C1524805|Chest vessels MRI angiogram WO and W contrast IV
C1524805|Chest ves MRI.Angio WO+W contr IV
C1524805|Multisection^WO & W contrast IV:Find:Pt:Chest vessels:Doc:MRI.angio
C1525097|Guidance for exchange of nephrostomy tube:Find:Pt:Kidney:Doc:CT
C1525097|Guidance for exchange of nephrostomy tube:Finding:Point in time:Kidney:Document:Computerized Tomography
C1525097|Kidney CT NT exchange guid
C1525097|CT Guidance for exchange of nephrostomy tube of Kidney
C1830179|Bone density:MAric:Pt:Hip.left:Qn:XR.DXA
C1830179|Bone density:Mass Aeric:Point in time:Hip.left:Quantitative:XR.DXA
C1830179|Hip - left DXA Bone density
C1830179|Hip-L DXA BDM
C1830203|UE a-Bl DOP Ltd
C1830203|Upper extremity artery - bilateral US.doppler limited
C1830203|Multisection limited:Find:Pt:Upper extremity artery.bilateral:Doc:US.doppler
C1830203|Multisection limited:Finding:Point in time:Upper extremity artery.bilateral:Document:Ultrasound.doppler
C1715422|Hrt SPECT W DIPY+Tc99mMIBI IV
C1715422|Heart SPECT W dipyridamole and W Tc-99m Sestamibi IV
C1715422|Multisection^W dipyridamole & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1715422|Multisection^W dipyridamole & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1715475|BDs Flr Endo guid W contr retro
C1715475|Fluoroscopy Guidance for endoscopy of Biliary ducts-- W contrast retrograde
C1715475|Guidance for endoscopy^W contrast retrograde:Finding:Point in time:Biliary ducts:Document:XR.fluor
C1715475|Guidance for endoscopy^W contrast retrograde:Find:Pt:Biliary ducts:Doc:XR.fluor
C1632800|Views^W contrast intra multiple ducts:Find:Pt:Breast.duct:Nar:XR
C1632800|Views^W contrast intra multiple ducts:Finding:Point in time:Breast.duct:Narrative:XR
C1632800|Deprecated Breast duct X-ray W contrast intra multiple ducts
C1632800|Deprecated Brst.duct XR W contr intra Dc
C1629070|Ft XR Obl+(AP+Lat) stand
C1629070|Foot X-ray oblique and (AP and lateral) standing
C1629070|Views oblique & (AP & lateral)^standing:Find:Pt:Foot:Doc:XR
C1629070|Views oblique & (AP & lateral)^standing:Finding:Point in time:Foot:Document:XR
C1636065|Foot sesamoid bones X-ray
C1636065|Ft.Sesamoids XR
C1636065|Views:Finding:Point in time:Foot.sesamoid bones:Document:XR
C1636065|Views:Find:Pt:Foot.sesamoid bones:Doc:XR
C1714814|BD+PDs Flr Endo guid 1h p contr retro
C1714814|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 1 hour post contrast retrograde
C1714814|Guidance for endoscopy^1 hour post contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1714814|Guidance for endoscopy^1H post contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1717249|Aorta abdominal Fluoroscopic angiogram runoff W contrast IA
C1717249|Ab Ao XRA Runoff W contr IA
C1717249|Views runoff^W contrast Intra-arterial:Finding:Point in time:Aorta.abdominal:Document:XR.fluor.angio
C1717249|Views runoff^W contrast IA:Find:Pt:Aorta.abdominal:Doc:XR.fluor.angio
C1715099|Brain+IAC MRI
C1715099|Brain and Internal auditory canal MRI
C1715099|Multisection:Find:Pt:Brain+Internal auditory canal:Doc:MRI
C1715099|Multisection:Finding:Point in time:Brain+Internal auditory canal:Document:MRI
C1636061|Spine Lumbar X-ray (AP^W R-bending and W L-bending) and (lateral^W flexion and W extension)
C1636061|L-spine XR (AP W R+L-bending)+(Lat W FE)
C1636061|Views (AP^W R-bending & W L-bending) & (lateral^W flexion & W extension):Find:Pt:Spine.lumbar:Doc:XR
C1636061|Views (AP^W R-bending & W L-bending) & (lateral^W flexion & W extension):Finding:Point in time:Spine.lumbar:Document:XR
C1636071|US Guidance for biopsy of Breast - left
C1636071|Brst-L US Bx guid
C1636071|Guidance for biopsy:Find:Pt:Breast.left:Doc:US
C1636071|Guidance for biopsy:Finding:Point in time:Breast.left:Document:Ultrasound
C1635015|US Guidance for placement of needle wire in Breast
C1635015|Brst US Needle Wire plac guid
C1635015|Guidance for placement of needle wire:Find:Pt:Breast:Doc:US
C1635015|Guidance for placement of needle wire:Finding:Point in time:Breast:Document:Ultrasound
C1630192|US Guidance for drainage of cyst of Kidney
C1630192|Kidney US cyst drain guid
C1630192|Guidance for drainage of cyst:Finding:Point in time:Kidney:Document:Ultrasound
C1630192|Guidance for drainage of cyst:Find:Pt:Kidney:Doc:US
C1638279|CT Guidance for biopsy of Heart
C1638279|Hrt CT Bx guid
C1638279|Guidance for biopsy:Find:Pt:Chest>Heart:Doc:CT
C1638279|Guidance for biopsy:Finding:Point in time:Chest>Heart:Document:Computerized Tomography
C1632989|Carotid artery - left US limited
C1632989|Carot a-L US Ltd
C1632989|Multisection limited:Find:Pt:Carotid artery.left:Doc:US
C1632989|Multisection limited:Finding:Point in time:Carotid artery.left:Document:Ultrasound
C1626770|Deprecated Views portable:Finding:Point in time:Tibia.left+Fibula.left:Narrative:XR
C1626770|Views portable:Find:Pt:Tibia.left+Fibula.left:Nar:XR
C1626770|Deprecated Tib+Fib-L XR port
C1626770|Deprecated Tibia Left & Fibula Left X-ray
C1626770|Views portable:Finding:Point in time:Tibia.left+Fibula.left:Narrative:XR
C1642591|Bone SPECT W In-111 WBC IV
C1642591|Bone SPECT W In-111 tagged WBC IV
C1642591|Multisection^W In-111 tagged WBC IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1642591|Multisection^W In-111 tagged WBC Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1643246|Wrist - right X-ray portable
C1643246|Wrist-R XR port
C1643246|Views portable:Finding:Point in time:Wrist.right:Document:XR
C1643246|Views portable:Find:Pt:Wrist.right:Doc:XR
C1953967|Neck MRI Ltd
C1953967|Neck MRI limited
C1953967|Multisection limited:Finding:Point in time:Neck:Document:MRI
C1953967|Multisection limited:Find:Pt:Neck:Doc:MRI
C1953985|Foot - left X-ray GE 3 views
C1953985|Ft-L XR GE 3V
C1953985|Views GE 3:Finding:Point in time:Foot.left:Document:XR
C1953985|Views GE 3:Find:Pt:Foot.left:Doc:XR
C1952657|TMJ-L XR Open+Closed Mouth
C1952657|Temporomandibular joint - left X-ray open and closed mouth
C1952657|Views open & closed mouth:Find:Pt:Temporomandibular joint.left:Doc:XR
C1952657|Views open & closed mouth:Finding:Point in time:Temporomandibular joint.left:Document:XR
C2923071|Head to thigh PET
C2923071|Multisection:Find:Pt:Head to thigh:Doc:Radnuc.PET
C2923071|Multisection:Finding:Point in time:Head to thigh:Document:Radnuc.PET
C3175183|Mammary artery.internal - right Fluoroscopic angiogram W contrast IA
C3175183|IMAl-R XRA W contr IA
C3175183|Views^W contrast IA:Find:Pt:Mammary artery.internal.right:Doc:XR.fluor.angio
C3175183|Views^W contrast Intra-arterial:Finding:Point in time:Mammary artery.internal.right:Document:XR.fluor.angio
C3169525|Head artery.left+Neck artery.left Fluoroscopic angiogram W contrast IA
C3169525|Head a+Neck a-L XRA W contr IA
C3169525|Views^W contrast Intra-arterial:Finding:Point in time:Head artery.left+Neck artery.left:Document:XR.fluor.angio
C3169525|Views^W contrast IA:Find:Pt:Head artery.left+Neck artery.left:Doc:XR.fluor.angio
C3169527|Fluoroscopic angiogram Guidance for placement of intraperitoneal catheter in Abdomen
C3169527|Abd XRA IP cath plac guide
C3169527|Guidance for placement of intraperitoneal catheter:Finding:Point in time:Abdomen:Document:XR.fluor.angio
C3169527|Guidance for placement of intraperitoneal catheter:Find:Pt:Abdomen:Doc:XR.fluor.angio
C2970309|Thyroid RI +Uptake W I-123 PO
C2970309|Thyroid Scan and uptake W I-123 PO
C2970309|Views & uptake^W I-123 PO:Find:Pt:Thyroid:Doc:Radnuc
C2970309|Views & uptake^W I-123 Oral:Finding:Point in time:Thyroid:Document:Radnuc
C3533554|Guidance for removal of catheter^W contrast Intravenous:Finding:Point in time:Central vein:Document:XR.fluor.angio
C3533554|Fluoroscopic angiogram Guidance for removal of catheter from Central vein-- W contrast IV
C3533554|Centl v XRA cath rem guid W contr IV
C3533554|Guidance for removal of catheter^W contrast IV:Find:Pt:Central vein:Doc:XR.fluor.angio
C3262986|Brst implant-Bl MRI WO+W contr IV
C3262986|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast implant.bilateral:Document:MRI
C3262986|Multisection^WO & W contrast IV:Find:Pt:Breast implant.bilateral:Doc:MRI
C3262986|Breast implant - bilateral MRI WO and W contrast IV
C3483137|L-spine Flr Inj guid
C3483137|Guidance for injection:Find:Pt:Spine.lumbar:Doc:XR.fluor
C3483137|Guidance for injection:Finding:Point in time:Spine.lumbar:Document:XR.fluor
C3483137|Fluoroscopy Guidance for injection of Lumbar spine
C3262468|MRI Guidance for needle biopsy of Thyroid
C3262468|Thyroid MRI Bx needle guid
C3262468|Guidance for biopsy.needle:Find:Pt:Thyroid:Doc:MRI
C3262468|Guidance for biopsy.needle:Finding:Point in time:Thyroid:Document:MRI
C3262470|Multisection^WO & W contrast Intravenous:Finding:Point in time:Finger.left:Document:MRI
C3262470|Multisection^WO & W contrast IV:Find:Pt:Finger.left:Doc:MRI
C3262470|Finger-L MRI WO+W contr IV
C3262470|Finger - left MRI WO and W contrast IV
C3263049|Thyroid RI +Uptake W I-131 PO
C3263049|Thyroid Scan and uptake W I-131 PO
C3263049|Views & uptake^W I-131 PO:Find:Pt:Thyroid:Doc:Radnuc
C3263049|Views & uptake^W I-131 Oral:Finding:Point in time:Thyroid:Document:Radnuc
C3263058|Fluoroscopy Guidance for percutaneous needle biopsy of Kidney
C3263058|Kidney Flr PC Bx needle guid
C3263058|Guidance for percutaneous biopsy.needle:Finding:Point in time:Kidney:Document:XR.fluor
C3263058|Guidance for percutaneous biopsy.needle:Find:Pt:Kidney:Doc:XR.fluor
C3263071|Brst implant-R Mam Dx
C3263071|Breast implant - right Mammogram diagnostic
C3263071|Views diagnostic:Finding:Point in time:Breast implant.right:Document:Mam
C3263071|Views diagnostic:Find:Pt:Breast implant.right:Doc:Mam
C3263079|Should XR Grashey+Ax+ Y
C3263079|Shoulder X-ray Grashey and axillary and Y
C3263079|Views Grashey & axillary & Y:Find:Pt:Shoulder:Doc:XR
C3263079|Views Grashey & axillary & Y:Finding:Point in time:Shoulder:Document:XR
C3263110|Tib+Fib-R XR 1V
C3263110|Tibia - right and Fibula - right X-ray Single view
C3263110|View 1:Finding:Point in time:Tibia.right+Fibula.right:Document:XR
C3263110|View 1:Find:Pt:Tibia.right+Fibula.right:Doc:XR
C3262920|CT Guidance for needle biopsy of Liver
C3262920|Liver CT Bx needle guid
C3262920|Guidance for biopsy.needle:Find:Pt:Abdomen>Liver:Doc:CT
C3262920|Guidance for biopsy.needle:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C0945318|Brst-R Mam Screening
C0945318|Breast - right Mammogram screening
C0945318|Views screening:Finding:Point in time:Breast.right:Document:Mam
C0945318|Views screening:Find:Pt:Breast.right:Doc:Mam
C0942191|Extr-R CT W contr IV
C0942191|Extremity - right CT W contrast IV
C0942191|Multisection^W contrast Intravenous:Finding:Point in time:Extremity.right:Document:Computerized Tomography
C0942191|Multisection^W contrast IV:Find:Pt:Extremity.right:Doc:CT
C0942222|Carot a-R US
C0942222|Carotid artery - right US
C0942222|Multisection:Finding:Point in time:Carotid artery.right:Document:Ultrasound
C0942222|Multisection:Find:Pt:Carotid artery.right:Doc:US
C0942285|Brst-L Mam Bx Str Guid
C0942285|Guidance for stereotactic biopsy:Finding:Point in time:Breast.left:Document:Mam
C0942285|Guidance for stereotactic biopsy:Find:Pt:Breast.left:Doc:Mam
C0942285|Mammogram Guidance for stereotactic biopsy of Breast - left
C0942297|Guidance for placement of large bore catheter into vessel in Central vein - right
C0942297|Cent v-R LB Cath plac guid into ves
C0942297|Guidance for placement of large bore catheter into vessel:Finding:Point in time:Central vein.right:Document
C0942297|Guidance for placement of large bore catheter into vessel:Find:Pt:Central vein.right:Doc
C0942301|Brst-L US Needle local guid
C0942301|US Guidance for needle localization of Breast - left
C0942301|Guidance for needle localization:Finding:Point in time:Breast.left:Document:Ultrasound
C0942301|Guidance for needle localization:Find:Pt:Breast.left:Doc:US
C0942311|Fluoroscopy Guidance for injection of Spine facet joint - right
C0942311|Spine facet joint-R Flr Inj guid
C0942311|Guidance for injection:Finding:Point in time:Spine facet joint.right:Document:XR.fluor
C0942311|Guidance for injection:Find:Pt:Spine facet joint.right:Doc:XR.fluor
C0942342|Knee-L XR AP+PA stand
C0942342|Knee - left X-ray AP and PA standing
C0942342|Views AP & PA^standing:Find:Pt:Knee.left:Doc:XR
C0942342|Views AP & PA^standing:Finding:Point in time:Knee.left:Document:XR
C0882541|Mandible X-ray panorex
C0882541|Mandible XR Panorex
C0882541|View panorex:Finding:Point in time:Mandible:Document:XR
C0882541|View panorex:Find:Pt:Mandible:Doc:XR
C0882028|Views:Finding:Point in time:Nasal bones:Narrative:XR
C0882028|Nasal bones X-ray
C0882028|Nasal bones XR
C0882028|Views:Find:Pt:Nasal bones:Doc:XR
C0882028|Views:Finding:Point in time:Nasal bones:Document:XR
C0882036|Neck US
C0882036|Multisection:Finding:Point in time:Neck:Document:Ultrasound
C0882036|Multisection:Find:Pt:Neck:Doc:US
C0882106|SB Flr W contr PO
C0882106|Small bowel Fluoroscopy W contrast PO
C0882106|Views^W contrast PO:Find:Pt:Small bowel:Doc:XR.fluor
C0882106|Views^W contrast Oral:Finding:Point in time:Small bowel:Document:XR.fluor
C0882116|C-spine MRI W anesthesia
C0882116|Multisection^W anesthesia:Finding:Point in time:Spine.cervical:Document:MRI
C0882116|Multisection^W anesthesia:Find:Pt:Spine.cervical:Doc:MRI
C0882116|Cervical spine MRI W anesthesia
C0882118|C-spine XR 5V
C0882118|Views 5:Finding:Point in time:Spine.cervical:Document:XR
C0882118|Views 5:Find:Pt:Spine.cervical:Doc:XR
C0882118|Cervical spine X-ray 5 views
C0882123|C-spine XR W FE
C0882123|Views^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C0882123|Views^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C0882123|Cervical spine X-ray W flexion and W extension
C0882559|US Guidance for biopsy of Thyroid
C0882559|Thyroid US Bx guid
C0882559|Guidance for biopsy:Find:Pt:Thyroid:Doc:US
C0882559|Guidance for biopsy:Finding:Point in time:Thyroid:Document:Ultrasound
C0882190|Views^W contrast IS:Find:Pt:Wrist:Doc:XR.fluor
C0882190|Wrist Fluoroscopy W contrast IS
C0882190|Wrist Flr W contr IS
C0882190|Views^W contrast Intrasynovial:Finding:Point in time:Wrist:Document:XR.fluor
C0942093|Hip-Bl Flr W contr IS
C0942093|Hip - bilateral Fluoroscopy W contrast IS
C0942093|Views^W contrast IS:Find:Pt:Hip.bilateral:Doc:XR.fluor
C0942093|Views^W contrast Intrasynovial:Finding:Point in time:Hip.bilateral:Document:XR.fluor
C0942123|Views:Find:Pt:Carpal bones.bilateral:Nar:XR
C0942123|Deprecated Carpal bones - bilateral X-ray
C0942123|Deprecated Carpal bones-Bl XR
C0942123|Views:Finding:Point in time:Carpal bones.bilateral:Narrative:XR
C0881805|Retroperitoneum CT
C0881805|Multisection:Find:Pt:Abdomen>Retroperitoneum:Doc:CT
C0881805|Multisection:Finding:Point in time:Abdomen>Retroperitoneum:Document:Computerized Tomography
C0881820|Multisection:Finding:Point in time:Thoracic outlet:Narrative:MRI
C0881820|TO MRI
C0881820|Thoracic outlet MRI
C0881820|Multisection:Find:Pt:Thoracic outlet:Doc:MRI
C0881820|Multisection:Finding:Point in time:Thoracic outlet:Document:MRI
C0881902|Pelvis US transvaginal
C0881902|Pelvis US Transvag
C0881902|Multisection transvaginal:Finding:Point in time:Pelvis:Document:Ultrasound
C0881902|Multisection transvaginal:Find:Pt:Pelvis:Doc:US
C0881925|Views:Finding:Point in time:Femur:Narrative:XR
C0881925|Femur XR
C0881925|Femur X-ray
C0881925|Views:Find:Pt:Femur:Doc:XR
C0881925|Views:Finding:Point in time:Femur:Document:XR
C0882531|Views:Finding:Point in time:Foot:Narrative:XR
C0882531|Ft XR
C0882531|Foot X-ray
C0882531|Views:Find:Pt:Foot:Doc:XR
C0882531|Views:Finding:Point in time:Foot:Document:XR
C0881962|XXX CT W contr IV
C0881962|Unspecified body region CT W contrast IV
C0881962|Multisection^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0881962|Multisection^W contrast IV:Find:Pt:XXX:Doc:CT
C0881998|Abd XR AP (Sup+Upr)
C0881998|Abdomen X-ray AP (supine and upright)
C0881998|Views AP (supine & upright):Finding:Point in time:Abdomen:Document:XR
C0881998|Views AP (supine & upright):Find:Pt:Abdomen:Doc:XR
C0882003|Knee RI W RNC IV
C0882003|Knee Scan
C0882003|Views^W radionuclide Intravenous:Finding:Point in time:Knee:Document:Radnuc
C0882003|Views^W radionuclide IV:Find:Pt:Knee:Doc:Radnuc
C1114580|L-spine XR 3V
C1114580|Views 3:Finding:Point in time:Spine.lumbar:Document:XR
C1114580|Views 3:Find:Pt:Spine.lumbar:Doc:XR
C1114580|Lumbar spine X-ray 3 views
C1114582|L-spine XR AP 1V
C1114582|View AP:Find:Pt:Spine.lumbar:Doc:XR
C1114582|View AP:Finding:Point in time:Spine.lumbar:Document:XR
C1114582|Lumbar spine X-ray AP single view
C1114602|L-spine XR 5V
C1114602|Views 5:Find:Pt:Spine.lumbar:Doc:XR
C1114602|Views 5:Finding:Point in time:Spine.lumbar:Document:XR
C1114602|Lumbar spine X-ray 5 views
C1114948|Maxillofacial region CT WO contrast
C1114948|Maxillofacial CT WO contr
C1114948|Multisection^WO contrast:Find:Pt:Head>Maxillofacial region:Doc:CT
C1114948|Multisection^WO contrast:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1114435|CT Guidance for biopsy of Kidney - bilateral
C1114435|Guidance for biopsy:Find:Pt:Kidney.bilateral:Doc:CT
C1114435|Guidance for biopsy:Finding:Point in time:Kidney.bilateral:Document:Computerized Tomography
C1114435|Kdny-Bl CT Bx guid
C1114476|TO MRI WO contr
C1114476|Thoracic outlet MRI WO contrast
C1114476|Multisection^WO contrast:Find:Pt:Thoracic outlet:Doc:MRI
C1114476|Multisection^WO contrast:Finding:Point in time:Thoracic outlet:Document:MRI
C1543455|Ankle-R XR AP+Lat+Obl stand
C1543455|Ankle - right X-ray AP and lateral and oblique standing
C1543455|Views AP & lateral & oblique^standing:Finding:Point in time:Ankle.right:Document:XR
C1543455|Views AP & lateral & oblique^standing:Find:Pt:Ankle.right:Doc:XR
C1543776|Hrt SPECT PF Rest+stress+W RNC IV
C1543776|Heart SPECT perfusion at rest and W stress and W radionuclide IV
C1543776|Multisection perfusion^at rest & W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543776|Multisection perfusion^at rest & W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543479|Should XR AP(w IR+ER)
C1543479|Shoulder X-ray AP (W internal rotation and W external rotation)
C1543479|View AP (W internal rotation & W external rotation):Finding:Point in time:Shoulder:Document:XR
C1543479|View AP (W internal rotation & W external rotation):Find:Pt:Shoulder:Doc:XR
C1543800|SPECT for Tumor W Tc99mMIBI IV
C1543800|SPECT for tumor W Tc-99m Sestamibi IV
C1543800|Multisection for tumor^W Tc-99m Sestamibi Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543800|Multisection for tumor^W Tc-99m Sestamibi IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543807|Vein RI W Tc99mDTPA IV
C1543807|Vein Scan W Tc-99m DTPA IV
C1543807|Views^W Tc-99m DTPA IV:Find:Pt:Vein:Doc:Radnuc
C1543807|Views^W Tc-99m DTPA Intravenous:Finding:Point in time:Vein:Document:Radnuc
C1542896|Lung RI V W Tc99mDTPA AeroIH
C1542896|Views ventilation^W Tc-99m DTPA aerosol Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1542896|Lung Scan ventilation W Tc-99m DTPA aerosol IH
C1542896|Views ventilation^W Tc-99m DTPA aerosol IH:Find:Pt:Lung:Doc:Radnuc
C1543892|Hrt SPECT BP Rest+W RNC IV
C1543892|Heart SPECT blood pool at rest and W radionuclide IV
C1543892|Multisection blood pool^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543892|Multisection blood pool^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543896|Head Cistern Scan delayed W radionuclide IT
C1543896|Head.cistern RI Delayed W RNC IT
C1543896|Views delayed^W radionuclide IT:Find:Pt:Head.cistern:Doc:Radnuc
C1543896|Views delayed^W radionuclide Intrathecal:Finding:Point in time:Head.cistern:Document:Radnuc
C1543911|Hrt RI FP+EF W RNC IV
C1543911|Heart Scan first pass and ejection fraction
C1543911|Views first pass & ejection fraction^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543911|Views first pass & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543932|Hrt RI FP+WM+EF W RNC IV
C1543932|Heart Scan first pass and wall motion and ejection fraction
C1543932|Views first pass & wall motion & ejection fraction^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543932|Views first pass & wall motion & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543161|AV fistula US
C1543161|AVF US
C1543161|Multisection:Finding:Point in time:AV fistula:Document:Ultrasound
C1543161|Multisection:Find:Pt:AV fistula:Doc:US
C1543184|L-spine XR 5V W FE
C1543184|Views 5^W flexion & W extension:Finding:Point in time:Spine.lumbar:Document:XR
C1543184|Views 5^W flexion & W extension:Find:Pt:Spine.lumbar:Doc:XR
C1543184|Lumbar spine X-ray 5 views W flexion and W extension
C1543216|Carot a+Cerebral a XRA W contr IA
C1543216|Carotid artery and Cerebral artery Fluoroscopic angiogram W contrast IA
C1543216|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Cerebral artery:Document:XR.fluor.angio
C1543216|Views^W contrast IA:Find:Pt:Carotid artery+Cerebral artery:Doc:XR.fluor.angio
C1526751|Should-R XR Grashey+West Point
C1526751|Shoulder - right X-ray Grashey and West Point
C1526751|Views Grashey & West Point:Finding:Point in time:Shoulder.right:Document:XR
C1526751|Views Grashey & West Point:Find:Pt:Shoulder.right:Doc:XR
C1524432|Mandible CT
C1524432|Multisection:Find:Pt:Mandible:Doc:CT
C1524432|Multisection:Finding:Point in time:Mandible:Document:Computerized Tomography
C1524174|Sacrum MRI
C1524174|Multisection:Finding:Point in time:Sacrum:Document:MRI
C1524174|Multisection:Find:Pt:Sacrum:Doc:MRI
C1524811|Ankle - left CT WO contrast
C1524811|Ankle-L CT WO contr
C1524811|Multisection^WO contrast:Finding:Point in time:Ankle.left:Document:Computerized Tomography
C1524811|Multisection^WO contrast:Find:Pt:Ankle.left:Doc:CT
C1524813|Ankle - right CT WO contrast
C1524813|Ankle-R CT WO contr
C1524813|Multisection^WO contrast:Finding:Point in time:Ankle.right:Document:Computerized Tomography
C1524813|Multisection^WO contrast:Find:Pt:Ankle.right:Doc:CT
C1524826|Multisection^WO contrast:Find:Pt:Calcaneus.right:Doc:CT
C1524826|Deprecated Calcaneus - right CT WO contrast
C1524826|Deprecated Heel-R CT WO contr
C1524826|Multisection^WO contrast:Finding:Point in time:Calcaneus.right:Document:Computerized Tomography
C1525176|Knee ves-L MRI.Angio
C1525176|Knee vessels - left MRI angiogram
C1525176|Multisection:Finding:Point in time:Knee vessels.left:Document:MRI.angio
C1525176|Multisection:Find:Pt:Knee vessels.left:Doc:MRI.angio
C1524449|UE joint MRI Ltd
C1524449|Multisection limited:Finding:Point in time:Upper extremity.joint:Document:MRI
C1524449|Multisection limited:Find:Pt:Upper extremity.joint:Doc:MRI
C1524449|Upper extremity.joint MRI limited
C1524450|Abd CT Ltd W contr IV
C1524450|Abdomen CT limited W contrast IV
C1524450|Multisection limited^W contrast IV:Find:Pt:Abdomen:Doc:CT
C1524450|Multisection limited^W contrast Intravenous:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1525283|Adrenal MRI WO+W contr IV
C1525283|Adrenal gland MRI WO and W contrast IV
C1525283|Multisection^WO & W contrast Intravenous:Finding:Point in time:Adrenal gland:Document:MRI
C1525283|Multisection^WO & W contrast IV:Find:Pt:Adrenal gland:Doc:MRI
C1525312|Elbow - left X-ray Jones
C1525312|Elbow-L XR Jones
C1525312|View Jones:Finding:Point in time:Elbow.left:Document:XR
C1525312|View Jones:Find:Pt:Elbow.left:Doc:XR
C1525313|Hip X-ray Judet
C1525313|Hip XR Judet
C1525313|View Judet:Finding:Point in time:Hip:Document:XR
C1525313|View Judet:Find:Pt:Hip:Doc:XR
C1525323|C-spine XR Lat Xtable port
C1525323|View lateral crosstable portable:Find:Pt:Spine.cervical:Doc:XR
C1525323|View lateral crosstable portable:Finding:Point in time:Spine.cervical:Document:XR
C1525323|Cervical spine X-ray lateral crosstable portable
C1525207|Orbit ves MRI.Angio W contr IV
C1525207|Orbit vessels MRI angiogram W contrast IV
C1525207|Multisection^W contrast IV:Find:Pt:Orbit vessels:Doc:MRI.angio
C1525207|Multisection^W contrast Intravenous:Finding:Point in time:Orbit vessels:Document:MRI.angio
C1527070|Salivary gland MRI
C1527070|Multisection:Find:Pt:Salivary gland:Doc:MRI
C1527070|Multisection:Finding:Point in time:Salivary gland:Document:MRI
C1525485|Wrist-L XR 6V
C1525485|Wrist - left X-ray 6 views
C1525485|Views 6:Finding:Point in time:Wrist.left:Document:XR
C1525485|Views 6:Find:Pt:Wrist.left:Doc:XR
C1525520|C-spine XR AP+Odont+Lat Xtable
C1525520|Views AP & odontoid & lateral crosstable:Finding:Point in time:Spine.cervical:Document:XR
C1525520|Views AP & odontoid & lateral crosstable:Find:Pt:Spine.cervical:Doc:XR
C1525520|Cervical spine X-ray AP and odontoid and lateral crosstable
C1525581|Views^W contrast Intrasynovial:Finding:Point in time:Ankle.bilateral:Document:XR.fluor
C1525581|Ankle-Bl Flr W contr IS
C1525581|Views^W contrast IS:Find:Pt:Ankle.bilateral:Doc:XR.fluor
C1525581|Ankle - bilateral Fluoroscopy W contrast IS
C1525589|C-spine Flr W contr ID
C1525589|Views^W contrast intradisc:Find:Pt:Spine.cervical:Doc:XR.fluor
C1525589|Views^W contrast intradisc:Finding:Point in time:Spine.cervical:Document:XR.fluor
C1525589|Cervical spine Fluoroscopy W contrast intradisc
C1525590|L-spine Flr W contr ID
C1525590|Views^W contrast intradisc:Finding:Point in time:Spine.lumbar:Document:XR.fluor
C1525590|Views^W contrast intradisc:Find:Pt:Spine.lumbar:Doc:XR.fluor
C1525590|Lumbar spine Fluoroscopy W contrast intradisc
C1525626|Temporomandibular joint - right MRI
C1525626|TMJ-R MRI
C1525626|Multisection:Find:Pt:Temporomandibular joint.right:Doc:MRI
C1525626|Multisection:Finding:Point in time:Temporomandibular joint.right:Document:MRI
C1525680|Wrist-Bl XR Scaphoid
C1525680|Wrist - bilateral X-ray scaphoid
C1525680|Views scaphoid:Find:Pt:Wrist.bilateral:Doc:XR
C1525680|Views scaphoid:Finding:Point in time:Wrist.bilateral:Document:XR
C1525687|Olecranon - left X-ray
C1525687|Olecranon-L XR
C1525687|Views:Finding:Point in time:Olecranon.left:Document:XR
C1525687|Views:Find:Pt:Olecranon.left:Doc:XR
C1525698|L-spine+Sacrum+SIJ+Coccyx XR 5V
C1525698|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray 5 views
C1525698|Views 5:Find:Pt:Spine.lumbar+Sacrum+Sacroiliac joint+Coccyx:Doc:XR
C1525698|Views 5:Finding:Point in time:Spine.lumbar+Sacrum+Sacroiliac joint+Coccyx:Document:XR
C1525726|Maxillary artery.internal Fluoroscopic angiogram W contrast IA
C1525726|Maxillary a.internal XRA W contr IA
C1525726|Views^W contrast IA:Find:Pt:Maxillary artery.internal:Doc:XR.fluor.angio
C1525726|Views^W contrast Intra-arterial:Finding:Point in time:Maxillary artery.internal:Document:XR.fluor.angio
C1527074|Wrist CT
C1527074|Multisection:Finding:Point in time:Wrist:Document:Computerized Tomography
C1527074|Multisection:Find:Pt:Wrist:Doc:CT
C1525797|Guidance for injection:Finding:Point in time:Spine.cervical>Intervertebral disc:Document:Computerized Tomography
C1525797|Guidance for injection:Find:Pt:Spine.cervical>Intervertebral disc:Doc:CT
C1525797|CT Guidance for injection of Cervical spine Intervertebral disc
C1525797|C-spine interv disc CT Inj guid
C1525844|Wrist-L XR PA+Lat
C1525844|Wrist - left X-ray PA and lateral
C1525844|Views PA & lateral:Finding:Point in time:Wrist.left:Document:XR
C1525844|Views PA & lateral:Find:Pt:Wrist.left:Doc:XR
C1525868|Spine Flr W contr IT
C1525868|Spine Fluoroscopy W contrast IT
C1525868|Views^W contrast Intrathecal:Finding:Point in time:Spine:Document:XR.fluor
C1525868|Views^W contrast IT:Find:Pt:Spine:Doc:XR.fluor
C1525876|Views^WO & W weight:Finding:Point in time:Acromioclavicular joint.bilateral:Document:XR
C1525876|AC joint-Bl XR WO+W Wt
C1525876|Views^WO & W weight:Find:Pt:Acromioclavicular joint.bilateral:Doc:XR
C1525876|Acromioclavicular joint - bilateral X-ray WO and W weight
C1525936|Pelvis XR AP+Inlet
C1525936|Pelvis X-ray AP and inlet
C1525936|Views AP & inlet:Find:Pt:Pelvis:Doc:XR
C1525936|Views AP & inlet:Finding:Point in time:Pelvis:Document:XR
C1526072|Knee-R XR V1 Tunnel stand
C1526072|Knee - right X-ray tunnel standing
C1526072|View tunnel^standing:Find:Pt:Knee.right:Doc:XR
C1526072|View tunnel^standing:Finding:Point in time:Knee.right:Document:XR
C1526080|Lower extremity - right X-ray Single view
C1526080|LE-R XR 1V
C1526080|View 1:Find:Pt:Lower extremity.right:Doc:XR
C1526080|View 1:Finding:Point in time:Lower extremity.right:Document:XR
C1525129|PA-R XRA W contr IA
C1525129|Views^W contrast Intra-arterial:Finding:Point in time:Pulmonary artery.right:Document:XR.fluor.angio
C1525129|Views^W contrast IA:Find:Pt:Pulmonary artery.right:Doc:XR.fluor.angio
C1525129|Right pulmonary artery Fluoroscopic angiogram W contrast IA
C1526140|AC joint XR Zanca
C1526140|Acromioclavicular Joint X-ray Zanca
C1526140|View Zanca:Find:Pt:Acromioclavicular joint:Doc:XR
C1526140|View Zanca:Finding:Point in time:Acromioclavicular joint:Document:XR
C1526171|Thumb XR Lat
C1526171|Thumb X-ray lateral
C1526171|View lateral:Find:Pt:Thumb:Doc:XR
C1526171|View lateral:Finding:Point in time:Thumb:Document:XR
C1526218|Extremity arteries - right Fluoroscopic angiogram W contrast IA
C1526218|Extr aa-R XRA W contr IA
C1526218|Views^W contrast IA:Find:Pt:Extremity arteries.right:Doc:XR.fluor.angio
C1526218|Views^W contrast Intra-arterial:Finding:Point in time:Extremity arteries.right:Document:XR.fluor.angio
C1526234|Sinus v XRA W contr IV
C1526234|Sinus vein Fluoroscopic angiogram W contrast IV
C1526234|Views^W contrast IV:Find:Pt:Sinus vein:Doc:XR.fluor.angio
C1526234|Views^W contrast Intravenous:Finding:Point in time:Sinus vein:Document:XR.fluor.angio
C1526273|XXX US Needle local guid
C1526273|US Guidance for needle localization of Unspecified body region
C1526273|Guidance for needle localization:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1526273|Guidance for needle localization:Find:Pt:XXX:Doc:US
C1526289|Breast implant - left MRI
C1526289|Brst implant-L MRI
C1526289|Multisection:Finding:Point in time:Breast implant.left:Document:MRI
C1526289|Multisection:Find:Pt:Breast implant.left:Doc:MRI
C1526343|Toe fourth - right X-ray
C1526343|Toe 4th-R XR
C1526343|Views:Find:Pt:Toe.fourth.right:Doc:XR
C1526343|Views:Finding:Point in time:Toe.fourth.right:Document:XR
C1526303|Brst specimen-Bl Mam
C1526303|Breast specimen - bilateral Mammogram
C1526303|Views:Find:Pt:Breast specimen.bilateral:Doc:Mam
C1526303|Views:Finding:Point in time:Breast specimen.bilateral:Document:Mam
C1524570|Pancreas MRI W contr IV
C1524570|Pancreas MRI W contrast IV
C1524570|Multisection^W contrast IV:Find:Pt:Pancreas:Doc:MRI
C1524570|Multisection^W contrast Intravenous:Finding:Point in time:Pancreas:Document:MRI
C1524572|Pituitary+ST MRI W contr IV
C1524572|Pituitary and Sella turcica MRI W contrast IV
C1524572|Multisection^W contrast IV:Find:Pt:Pituitary+Sella turcica:Doc:MRI
C1524572|Multisection^W contrast Intravenous:Finding:Point in time:Pituitary+Sella turcica:Document:MRI
C1524582|Scapula-L MRI W contr IV
C1524582|Scapula - left MRI W contrast IV
C1524582|Multisection^W contrast Intravenous:Finding:Point in time:Scapula.left:Document:MRI
C1524582|Multisection^W contrast IV:Find:Pt:Scapula.left:Doc:MRI
C1524211|Hip XR AP 1V
C1524211|Hip X-ray AP single view
C1524211|View AP:Find:Pt:Hip:Doc:XR
C1524211|View AP:Finding:Point in time:Hip:Document:XR
C1524985|Views:Finding:Point in time:Maxilla:Narrative:XR
C1524985|Maxilla X-ray
C1524985|Maxilla XR
C1524985|Views:Finding:Point in time:Maxilla:Document:XR
C1524985|Views:Find:Pt:Maxilla:Doc:XR
C1524324|Stom Flr Endo guid
C1524324|Fluoroscopy Guidance for endoscopy of Stomach
C1524324|Guidance for endoscopy:Find:Pt:Stomach:Doc:XR.fluor
C1524324|Guidance for endoscopy:Finding:Point in time:Stomach:Document:XR.fluor
C1524325|Stom Flr Gastrostomy guid
C1524325|Fluoroscopy Guidance for gastrostomy of Stomach
C1524325|Guidance for gastrostomy:Find:Pt:Stomach:Doc:XR.fluor
C1524325|Guidance for gastrostomy:Finding:Point in time:Stomach:Document:XR.fluor
C1524341|Ankle - left X-ray tomograph
C1524341|Ankle-L XRTomo
C1524341|Multisection:Find:Pt:Ankle.left:Doc:XR.tomo
C1524341|Multisection:Finding:Point in time:Ankle.left:Document:XR.tomo
C1524745|Multisection^WO & W contrast IV:Find:Pt:Hip:Doc:CT
C1524745|Hip CT WO and W contrast IV
C1524745|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip:Document:Computerized Tomography
C1524745|Hip CT WO+W contr IV
C1524754|Upper arm - left MRI WO and W contrast IV
C1524754|Upper arm-L MRI WO+W contr IV
C1524754|Multisection^WO & W contrast IV:Find:Pt:Upper arm.left:Doc:MRI
C1524754|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper arm.left:Document:MRI
C1524764|Multisection^WO & W contrast IV:Find:Pt:Kidney.bilateral:Doc:MRI
C1524764|Kidney - bilateral MRI WO and W contrast IV
C1524764|Multisection^WO & W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:MRI
C1524764|Kdny-Bl MRI WO+W contr IV
C1524391|Forearm - left CT
C1524391|Forearm-L CT
C1524391|Multisection:Find:Pt:Forearm.left:Doc:CT
C1524391|Multisection:Finding:Point in time:Forearm.left:Document:Computerized Tomography
C1524800|Renal vein MRI angiogram WO and W contrast IV
C1524800|Multisection^WO & W contrast Intravenous:Finding:Point in time:Renal vein:Document:MRI.angio
C1524800|Renal v MRI.Angio WO+W contr IV
C1524800|Multisection^WO & W contrast IV:Find:Pt:Renal vein:Doc:MRI.angio
C1830232|Orbit CT WO contrast
C1830232|Orbit CT WO contr
C1830232|Multisection^WO contrast:Find:Pt:Head>Orbit:Doc:CT
C1830232|Multisection^WO contrast:Finding:Point in time:Head>Orbit:Document:Computerized Tomography
C1715374|CT Guidance for procedure of Joint space
C1715374|Joint space CT Procedure guid
C1715374|Guidance for procedure:Finding:Point in time:Joint space:Document:Computerized Tomography
C1715374|Guidance for procedure:Find:Pt:Joint space:Doc:CT
C1715468|Deprecated Knee - bilateral X-ray AP standing
C1715468|Views AP^standing:Find:Pt:Knee.bilateral:Nar:XR
C1715468|Deprecated Knee-Bl XR AP stand
C1715468|Views AP^standing:Finding:Point in time:Knee.bilateral:Narrative:XR
C1715473|C-spine XR GE 4V
C1715473|Views GE 4:Finding:Point in time:Spine.cervical:Document:XR
C1715473|Views GE 4:Find:Pt:Spine.cervical:Doc:XR
C1715473|Cervical spine X-ray GE 4 views
C1715476|Fluoroscopy Guidance for fine needle aspiration of Unspecified body region
C1715476|XXX Flr FNA Asp
C1715476|Guidance for aspiration.fine needle:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1715476|Guidance for aspiration.fine needle:Find:Pt:XXX:Doc:XR.fluor
C1714791|Knee-R MRI Dyn W contr IV
C1714791|Knee - right MRI dynamic W contrast IV
C1714791|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Knee.right:Document:MRI
C1714791|Multisection dynamic^W contrast IV:Find:Pt:Knee.right:Doc:MRI
C1706618|Finger fifth - left X-ray GE 3 views
C1706618|Finger.5th-L XR GE 3V
C1706618|Finger fifth - left Narrative X-ray GE 3 views
C1706618|Views GE 3:Finding:Point in time:Finger.fifth.left:Document:XR
C1706618|Views GE 3:Find:Pt:Finger.fifth.left:Doc:XR
C1714914|Lower leg ves-L MRI.Angio
C1714914|Lower leg vessels - left MRI angiogram
C1714914|Multisection:Find:Pt:Lower leg vessels.left:Doc:MRI.angio
C1714914|Multisection:Finding:Point in time:Lower leg vessels.left:Document:MRI.angio
C1714925|Multisection^W radionuclide Intravenous:Finding:Point in time:To be specified in another part of the message:Narrative:Radnuc.SPECT
C1714925|Unspecified body region SPECT
C1714925|XXX SPECT W RNC IV
C1714925|Multisection^W radionuclide IV:Find:Pt:XXX:Doc:Radnuc.SPECT
C1714925|Multisection^W radionuclide Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Radnuc.SPECT
C1714953|Hip+Thigh US
C1714953|Hip and Thigh US
C1714953|Multisection:Find:Pt:Hip+Thigh:Doc:US
C1714953|Multisection:Finding:Point in time:Hip+Thigh:Document:Ultrasound
C1717222|Brst-Bl US Localization guid
C1717222|US Guidance for localization of Breast - bilateral
C1717222|Guidance for localization:Find:Pt:Breast.bilateral:Doc:US
C1717222|Guidance for localization:Finding:Point in time:Breast.bilateral:Document:Ultrasound
C1715103|Iliac a DOP Ltd
C1715103|Iliac artery US.doppler limited
C1715103|Multisection limited:Finding:Point in time:Iliac artery:Document:Ultrasound.doppler
C1715103|Multisection limited:Find:Pt:Iliac artery:Doc:US.doppler
C1717276|Hrt RI PF Rest+W ADE+Tl201 IV
C1717276|Heart Scan perfusion at rest and W adenosine and W Tl-201 IV
C1717276|Views perfusion^at rest & W adenosine & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1717276|Views perfusion^at rest & W adenosine & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1637280|Brst Flr PC Abscess Drain guid
C1637280|Fluoroscopy Guidance for percutaneous drainage of abscess of Breast
C1637280|Guidance for percutaneous drainage of abscess:Find:Pt:Breast:Doc:XR.fluor
C1637280|Guidance for percutaneous drainage of abscess:Finding:Point in time:Breast:Document:XR.fluor
C1635012|T-spine XR AP W+WO L-bending
C1635012|Views AP^W L-bending & WO bending:Find:Pt:Spine.thoracic:Doc:XR
C1635012|Views AP^W L-bending & WO bending:Finding:Point in time:Spine.thoracic:Document:XR
C1635012|Thoracic spine X-ray AP W left bending and WO bending
C1639903|US Guidance for removal of catheter from Central vein-- Tunneled
C1639903|Centl v US cath rem guid Tunneled
C1639903|Guidance for removal of catheter^tunneled:Finding:Point in time:Central vein:Document:Ultrasound
C1639903|Guidance for removal of catheter^tunneled:Find:Pt:Central vein:Doc:US
C1641048|Deprecated View AP lateral-decubitus:Find:Pt:Chest:Nar:XR
C1641048|View AP lateral-decubitus:Find:Pt:Chest:Nar:XR
C1641048|Deprecated Chest X-ray AP lateral-decubitus
C1641048|Deprecated Chest XR AP Lat Decub
C1641048|View AP lateral-decubitus:Finding:Point in time:Chest:Narrative:XR
C1632380|Views:Finding:Point in time:Sella turcica:Narrative:XR
C1632380|Sella turcica X-ray
C1632380|ST XR
C1632380|Views:Finding:Point in time:Sella turcica:Document:XR
C1632380|Views:Find:Pt:Sella turcica:Doc:XR
C1633478|Breast - left FFD mammogram diagnostic
C1633478|Views diagnostic:Finding:Point in time:Breast.left:Document:Mam.FFD
C1633478|Brst-L FFDM Dx
C1633478|Views diagnostic:Find:Pt:Breast.left:Doc:Mam.FFD
C1624128|Brst Mam XCCL
C1624128|Breast Mammogram XCCL
C1624128|View XCCL:Find:Pt:Breast:Doc:Mam
C1624128|View XCCL:Finding:Point in time:Breast:Document:Mam
C1630180|CT Guidance for needle biopsy of Kidney
C1630180|Kidney CT Bx needle guid
C1630180|Guidance for biopsy.needle:Find:Pt:Kidney:Doc:CT
C1630180|Guidance for biopsy.needle:Finding:Point in time:Kidney:Document:Computerized Tomography
C1624698|Chest and Abdomen X-ray Single view
C1624698|Chest+Abd XR 1V
C1624698|View 1:Find:Pt:Chest+Abdomen:Doc:XR
C1624698|View 1:Finding:Point in time:Chest+Abdomen:Document:XR
C1953969|Knee-R XR AP 1V
C1953969|Knee - right X-ray AP single view
C1953969|View AP:Find:Pt:Knee.right:Doc:XR
C1953969|View AP:Finding:Point in time:Knee.right:Document:XR
C1953972|Skull XR Ltd
C1953972|Skull X-ray limited
C1953972|Views limited:Find:Pt:Skull:Doc:XR
C1953972|Views limited:Finding:Point in time:Skull:Document:XR
C3174153|Lung-R XR W contr IB
C3174153|Lung - right X-ray W contrast intrabronchial
C3174153|Views^W contrast intrabronchial:Finding:Point in time:Lung.right:Document:XR
C3174153|Views^W contrast intrabronchial:Find:Pt:Lung.right:Doc:XR
C3533562|Guidance for facet joint denervation:Find:Pt:Spine.XXX:Doc:XR.fluor
C3533562|Spine Flr FJ DN guid
C3533562|Fluoroscopy Guidance for facet joint denervation of Spine
C3533562|Guidance for facet joint denervation:Finding:Point in time:Spine.To be specified in another part of the message:Document:XR.fluor
C3533800|Pelvis MRI W contrast PR at rest and maxmal sphincter contraction during straining and defecation
C3533800|Multisection^W contrast Rectal at rest & maxmal sphincter contraction during straining & defecation:Finding:Point in time:Pelvis:Document:MRI
C3533800|Multisection^W contrast PR at rest & maxmal sphincter contraction during straining & defecation:Find:Pt:Pelvis:Doc:MRI
C3533800|Pelvis MRI W cntr PR rest+MASC
C3533795|Chst Pulm art CT for PE
C3533795|Multisection for pulmonary embolus:Find:Pt:Chest>Pulmonary arteries:Doc:CT
C3533795|Chest Pulmonary arteries CT for pulmonary embolus
C3533795|Multisection for pulmonary embolus:Finding:Point in time:Chest>Pulmonary arteries:Document:Computerized Tomography
C1525468|Knee - left X-ray tunnel
C1525468|Knee-L XR V1 Tunnel
C1525468|Knee - left X-ray and tunnel
C1525468|Knee-L XR +Tunnel
C1525468|View tunnel:Find:Pt:Knee.left:Doc:XR
C1525468|View tunnel:Finding:Point in time:Knee.left:Document:XR
C1525468|Views & tunnel:Find:Pt:Knee.left:Doc:XR
C1525468|Views & tunnel:Finding:Point in time:Knee.left:Document:XR
C3262473|Hip - left MRI WO and W contrast IS
C3262473|Hip-L MRI WO+W contr IS
C3262473|Multisection^WO & W contrast IS:Find:Pt:Hip.left:Doc:MRI
C3262473|Multisection^WO & W contrast Intrasynovial:Finding:Point in time:Hip.left:Document:MRI
C3263022|Wrist - left and Hand - left MRI
C3263022|Wrist+Hand-L MRI
C3263022|Multisection:Finding:Point in time:Wrist.left+Hand.left:Document:MRI
C3263022|Multisection:Find:Pt:Wrist.left+Hand.left:Doc:MRI
C3263029|Finger-R MRI WO contr
C3263029|Finger - right MRI WO contrast
C3263029|Multisection^WO contrast:Finding:Point in time:Finger.right:Document:MRI
C3263029|Multisection^WO contrast:Find:Pt:Finger.right:Doc:MRI
C3263044|Hrt RI W Stress+W Tc-99m IV
C3263044|Heart Scan W stress and W Tc-99m IV
C3263044|Views^W stress & W Tc-99m Intravenous:Finding:Point in time:Heart:Document:Radnuc
C3263044|Views^W stress & W Tc-99m IV:Find:Pt:Heart:Doc:Radnuc
C3263059|Fluoroscopy Guidance for percutaneous needle biopsy of Liver
C3263059|Liver Flr PC Bx needle guid
C3263059|Guidance for percutaneous biopsy.needle:Finding:Point in time:Liver:Document:XR.fluor
C3263059|Guidance for percutaneous biopsy.needle:Find:Pt:Liver:Doc:XR.fluor
C3263082|Skull X-ray PA
C3263082|Skull XR PA V1
C3263082|View PA:Find:Pt:Skull:Doc:XR
C3263082|View PA:Finding:Point in time:Skull:Document:XR
C3261718|Portal+Hepatic v DOP
C3261718|Portal vein and Hepatic vein US.doppler
C3261718|Multisection:Find:Pt:Portal vein+Hepatic vein:Doc:US.doppler
C3261718|Multisection:Finding:Point in time:Portal vein+Hepatic vein:Document:Ultrasound.doppler
C3263088|Muscle US Bx needle guid
C3263088|US Guidance for needle biopsy of Muscle
C3263088|Guidance for biopsy.needle:Find:Pt:Muscle:Doc:US
C3263088|Guidance for biopsy.needle:Finding:Point in time:Muscle:Document:Ultrasound
C3261476|Hand-R XR 1V
C3261476|Hand - right X-ray Single view
C3261476|View 1:Finding:Point in time:Hand.right:Document:XR
C3261476|View 1:Find:Pt:Hand.right:Doc:XR
C3263221|Kidney Bilateral and Bladder US
C3263221|Multisection:Find:Pt:Kidney.bilateral+Bladder:Doc:US
C3263221|Multisection:Finding:Point in time:Kidney.bilateral+Bladder:Document:Ultrasound
C3263221|Kidney-Bl+Bladder US
C3262898|Fluoroscopy Guidance for biopsy of Salivary gland
C3262898|Salivary gland Flr Bx guid
C3262898|Guidance for biopsy:Find:Pt:Salivary gland:Doc:XR.fluor
C3262898|Guidance for biopsy:Finding:Point in time:Salivary gland:Document:XR.fluor
C3262909|Multisection^WO & W contrast:Find:Pt:Chest+Abdomen>Aorta:Doc:CT
C3262909|Multisection^WO & W contrast:Finding:Point in time:Chest+Abdomen>Aorta:Document:Computerized Tomography
C3262909|Deprecated Chest+Abd>Aorta CT WO+W contr
C3262909|Deprecated Chest+Abdomen>Aorta CT WO and W contrast
C0942181|Wrist-R XR
C0942181|Wrist - right X-ray
C0942181|Views:Finding:Point in time:Wrist.right:Document:XR
C0942181|Views:Find:Pt:Wrist.right:Doc:XR
C0942182|Zygomatic arch-Bl XR
C0942182|Zygomatic arch - bilateral X-ray
C0942182|Views:Find:Pt:Zygomatic arch.bilateral:Doc:XR
C0942182|Views:Finding:Point in time:Zygomatic arch.bilateral:Document:XR
C0942183|Views:Finding:Point in time:Zygomatic arch.leftTiss fixed:Narrative:XR
C0942183|Zygomatic arch-L XR
C0942183|Zygomatic arch - left X-ray
C0942183|Views:Find:Pt:Zygomatic arch.left:Doc:XR
C0942183|Views:Finding:Point in time:Zygomatic arch.left:Document:XR
C0942186|Femoral artery - bilateral Fluoroscopic angiogram runoff W contrast IA
C0942186|Fem a-Bl XRA Runoff W contr IA
C0942186|View runoff^W contrast IA:Find:Pt:Femoral artery.bilateral:Doc:XR.fluor.angio
C0942186|View runoff^W contrast Intra-arterial:Finding:Point in time:Femoral artery.bilateral:Document:XR.fluor.angio
C0942259|Popliteal space-R US
C0942259|Popliteal space - right US
C0942259|Multisection:Finding:Point in time:Popliteal space.right:Document:Ultrasound
C0942259|Multisection:Find:Pt:Popliteal space.right:Doc:US
C0942267|Scrotum+Test-L US
C0942267|Scrotum and Testicle - left US
C0942267|Multisection:Finding:Point in time:Scrotum+Testicle.left:Document:Ultrasound
C0942267|Multisection:Find:Pt:Scrotum+Testicle.left:Doc:US
C0942300|US Guidance for needle localization of Breast - bilateral
C0942300|Brst-Bl US Needle local guid
C0942300|Guidance for needle localization:Find:Pt:Breast.bilateral:Doc:US
C0942300|Guidance for needle localization:Finding:Point in time:Breast.bilateral:Document:Ultrasound
C0942349|BrachCeph a-R XRA Angpsty W contr IA
C0942349|Brachiocephalic artery - right Fluoroscopic angiogram Angioplasty W contrast IA
C0942349|Angioplasty^W contrast IA:Find:Pt:Brachiocephalic artery.right:Doc:XR.fluor.angio
C0942349|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Brachiocephalic artery.right:Document:XR.fluor.angio
C0942366|Ankle - right X-ray 2 views
C0942366|Ankle-R XR 2V
C0942366|Views 2:Finding:Point in time:Ankle.right:Document:XR
C0942366|Views 2:Find:Pt:Ankle.right:Doc:XR
C0882033|Neck MRI
C0882033|Multisection:Finding:Point in time:Neck:Narrative:MRI
C0882033|Multisection:Find:Pt:Neck:Doc:MRI
C0882033|Multisection:Finding:Point in time:Neck:Document:MRI
C0882553|Multisection^WO & W contrast IV:Find:Pt:Spine.cervical:Doc:MRI
C0882553|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.cervical:Document:MRI
C0882553|C-spine MRI WO+W contr IV
C0882553|Cervical spine MRI WO and W contrast IV
C0882141|Multisection^WO & W contrast IV:Find:Pt:Spine.thoracic:Doc:MRI
C0882141|T-spine MRI WO+W contr IV
C0882141|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.thoracic:Document:MRI
C0882141|Thoracic spine MRI WO and W contrast IV
C0882558|Thigh ves MRI.Angio W contr IV
C0882558|Thigh vessels MRI angiogram W contrast IV
C0882558|Multisection^W contrast Intravenous:Finding:Point in time:Thigh vessels:Document:MRI.angio
C0882558|Multisection^W contrast IV:Find:Pt:Thigh vessels:Doc:MRI.angio
C0882215|Vessel Fluoroscopic angiogram Angioplasty W contrast IA
C0882215|Angioplasty^W contrast IA:Find:Pt:Vessel:Doc:XR.fluor.angio
C0882215|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Vessel:Document:XR.fluor.angio
C0882215|Vesl XRA Angpsty W contr IA
C0942110|Knee - right Scan
C0942110|Knee-R RI W RNC IV
C0942110|Views^W radionuclide Intravenous:Finding:Point in time:Knee.right:Document:Radnuc
C0942110|Views^W radionuclide IV:Find:Pt:Knee.right:Doc:Radnuc
C0942120|Deprecated Calcaneus - bilateral X-ray standing
C0942120|Views:Finding:Point in time:Calcaneus.bilateral:Document:XR
C0942120|Deprecated Heel-Bl XR stand
C0942120|Views:Find:Pt:Calcaneus.bilateral:Doc:XR
C0942120|Deprecated Views:Find:Pt:Calcaneus.bilateral:Doc:XR
C0942146|Acetabulum-L XR
C0942146|Acetabulum - left X-ray
C0942146|Views:Find:Pt:Acetabulum.left:Doc:XR
C0942146|Views:Finding:Point in time:Acetabulum.left:Document:XR
C0881774|Abdomen RUQ US
C0881774|Abd.RUQ US
C0881774|Multisection:Find:Pt:Abdomen.RUQ:Doc:US
C0881774|Multisection:Finding:Point in time:Abdomen.RUQ:Document:Ultrasound
C0881797|Abdomen US
C0881797|Abd US
C0881797|Multisection:Find:Pt:Abdomen:Doc:US
C0881797|Multisection:Finding:Point in time:Abdomen:Document:Ultrasound
C0881957|Head.SS MRI.Angio W contr IV
C0881957|Head Sagittal Sinus MRI angiogram W contrast IV
C0881957|Multisection^W contrast IV:Find:Pt:Head.sagittal sinus:Doc:MRI.angio
C0881957|Multisection^W contrast Intravenous:Finding:Point in time:Head.sagittal sinus:Document:MRI.angio
C0881973|Kidney US Bx guid
C0881973|US Guidance for biopsy of Kidney
C0881973|Guidance for biopsy:Finding:Point in time:Kidney:Document:Ultrasound
C0881973|Guidance for biopsy:Find:Pt:Kidney:Doc:US
C1114484|Sinuses MRI WO contrast
C1114484|Sinuses MRI WO contr
C1114484|Multisection^WO contrast:Finding:Point in time:Sinuses:Document:MRI
C1114484|Multisection^WO contrast:Find:Pt:Sinuses:Doc:MRI
C1114527|Views^W R-bending & W L-bending:Finding:Point in time:Spine:Narrative:XR
C1114527|Spine XR W R+L-bending
C1114527|Spine X-ray W right bending and W left bending
C1114527|Views^W R-bending & W L-bending:Find:Pt:Spine:Doc:XR
C1114527|Views^W R-bending & W L-bending:Finding:Point in time:Spine:Document:XR
C1114578|L-spine XR 1V
C1114578|View 1:Find:Pt:Spine.lumbar:Doc:XR
C1114578|View 1:Finding:Point in time:Spine.lumbar:Document:XR
C1114578|Lumbar spine X-ray Single view
C1114588|Finger fifth X-ray
C1114588|Finger.5th XR
C1114588|Views:Find:Pt:Finger.fifth:Doc:XR
C1114588|Views:Finding:Point in time:Finger.fifth:Document:XR
C1114676|Lower extremity vein US.doppler
C1114676|LE v DOP
C1114676|Multisection:Finding:Point in time:Lower extremity vein:Document:Ultrasound.doppler
C1114676|Multisection:Find:Pt:Lower extremity vein:Doc:US.doppler
C1114417|Multisection^WO & W contrast IV:Find:Pt:Neck:Doc:CT
C1114417|Neck CT WO and W contrast IV
C1114417|Neck CT WO+W contr IV
C1114417|Multisection^WO & W contrast Intravenous:Finding:Point in time:Neck:Document:Computerized Tomography
C1114436|CT Guidance for fine needle aspiration of Kidney - bilateral
C1114436|Guidance for aspiration.fine needle:Finding:Point in time:Kidney.bilateral:Document:Computerized Tomography
C1114436|Guidance for aspiration.fine needle:Find:Pt:Kidney.bilateral:Doc:CT
C1114436|Kdny-Bl CT FNA Asp
C1114441|Pancreas CT WO contr
C1114441|Pancreas CT WO contrast
C1114441|Multisection^WO contrast:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C1114441|Multisection^WO contrast:Find:Pt:Abdomen>Pancreas:Doc:CT
C1543756|Hrt RI PF W Tc99mMIBI IV
C1543756|Heart Scan perfusion W Tc-99m Sestamibi IV
C1543756|Views perfusion^W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543756|Views perfusion^W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543758|Deprecated Views perfusion^W dipyridamole & W 99m Tc mibi IV:Find:Pt:Heart:Nar:Radnuc
C1543758|Views perfusion^W dipyridamole & W 99m Tc mibi IV:Find:Pt:Heart:Nar:Radnuc
C1543758|Deprecated Hrt RI PF
C1543758|Deprecated Heart Scintigraphy perfusion W dipyridamole & W Tc-99m Sestamibi IV
C1543758|Views perfusion^W dipyridamole & W 99m Tc mibi Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1543772|Hrt RI PF Rest+W DPY+Tc99mMIBI IV
C1543772|Heart Scan perfusion at rest and W dipyridamole and W Tc-99m Sestamibi IV
C1543772|Views perfusion^at rest & W dipyridamole & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543772|Views perfusion^at rest & W dipyridamole & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543488|T-spine XR AP 1V W R-bending
C1543488|View AP^W R-bending:Find:Pt:Spine.thoracic:Doc:XR
C1543488|View AP^W R-bending:Finding:Point in time:Spine.thoracic:Document:XR
C1543488|Thoracic spine X-ray AP single view W right bending
C1543490|T-spine XR 4V+Obl
C1543490|Views 4 & oblique:Finding:Point in time:Spine.thoracic:Document:XR
C1543490|Views 4 & oblique:Find:Pt:Spine.thoracic:Doc:XR
C1543490|Thoracic spine X-ray 4 views and oblique
C1543792|Parathyroid SPECT
C1543792|Parathyroid SPECT W RNC IV
C1543792|Multisection^W radionuclide Intravenous:Finding:Point in time:Parathyroid:Document:Radnuc.SPECT
C1543792|Multisection^W radionuclide IV:Find:Pt:Parathyroid:Doc:Radnuc.SPECT
C1543530|Liver Transplant US
C1543530|Multisection:Finding:Point in time:Liver transplant:Document:Ultrasound
C1543530|Multisection:Find:Pt:Liver transplant:Doc:US
C1543578|Ovarian vessels US.doppler
C1543578|Ovarian ves DOP
C1543578|Multisection:Finding:Point in time:Ovarian vessels:Document:Ultrasound.doppler
C1543578|Multisection:Find:Pt:Ovarian vessels:Doc:US.doppler
C1543587|Hip-R XR AP+Danelius Miller
C1543587|Hip - right X-ray AP and Danelius Miller
C1543587|Views AP & Danelius Miller:Finding:Point in time:Hip.right:Document:XR
C1543587|Views AP & Danelius Miller:Find:Pt:Hip.right:Doc:XR
C1525164|Femur - right X-ray tomograph
C1525164|Femur-R XRTomo
C1525164|Multisection:Finding:Point in time:Femur.right:Document:XR.tomo
C1525164|Multisection:Find:Pt:Femur.right:Doc:XR.tomo
C1543681|Pulmonary system Scan
C1543681|Pulm RI W RNC IV
C1543681|Views^W radionuclide Intravenous:Finding:Point in time:Pulmonary system:Document:Radnuc
C1543681|Views^W radionuclide IV:Find:Pt:Pulmonary system:Doc:Radnuc
C1525931|Views ski jump:Finding:Point in time:Calcaneus.right:Document:XR
C1525931|Views ski jump:Find:Pt:Calcaneus.right:Doc:XR
C1525931|Deprecated Heel-R XR Ski Jump
C1525931|Deprecated Calcaneus - right X-ray ski jump
C1526753|Humerus bicipital groove - right X-ray
C1526753|Humerus bicipital groove-R XR
C1526753|Views:Finding:Point in time:Humerus.bicipital groove.right:Document:XR
C1526753|Views:Find:Pt:Humerus.bicipital groove.right:Doc:XR
C1526770|Deprecated Calcaneus - right X-ray Broden
C1526770|Views Broden:Finding:Point in time:Calcaneus.right:Document:XR
C1526770|Views Broden:Find:Pt:Calcaneus.right:Doc:XR
C1526770|Deprecated Heel-R XR Broden
C1526783|Lacrimal duct - right Fluoroscopy W contrast intra lacrimal duct
C1526783|Lacrimal Duct-R Flr W contr intra LD
C1526783|Views^W contrast intra lacrimal duct:Find:Pt:Lacrimal duct.right:Doc:XR.fluor
C1526783|Views^W contrast intra lacrimal duct:Finding:Point in time:Lacrimal duct.right:Document:XR.fluor
C1524827|Chest MRI WO contr
C1524827|Chest MRI WO contrast
C1524827|Multisection^WO contrast:Finding:Point in time:Chest:Document:MRI
C1524827|Multisection^WO contrast:Find:Pt:Chest:Doc:MRI
C1525111|Lower extremity veins - right MRI angiogram
C1525111|LE vv-R MRI.Angio
C1525111|Multisection:Finding:Point in time:Lower extremity veins.right:Document:MRI.angio
C1525111|Multisection:Find:Pt:Lower extremity veins.right:Doc:MRI.angio
C1525115|Pelvis vv MRI.Angio
C1525115|Pelvis veins MRI angiogram
C1525115|Multisection:Finding:Point in time:Pelvis veins:Document:MRI.angio
C1525115|Multisection:Find:Pt:Pelvis veins:Doc:MRI.angio
C1525184|Head vessels MRI angiogram limited
C1525184|Head ves MRI.Angio Ltd
C1525184|Multisection limited:Finding:Point in time:Head vessels:Document:MRI.angio
C1525184|Multisection limited:Find:Pt:Head vessels:Doc:MRI.angio
C1524458|Abdomen CT limited WO contrast
C1524458|Abd CT Ltd WO contr
C1524458|Multisection limited^WO contrast:Find:Pt:Abdomen:Doc:CT
C1524458|Multisection limited^WO contrast:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524235|LE CT Ltd WO contr
C1524235|Lower extremity CT limited WO contrast
C1524235|Multisection limited^WO contrast:Find:Pt:Lower extremity:Doc:CT
C1524235|Multisection limited^WO contrast:Finding:Point in time:Lower extremity:Document:Computerized Tomography
C1525286|Adrenal gland MRI WO contrast
C1525286|Adrenal MRI WO contr
C1525286|Multisection^WO contrast:Find:Pt:Adrenal gland:Doc:MRI
C1525286|Multisection^WO contrast:Finding:Point in time:Adrenal gland:Document:MRI
C1525305|Hip XR Friedman
C1525305|Hip X-ray Friedman
C1525305|View Friedman:Finding:Point in time:Hip:Document:XR
C1525305|View Friedman:Find:Pt:Hip:Doc:XR
C1525208|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen>Renal vessels:Document:Computerized Tomography.angio
C1525208|Multisection^W contrast IV:Find:Pt:Abdomen>Renal vessels:Doc:CT.angio
C1525208|Abd>Renal vls CT.Angio W contr IV
C1525208|Abdominal Renal vessels CT angiogram W contrast IV
C1525230|Multisection^WO & W contrast Intravenous:Finding:Point in time:Carotid vessel:Document:MRI.angio
C1525230|Carotid vessel MRI angiogram WO and W contrast IV
C1525230|Multisection^WO & W contrast IV:Find:Pt:Carotid vessel:Doc:MRI.angio
C1525230|Carot ves MRI.Angio WO+W contr IV
C1525273|Salivary gland CT W contrast intra salivary duct
C1525273|Salivary gland CT W contr intra SD
C1525273|Multisection^W contrast intra salivary duct:Finding:Point in time:Salivary gland:Document:Computerized Tomography
C1525273|Multisection^W contrast intra salivary duct:Find:Pt:Salivary gland:Doc:CT
C1524680|Shoulder - bilateral X-ray outlet
C1524680|Should-Bl XR Outlet
C1524680|View outlet:Find:Pt:Shoulder.bilateral:Doc:XR
C1524680|View outlet:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525492|Should-Bl XR AP+Ax+Outlet
C1525492|Shoulder - bilateral X-ray AP and axillary and outlet
C1525492|Views AP & axillary & outlet:Find:Pt:Shoulder.bilateral:Doc:XR
C1525492|Views AP & axillary & outlet:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525521|Clavicle-L XR AP+Serendipity
C1525521|Clavicle - left X-ray AP and Serendipity
C1525521|Views AP & Serendipity:Find:Pt:Clavicle.left:Doc:XR
C1525521|Views AP & Serendipity:Finding:Point in time:Clavicle.left:Document:XR
C1525540|Chest XR PA+R-Lat
C1525540|Chest X-ray PA and right lateral
C1525540|Views PA & R-lateral:Find:Pt:Chest:Doc:XR
C1525540|Views PA & R-lateral:Finding:Point in time:Chest:Document:XR
C1525622|Temporomandibular joint - bilateral X-ray tomograph
C1525622|TMJ-Bl XRTomo
C1525622|Multisection:Finding:Point in time:Temporomandibular joint.bilateral:Document:XR.tomo
C1525622|Multisection:Find:Pt:Temporomandibular joint.bilateral:Doc:XR.tomo
C1525624|Temporomandibular joint - left X-ray tomograph
C1525624|TMJ-L XRTomo
C1525624|Multisection:Find:Pt:Temporomandibular joint.left:Doc:XR.tomo
C1525624|Multisection:Finding:Point in time:Temporomandibular joint.left:Document:XR.tomo
C1525629|Circle of Willis MRI.Angio
C1525629|Circle of Willis MRI angiogram
C1525629|Multisection:Finding:Point in time:Head+Neck>Circle of Willis:Document:MRI.angio
C1525629|Multisection:Find:Pt:Head+Neck>Circle of Willis:Doc:MRI.angio
C1525647|L-spine+SIJ XR 3V
C1525647|Spine Lumbar and Sacroiliac Joint X-ray 3 views
C1525647|Views 3:Finding:Point in time:Spine.lumbar+Sacroiliac joint:Document:XR
C1525647|Views 3:Find:Pt:Spine.lumbar+Sacroiliac joint:Doc:XR
C1525652|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sternoclavicular joint:Document:Computerized Tomography
C1525652|Multisection^WO & W contrast IV:Find:Pt:Sternoclavicular joint:Doc:CT
C1525652|SC joint CT WO+W contr IV
C1525652|Sternoclavicular Joint CT WO and W contrast IV
C1525705|Ac arch+UE a XRA W contr IA
C1525705|Aortic arch and Upper Extremity artery Fluoroscopic angiogram W contrast IA
C1525705|Views^W contrast IA:Find:Pt:Aortic arch+Upper extremity artery:Doc:XR.fluor.angio
C1525705|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Upper extremity artery:Document:XR.fluor.angio
C1525740|Fem v XRA W contr IV
C1525740|Femoral vein Fluoroscopic angiogram W contrast IV
C1525740|Views^W contrast Intravenous:Finding:Point in time:Femoral vein:Document:XR.fluor.angio
C1525740|Views^W contrast IV:Find:Pt:Femoral vein:Doc:XR.fluor.angio
C1525766|Wrist CT WO contrast
C1525766|Wrist CT WO contr
C1525766|Multisection^WO contrast:Find:Pt:Wrist:Doc:CT
C1525766|Multisection^WO contrast:Finding:Point in time:Wrist:Document:Computerized Tomography
C1525783|Knee X-ray PA W 45 degree flexion
C1525783|Knee XR PA V1 W 45 deg Flx
C1525783|View PA^W 45 degree flexion:Find:Pt:Knee:Doc:XR
C1525783|View PA^W 45 degree flexion:Finding:Point in time:Knee:Document:XR
C1525793|Tibioperon aa XRA W contr IA
C1525793|Tibioperoneal arteries Fluoroscopic angiogram W contrast IA
C1525793|Views^W contrast Intra-arterial:Finding:Point in time:Tibioperoneal arteries:Document:XR.fluor.angio
C1525793|Views^W contrast IA:Find:Pt:Tibioperoneal arteries:Doc:XR.fluor.angio
C1525795|CT Guidance for aspiration of Pleural space
C1525795|Pl space CT Asp guid
C1525795|Guidance for aspiration:Find:Pt:Chest>Pleural space:Doc:CT
C1525795|Guidance for aspiration:Finding:Point in time:Chest>Pleural space:Document:Computerized Tomography
C1525862|Unspecified body region Fluoroscopy W contrast via catheter
C1525862|XXX Flr W contr via cath
C1525862|Views^W contrast via catheter:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1525862|Views^W contrast via catheter:Find:Pt:XXX:Doc:XR.fluor
C1525880|Great toe-L XR stand
C1525880|Great toe - left X-ray standing
C1525880|Views^standing:Find:Pt:Great toe.left:Doc:XR
C1525880|Views^standing:Finding:Point in time:Great toe.left:Document:XR
C1525882|Penis Fluoroscopy W contrast intra corpus cavernosum
C1525882|Penis Flr W contr intra CC
C1525882|Views^W contrast intra corpus cavernosum:Finding:Point in time:Penis:Document:XR.fluor
C1525882|Views^W contrast intra corpus cavernosum:Find:Pt:Penis:Doc:XR.fluor
C1524144|Lymph Pelvic-Bl Flr W contr IL
C1524144|Lymphatics pelvic - bilateral Fluoroscopy W contrast intra lymphatic
C1524144|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.pelvic.bilateral:Document:XR.fluor
C1524144|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.pelvic.bilateral:Doc:XR.fluor
C1525889|Nasal bones XR Lat+Waters
C1525889|Nasal bones X-ray lateral and Waters
C1525889|Views lateral & Waters:Find:Pt:Nasal bones:Doc:XR
C1525889|Views lateral & Waters:Finding:Point in time:Nasal bones:Document:XR
C1525942|Pelvis XR AP+Lat+Obl
C1525942|Pelvis X-ray AP and lateral and oblique
C1525942|Views AP & lateral & oblique:Find:Pt:Pelvis:Doc:XR
C1525942|Views AP & lateral & oblique:Finding:Point in time:Pelvis:Document:XR
C1525812|L-spine CT W contr ID
C1525812|Multisection^W contrast intradisc:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1525812|Multisection^W contrast intradisc:Find:Pt:Spine.lumbar:Doc:CT
C1525812|Lumbar spine CT W contrast intradisc
C1525813|Spine ves MRI.Angio WO contr
C1525813|Spine vessels MRI angiogram WO contrast
C1525813|Multisection^WO contrast:Finding:Point in time:Spine vessels:Document:MRI.angio
C1525813|Multisection^WO contrast:Find:Pt:Spine vessels:Doc:MRI.angio
C1525975|T+L-spine XR Scoli AP 1V stand
C1525975|View scoliosis AP^standing:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1525975|View scoliosis AP^standing:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1525975|Spine Thoracic and Lumbar X-ray scoliosis AP standing
C1526021|Ft-R XR W Stress
C1526021|Foot - right X-ray W manual stress
C1526021|Views^W manual stress:Finding:Point in time:Foot.right:Document:XR
C1526021|Views^W manual stress:Find:Pt:Foot.right:Doc:XR
C1526105|Shoulder - right X-ray axillary
C1526105|Should-R XR Ax
C1526105|View axillary:Finding:Point in time:Shoulder.right:Document:XR
C1526105|View axillary:Find:Pt:Shoulder.right:Doc:XR
C1526126|Toes - right X-ray 2 views
C1526126|Toes-R XR 2V
C1526126|Views 2:Finding:Point in time:Toes.right:Document:XR
C1526126|Views 2:Find:Pt:Toes.right:Doc:XR
C1525905|Wrist-R XR PA+Lat
C1525905|Wrist - right X-ray PA and lateral
C1525905|Views PA & lateral:Finding:Point in time:Wrist.right:Document:XR
C1525905|Views PA & lateral:Find:Pt:Wrist.right:Doc:XR
C1526084|Brst-R Mam 2V
C1526084|Breast - right Mammogram 2 views
C1526084|Views 2:Find:Pt:Breast.right:Doc:Mam
C1526084|Views 2:Finding:Point in time:Breast.right:Document:Mam
C1526183|T-spine XR Lat Xtable
C1526183|View lateral crosstable:Find:Pt:Spine.thoracic:Doc:XR
C1526183|View lateral crosstable:Finding:Point in time:Spine.thoracic:Document:XR
C1526183|Thoracic spine X-ray lateral crosstable
C1526196|US Guidance for needle biopsy of Lymph node
C1526196|LN US Bx needle guid
C1526196|Guidance for biopsy.needle:Find:Pt:Lymph node:Doc:US
C1526196|Guidance for biopsy.needle:Finding:Point in time:Lymph node:Document:Ultrasound
C1526204|Zygomatic arch XR 4V
C1526204|Zygomatic arch X-ray 4 views
C1526204|Views 4:Find:Pt:Zygomatic arch:Doc:XR
C1526204|Views 4:Finding:Point in time:Zygomatic arch:Document:XR
C1526240|Spine thoracolumbar junction XR
C1526240|Spine Thoracolumbar Junction X-ray
C1526240|Views:Find:Pt:Spine.thoracolumbar junction:Doc:XR
C1526240|Views:Finding:Point in time:Spine.thoracolumbar junction:Document:XR
C1526256|Views Grashey^WO & W weight:Find:Pt:Shoulder.left:Doc:XR
C1526256|Should-L XR Grashey WO+W Wt
C1526256|Shoulder - left X-ray Grashey WO and W weight
C1526256|Views Grashey^WO & W weight:Finding:Point in time:Shoulder.left:Document:XR
C1526279|Pelvis US limited
C1526279|Pelvis US Ltd
C1526279|Multisection limited:Find:Pt:Pelvis:Doc:US
C1526279|Multisection limited:Finding:Point in time:Pelvis:Document:Ultrasound
C1524478|Abd MRI W contr IV
C1524478|Abdomen MRI W contrast IV
C1524478|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen:Document:MRI
C1524478|Multisection^W contrast IV:Find:Pt:Abdomen:Doc:MRI
C1524506|Elbow-R MRI W contr IV
C1524506|Elbow - right MRI W contrast IV
C1524506|Multisection^W contrast IV:Find:Pt:Elbow.right:Doc:MRI
C1524506|Multisection^W contrast Intravenous:Finding:Point in time:Elbow.right:Document:MRI
C1524884|LE.joint-R MRI WO contr
C1524884|Lower extremity joint - right MRI WO contrast
C1524884|Multisection^WO contrast:Finding:Point in time:Lower extremity.joint.right:Document:MRI
C1524884|Multisection^WO contrast:Find:Pt:Lower extremity.joint.right:Doc:MRI
C1524526|Ft-L MRI W contr IV
C1524526|Foot - left MRI W contrast IV
C1524526|Multisection^W contrast IV:Find:Pt:Foot.left:Doc:MRI
C1524526|Multisection^W contrast Intravenous:Finding:Point in time:Foot.left:Document:MRI
C1524146|Sacrum+Coccyx MRI WO contr
C1524146|Sacrum and Coccyx MRI WO contrast
C1524146|Multisection^WO contrast:Finding:Point in time:Sacrum+Coccyx:Document:MRI
C1524146|Multisection^WO contrast:Find:Pt:Sacrum+Coccyx:Doc:MRI
C1524148|Should CT WO contr
C1524148|Shoulder CT WO contrast
C1524148|Multisection^WO contrast:Finding:Point in time:Shoulder:Document:Computerized Tomography
C1524148|Multisection^WO contrast:Find:Pt:Shoulder:Doc:CT
C1524583|Scapula-R MRI W contr IV
C1524583|Scapula - right MRI W contrast IV
C1524583|Multisection^W contrast Intravenous:Finding:Point in time:Scapula.right:Document:MRI
C1524583|Multisection^W contrast IV:Find:Pt:Scapula.right:Doc:MRI
C1524937|View 1:Find:Pt:Calcaneus:Doc:XR
C1524937|Deprecated Calcaneus X-ray Single view
C1524937|Deprecated Heel XR 1V
C1524937|View 1:Finding:Point in time:Calcaneus:Document:XR
C1524592|Lower leg CT W contr IV
C1524592|Lower leg CT W contrast IV
C1524592|Multisection^W contrast IV:Find:Pt:Lower leg:Doc:CT
C1524592|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg:Document:Computerized Tomography
C1524628|Femur XR 3V
C1524628|Femur X-ray 3 views
C1524628|Views 3:Finding:Point in time:Femur:Document:XR
C1524628|Views 3:Find:Pt:Femur:Doc:XR
C1524634|Hip - bilateral X-ray 3 views
C1524634|Hip-Bl XR 3V
C1524634|Views 3:Find:Pt:Hip.bilateral:Doc:XR
C1524634|Views 3:Finding:Point in time:Hip.bilateral:Document:XR
C1524635|Hip-L XR 3V
C1524635|Hip - left X-ray 3 views
C1524635|Views 3:Find:Pt:Hip.left:Doc:XR
C1524635|Views 3:Finding:Point in time:Hip.left:Document:XR
C1525006|Shoulder - bilateral X-ray 2 views
C1525006|Should-Bl XR 2V
C1525006|Views 2:Find:Pt:Shoulder.bilateral:Doc:XR
C1525006|Views 2:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525019|C-spine XR 7V
C1525019|Views 7:Find:Pt:Spine.cervical:Doc:XR
C1525019|Views 7:Finding:Point in time:Spine.cervical:Document:XR
C1525019|Cervical spine X-ray 7 views
C1525067|Ft XR AP+Lat+Obl
C1525067|Foot X-ray AP and lateral and oblique
C1525067|Views AP & lateral & oblique:Find:Pt:Foot:Doc:XR
C1525067|Views AP & lateral & oblique:Finding:Point in time:Foot:Document:XR
C1830191|CT Guidance for biopsy of Unspecified body region-- WO contrast
C1830191|XXX CT Bx guid WO contr
C1830191|Guidance for biopsy^WO contrast:Find:Pt:XXX:Doc:CT
C1830191|Guidance for biopsy^WO contrast:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1830239|Breast - unilateral Mammogram Single view
C1830239|Brst-UL Mam 1V
C1830239|View 1:Finding:Point in time:Breast.unilateral:Document:Mam
C1830239|View 1:Find:Pt:Breast.unilateral:Doc:Mam
C1830246|Elbow - right X-ray GE 3 views
C1830246|Elbow-R XR GE 3V
C1830246|Views GE 3:Find:Pt:Elbow.right:Doc:XR
C1830246|Views GE 3:Finding:Point in time:Elbow.right:Document:XR
C1830257|Breast - unilateral Mammogram screening
C1830257|Brst-UL Mam Screening
C1830257|Views screening:Find:Pt:Breast.unilateral:Doc:Mam
C1830257|Views screening:Finding:Point in time:Breast.unilateral:Document:Mam
C1830074|Mandible X-ray LE 3 views
C1830074|Mandible XR LE 3V
C1830074|Views LE 3:Finding:Point in time:Mandible:Document:XR
C1830074|Views LE 3:Find:Pt:Mandible:Doc:XR
C1715409|PET WB
C1715409|PET whole body
C1715409|Multisection whole body:Finding:Point in time:^Patient:Document:Radnuc.PET
C1715409|Multisection whole body:Find:Pt:^Patient:Doc:Radnuc.PET
C1715435|Guidance for drainage of abscess:Finding:Point in time:Peritoneal space:Document:Ultrasound
C1715435|Peritoneal space US Abscess drain guid
C1715435|Guidance for drainage of abscess:Find:Pt:Peritoneal space:Doc:US
C1715435|US Guidance for drainage of abscess of Peritoneal space
C1715452|C-spine XR AP+Obl+Odont+Lat Port W FE
C1715452|Views AP & oblique & odontoid & lateral portable^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C1715452|Views AP & oblique & odontoid & lateral portable^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C1715452|Cervical spine X-ray AP and oblique and odontoid and lateral portable W flexion and W extension
C1715460|Knee - bilateral X-ray GE 5 views standing
C1715460|Knee-Bl XR GE 5V stand
C1715460|Views GE 5^standing:Finding:Point in time:Knee.bilateral:Document:XR
C1715460|Views GE 5^standing:Find:Pt:Knee.bilateral:Doc:XR
C1715461|Knee XR 1V or 2V
C1715461|Knee X-ray 1 or 2 views
C1715461|Views 1 or 2:Find:Pt:Knee:Doc:XR
C1715461|Views 1 or 2:Finding:Point in time:Knee:Document:XR
C1715462|Face XR 1V or 2V
C1715462|Facial bones X-ray 1 or 2 views
C1715462|Views 1 or 2:Finding:Point in time:Facial bones:Document:XR
C1715462|Views 1 or 2:Find:Pt:Facial bones:Doc:XR
C1715464|Pelvis X-ray 1 or 2 views portable
C1715464|Pelvis XR 1V or 2V Port
C1715464|Views 1 or 2 portable:Finding:Point in time:Pelvis:Document:XR
C1715464|Views 1 or 2 portable:Find:Pt:Pelvis:Doc:XR
C1715486|Colon Flr Reduction W views W Ba PR
C1715486|Colon Fluoroscopy Reduction W views W barium contrast PR
C1715486|Reduction W views^W barium contrast PR:Find:Pt:Colon:Doc:XR.fluor
C1715486|Reduction W views^W barium contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C1717322|Multisection^WO & W contrast IV:Find:Pt:Superior mesenteric vessels:Doc:MRI.angio
C1717322|Superior mesenteric vessels MRI angiogram WO and W contrast IV
C1717322|Multisection^WO & W contrast Intravenous:Finding:Point in time:Superior mesenteric vessels:Document:MRI.angio
C1717322|SM ves MRI.Angio WO+W contr IV
C1644648|Humerus - left X-ray portable
C1644648|Humerus-L XR port
C1644648|Views portable:Find:Pt:Humerus.left:Doc:XR
C1644648|Views portable:Finding:Point in time:Humerus.left:Document:XR
C1643600|Extr vv-L US
C1643600|Extremity veins - left US
C1643600|Multisection:Finding:Point in time:Extremity veins.left:Document:Ultrasound
C1643600|Multisection:Find:Pt:Extremity veins.left:Doc:US
C1625228|AV shunt RI W RNC IV
C1625228|AV shunt Scan
C1625228|Views^W radionuclide IV:Find:Pt:AV shunt:Doc:Radnuc
C1625228|Views^W radionuclide Intravenous:Finding:Point in time:AV shunt:Document:Radnuc
C1714527|Guidance for localization of bleeding site^W radionuclide Intravenous:Finding:Point in time:^Patient:Narrative:Radnuc
C1714527|Deprecated RI Bleeding local guid W RNC
C1714527|Deprecated Scan Guidance for localization of bleeding site
C1714527|Guidance for localization of bleeding site^W radionuclide IV:Find:Pt:^Patient:Nar:Radnuc
C1714931|Chest and Abdomen X-ray upright and PA chest
C1714931|Chest+Abd XR upright+PA chst
C1714931|Views upright & PA chest:Finding:Point in time:Chest+Abdomen:Document:XR
C1714931|Views upright & PA chest:Find:Pt:Chest+Abdomen:Doc:XR
C1715021|RI for ETr Mul Areas W In-111-P IV
C1715021|Scan for endocrine tumor multiple areas W In-111 pentetreotide IV
C1715021|Views for endocrine tumor multiple areas^W In-111 pentetreotide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1715021|Views for endocrine tumor multiple areas^W In-111 pentetreotide IV:Find:Pt:^Patient:Doc:Radnuc
C1715022|Liver+BDs+GB RI W CCK+RNC IV
C1715022|Liver and Biliary ducts and Gallbladder Scan W cholecystokinin and W radionuclide IV
C1715022|Views^W cholecystokinin & W radionuclide Intravenous:Finding:Point in time:Liver+Biliary ducts+Gallbladder:Document:Radnuc
C1715022|Views^W cholecystokinin & W radionuclide IV:Find:Pt:Liver+Biliary ducts+Gallbladder:Doc:Radnuc
C1639942|L-spine XR W R+L-bending
C1639942|Views^W R-bending & W L-bending:Finding:Point in time:Spine.lumbar:Document:XR
C1639942|Views^W R-bending & W L-bending:Find:Pt:Spine.lumbar:Doc:XR
C1639942|Lumbar spine X-ray W right bending and W left bending
C1624109|Views^W non-ionic contrast IT:Find:Pt:Spine.cervical:Nar:XR.fluor
C1624109|Deprecated C-spine Flr W Non-ionic contr
C1624109|Deprecated Spine Cervical X-ray fluoroscopy W contrast IT
C1624109|Views^W non-ionic contrast Intrathecal:Finding:Point in time:Spine.cervical:Narrative:XR.fluor
C1632785|Views^W non-ionic contrast IT:Find:Pt:Spine.thoracic:Nar:XR.fluor
C1632785|Deprecated T-spine Flr W Non-ionic contr
C1632785|Deprecated Spine Thoracic X-ray fluoroscopy W contrast IT
C1632785|Views^W non-ionic contrast Intrathecal:Finding:Point in time:Spine.thoracic:Narrative:XR.fluor
C1636072|US Guidance for aspiration of cyst of Breast - left
C1636072|Brst-L US Cyst Asp guid
C1636072|Guidance for aspiration of cyst:Finding:Point in time:Breast.left:Document:Ultrasound
C1636072|Guidance for aspiration of cyst:Find:Pt:Breast.left:Doc:US
C1631256|Views:Finding:Point in time:Abdomen+Chest:Narrative:XR
C1631256|Chest+Abd XR
C1631256|Chest and Abdomen X-ray
C1631256|Views:Find:Pt:Chest+Abdomen:Doc:XR
C1631256|Views:Finding:Point in time:Chest+Abdomen:Document:XR
C1633469|Prostate US Drain guid
C1633469|US Guidance for drainage of Prostate
C1633469|Guidance for drainage:Finding:Point in time:Prostate:Document:Ultrasound
C1633469|Guidance for drainage:Find:Pt:Prostate:Doc:US
C1953940|Kidney US Asp guid
C1953940|US Guidance for aspiration of Kidney
C1953940|Guidance for aspiration:Find:Pt:Kidney:Doc:US
C1953940|Guidance for aspiration:Finding:Point in time:Kidney:Document:Ultrasound
C3533790|Views for motility^W radioopaque markers:Find:Pt:Abdomen:Doc:XR
C3533790|Abd XR for Motility W ROMS
C3533790|Views for motility^W radioopaque markers:Finding:Point in time:Abdomen:Document:XR
C3533790|Abdomen X-ray for motility W radioopaque markers
C3262937|Multisection^W contrast IS:Find:Pt:Knee.right:Doc:CT
C3262937|Knee - right CT W contrast IS
C3262937|Knee-R CT W contr IS
C3262937|Multisection^W contrast Intrasynovial:Finding:Point in time:Knee.right:Document:Computerized Tomography
C3262941|Scapula CT WO contr
C3262941|Scapula CT WO contrast
C3262941|Multisection^WO contrast:Finding:Point in time:Scapula:Document:Computerized Tomography
C3262941|Multisection^WO contrast:Find:Pt:Scapula:Doc:CT
C3262944|Fluoroscopy Guidance for aspiration of cyst of Ovary
C3262944|Ovary Flr Cyst Asp guid
C3262944|Guidance for aspiration of cyst:Find:Pt:Ovary:Doc:XR.fluor
C3262944|Guidance for aspiration of cyst:Finding:Point in time:Ovary:Document:XR.fluor
C3262959|Ankle - left X-ray AP and lateral and oblique standing
C3262959|Ankle-L XR AP+Lat+Obl stand
C3262959|Views AP & lateral & oblique^standing:Find:Pt:Ankle.left:Doc:XR
C3262959|Views AP & lateral & oblique^standing:Finding:Point in time:Ankle.left:Document:XR
C3262998|Hand-Bl MRI W contr IV
C3262998|Hand - bilateral MRI W contrast IV
C3262998|Multisection^W contrast Intravenous:Finding:Point in time:Hand.bilateral:Document:MRI
C3262998|Multisection^W contrast IV:Find:Pt:Hand.bilateral:Doc:MRI
C3263101|Upper extremity vein Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IV
C3263101|UE v XRA PTA of ves W contr IV
C3263101|Percutaneous transluminal angioplasty of vessel^W contrast Intravenous:Finding:Point in time:Upper extremity vein:Document:XR.fluor.angio
C3263101|Percutaneous transluminal angioplasty of vessel^W contrast IV:Find:Pt:Upper extremity vein:Doc:XR.fluor.angio
C3263214|Breast v DOP
C3263214|Breast vessels US.doppler
C3263214|Multisection:Find:Pt:Breast vessels:Doc:US.doppler
C3263214|Multisection:Finding:Point in time:Breast vessels:Document:Ultrasound.doppler
C3262914|Wrist-Bl CT W contr IV
C3262914|Wrist - bilateral CT W contrast IV
C3262914|Multisection^W contrast Intravenous:Finding:Point in time:Wrist.bilateral:Document:Computerized Tomography
C3262914|Multisection^W contrast IV:Find:Pt:Wrist.bilateral:Doc:CT
C0942206|Multisection^WO & W contrast IV:Find:Pt:Shoulder.bilateral:Doc:MRI
C0942206|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder.bilateral:Document:MRI
C0942206|Should-Bl MRI WO+W contr IV
C0942206|Shoulder - bilateral MRI WO and W contrast IV
C0942268|Multisection:Finding:Point in time:Thigh.bilateral:Narrative:MRI
C0942268|Thigh - bilateral MRI
C0942268|Thigh-Bl MRI
C0942268|Multisection:Find:Pt:Thigh.bilateral:Doc:MRI
C0942268|Multisection:Finding:Point in time:Thigh.bilateral:Document:MRI
C0945327|Foot - left MRI
C0945327|Ft-L MRI
C0945327|Multisection:Finding:Point in time:Foot.left:Document:MRI
C0945327|Multisection:Find:Pt:Foot.left:Doc:MRI
C0942310|Spine facet joint-L Flr Inj guid
C0942310|Fluoroscopy Guidance for injection of Spine facet joint - left
C0942310|Guidance for injection:Finding:Point in time:Spine facet joint.left:Document:XR.fluor
C0942310|Guidance for injection:Find:Pt:Spine facet joint.left:Doc:XR.fluor
C0942359|Hand - left X-ray 3 views
C0942359|Hand-L XR 3V
C0942359|Views 3:Find:Pt:Hand.left:Doc:XR
C0942359|Views 3:Finding:Point in time:Hand.left:Document:XR
C0882052|Pancreas US
C0882052|Multisection:Find:Pt:Pancreas:Doc:US
C0882052|Multisection:Finding:Point in time:Pancreas:Document:Ultrasound
C0882119|C-spine XR 1V
C0882119|View 1:Finding:Point in time:Spine.cervical:Narrative:XR
C0882119|View 1:Finding:Point in time:Spine.cervical:Document:XR
C0882119|View 1:Find:Pt:Spine.cervical:Doc:XR
C0882119|Cervical spine X-ray Single view
C0882169|Tib+Fib XR
C0882169|Tibia and Fibula X-ray
C0882169|Views:Finding:Point in time:Tibia+Fibula:Narrative:XR
C0882169|Views:Finding:Point in time:Tibia+Fibula:Document:XR
C0882169|Views:Find:Pt:Tibia+Fibula:Doc:XR
C0882184|Fluoroscopic angiogram Guidance for placement of catheter for adminstration of thrombolytic in Vessel-- W contrast intravascular
C0882184|Guidance for placement of catheter for adminstration of thrombolytic^W contrast intravascular:Find:Pt:Vessel:Doc:XR.fluor.angio
C0882184|Guidance for placement of catheter for adminstration of thrombolytic^W contrast intravascular:Finding:Point in time:Vessel:Document:XR.fluor.angio
C0882184|Vesl XRA Cath plac gd Tl admn W contr IV
C2709246|Deprecated Views:Finding:Point in time:Wrist:Narrative:XR
C2709246|Views:Find:Pt:Wrist:Nar:XR
C2709246|Deprecated Wrist X-ray
C2709246|Deprecated Wrist XR
C2709246|Views:Finding:Point in time:Wrist:Narrative:XR
C0882199|CT Guidance for aspiration of Unspecified body region
C0882199|XXX CT Asp guid
C0882199|Guidance for aspiration:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882199|Guidance for aspiration:Find:Pt:XXX:Doc:CT
C0942094|Hip - left Fluoroscopy W contrast IS
C0942094|Views^W contrast IS:Find:Pt:Hip.left:Doc:XR.fluor
C0942094|Views^W contrast Intrasynovial:Finding:Point in time:Hip.left:Document:XR.fluor
C0942094|Hip-L Flr W contr IS
C0942128|Elbow-Bl XR
C0942128|Elbow - bilateral X-ray
C0942128|Views:Finding:Point in time:Elbow.bilateral:Document:XR
C0942128|Views:Find:Pt:Elbow.bilateral:Doc:XR
C0942136|Femur-L XR
C0942136|Femur - left X-ray
C0942136|Views:Find:Pt:Femur.left:Doc:XR
C0942136|Views:Finding:Point in time:Femur.left:Document:XR
C0942138|Femur - right X-ray
C0942138|Femur-R XR
C0942138|Views:Find:Pt:Femur.right:Doc:XR
C0942138|Views:Finding:Point in time:Femur.right:Document:XR
C0942143|Hip - bilateral X-ray
C0942143|Hip-Bl XR
C0942143|Views:Find:Pt:Hip.bilateral:Doc:XR
C0942143|Views:Finding:Point in time:Hip.bilateral:Document:XR
C0881778|US Guidance for removal of amniotic fluid from Uterus
C0881778|Uterus US Amn fld rem guid
C0881778|Guidance for removal of amniotic fluid:Finding:Point in time:Uterus:Document:Ultrasound
C0881778|Guidance for removal of amniotic fluid:Find:Pt:Uterus:Doc:US
C0881876|Chest XR AP (R+L-Lat Decub) Port
C0881876|Chest X-ray AP (right lateral-decubitus and left lateral-decubitus) portable
C0881876|Views AP (R-lateral-decubitus & L-lateral-decubitus) portable:Find:Pt:Chest:Doc:XR
C0881876|Views AP (R-lateral-decubitus & L-lateral-decubitus) portable:Finding:Point in time:Chest:Document:XR
C0881908|Esoph+Stom RI W Tc99mSC PO
C0881908|Esophagus and Stomach Scan W Tc-99m SC PO
C0881908|Views^W Tc-99m SC PO:Find:Pt:Esophagus+Stomach:Doc:Radnuc
C0881908|Views^W Tc-99m Subcutaneous Oral:Finding:Point in time:Esophagus+Stomach:Document:Radnuc
C0881920|Fem a XRA Angpsty W contr IA
C0881920|Femoral artery Fluoroscopic angiogram Angioplasty W contrast IA
C0881920|Angioplasty^W contrast IA:Find:Pt:Femoral artery:Doc:XR.fluor.angio
C0881920|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Femoral artery:Document:XR.fluor.angio
C0881922|Femur+Tib XR Leg Length
C0881922|Femur and Tibia X-ray for leg length
C0881922|Views for leg length:Finding:Point in time:Femur+Tibia:Document:XR
C0881922|Views for leg length:Find:Pt:Femur+Tibia:Doc:XR
C0881926|Multisection:Finding:Point in time:Finger:Narrative:MRI
C0881926|Finger MRI
C0881926|Multisection:Find:Pt:Finger:Doc:MRI
C0881926|Multisection:Finding:Point in time:Finger:Document:MRI
C0881938|Groin US
C0881938|Multisection:Find:Pt:Groin:Doc:US
C0881938|Multisection:Finding:Point in time:Groin:Document:Ultrasound
C0881939|Hand MRI
C0881939|Multisection:Finding:Point in time:Hand:Document:MRI
C0881939|Multisection:Find:Pt:Hand:Doc:MRI
C0881940|Hand X-ray 3 views
C0881940|Hand XR 3V
C0881940|Views 3:Find:Pt:Hand:Doc:XR
C0881940|Views 3:Finding:Point in time:Hand:Document:XR
C0881949|Head US
C0881949|Multisection:Finding:Point in time:Head:Document:Ultrasound
C0881949|Multisection:Find:Pt:Head:Doc:US
C0881991|MULTISECTION:FINDING:POINT IN TIME:KIDNEY.BILATERAL AND COLLECTING SYSTEM:NARRATIVE:XR.TOMO
C0881991|Deprecated KD-Bl+CS XR.Tomo
C0881991|Deprecated Kidney Bilateral & Collecting system X-ray tomograph Multisection
C0881991|Multisection:Find:Pt:Kidney.bilateral+Collecting system:Nar:XR.tomo
C0881991|Multisection:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:XR.tomo
C0882004|Knee XR AP+Lat stand
C0882004|Knee X-ray AP and lateral standing
C0882004|Views AP & lateral^standing:Find:Pt:Knee:Doc:XR
C0882004|Views AP & lateral^standing:Finding:Point in time:Knee:Document:XR
C1114933|Multisection^WO & W contrast IV:Find:Pt:Foot:Doc:MRI
C1114933|Foot MRI WO and W contrast IV
C1114933|Multisection^WO & W contrast Intravenous:Finding:Point in time:Foot:Document:MRI
C1114933|Ft MRI WO+W contr IV
C1114935|Should MRI WO contr
C1114935|Shoulder MRI WO contrast
C1114935|Multisection^WO contrast:Finding:Point in time:Shoulder:Document:MRI
C1114935|Multisection^WO contrast:Find:Pt:Shoulder:Doc:MRI
C1114512|Thyroid RI +Single Uptake W RNC IV
C1114512|Thyroid Scan and uptake.single
C1114512|Views & uptake.single^W radionuclide IV:Find:Pt:Thyroid:Doc:Radnuc
C1114512|Views & uptake.single^W radionuclide Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1114595|Knee X-ray tunnel
C1114595|Knee XR V1 Tunnel
C1114595|View tunnel:Finding:Point in time:Knee:Document:XR
C1114595|View tunnel:Find:Pt:Knee:Doc:XR
C1114627|SS v XRA W contr IV
C1114627|Sagittal sinus vein Fluoroscopic angiogram W contrast IV
C1114627|Views^W contrast Intravenous:Finding:Point in time:Sagittal sinus vein:Document:XR.fluor.angio
C1114627|Views^W contrast IV:Find:Pt:Sagittal sinus vein:Doc:XR.fluor.angio
C1114423|Multisection^WO & W contrast IV:Find:Pt:Neck>Vessels:Doc:CT.angio
C1114423|Multisection^WO & W contrast Intravenous:Finding:Point in time:Neck>Vessels:Document:Computerized Tomography.angio
C1114423|Neck ves CT.Angio WO+W contr IV
C1114423|Neck vessels CT angiogram WO and W contrast IV
C1114445|Multisection^WO contrast:Find:Pt:Kidney.bilateral+Collecting system:Nar:CT
C1114445|Multisection^WO contrast:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:Computerized Tomography
C1114445|Deprecated Kidney - bilateral and Collecting system CT WO contrast
C1114445|Deprecated KD-Bl+CS CT WO contr
C1114459|Esoph Flr W Ba PO
C1114459|Esophagus Fluoroscopy W barium contrast PO
C1114459|Views^W barium contrast PO:Find:Pt:Esophagus:Doc:XR.fluor
C1114459|Views^W barium contrast Oral:Finding:Point in time:Esophagus:Document:XR.fluor
C1114459|VIEWS^W BARIUM CONTRAST ORAL:FINDING:POINT IN TIME:ESOPHAGUS:NARRATIVE:XR.FLUOR
C1543444|Kidney - bilateral X-ray tomograph WO contrast
C1543444|Multisection^WO contrast:Find:Pt:Kidney.bilateral:Doc:XR.tomo
C1543444|Multisection^WO contrast:Finding:Point in time:Kidney.bilateral:Document:XR.tomo
C1543444|Kdny-Bl XRTomo WO contr
C1543454|Ankle-R XR & (view W Stress)
C1543454|Ankle - right X-ray and (view W manual stress)
C1543454|Views & (view^W manual stress):Find:Pt:Ankle.right:Doc:XR
C1543454|Views & (view^W manual stress):Finding:Point in time:Ankle.right:Document:XR
C1543757|Hrt RI PF W DIPY+Tc99mMIBI IV
C1543757|Heart Scan perfusion W dipyridamole and W Tc-99m Sestamibi IV
C1543757|Views perfusion^W dipyridamole & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543757|Views perfusion^W dipyridamole & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543467|Knee-R XR 4V+Sunrise+Tunnel
C1543467|Knee - right X-ray 4 views and Sunrise and tunnel
C1543467|Views 4 & Sunrise & tunnel:Finding:Point in time:Knee.right:Document:XR
C1543467|Views 4 & Sunrise & tunnel:Find:Pt:Knee.right:Doc:XR
C1542924|Hrt RI FP W Stress+W RNC IV
C1542924|Heart Scan first pass W stress and W radionuclide IV
C1542924|Views first pass^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1542924|Views first pass^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543913|Hrt RI for Infarct+FP W Tc99mPyp IV
C1543913|Heart Scan for infarct and first pass W Tc-99m PYP IV
C1543913|Views for infarct & first pass^W Tc-99m PYP IV:Find:Pt:Heart:Doc:Radnuc
C1543913|Views for infarct & first pass^W Tc-99m PYP Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543920|Lung SPECT ventilation W radionuclide aerosol IH
C1543920|Lung SPECT V W RNC Aero IH
C1543920|Multisection ventilation^W radionuclide aerosol IH:Find:Pt:Lung:Doc:Radnuc.SPECT
C1543920|Multisection ventilation^W radionuclide aerosol Inhalation:Finding:Point in time:Lung:Document:Radnuc.SPECT
C1543151|Vein - bilateral US
C1543151|Vein-Bl US
C1543151|Multisection:Find:Pt:Vein.bilateral:Doc:US
C1543151|Multisection:Finding:Point in time:Vein.bilateral:Document:Ultrasound
C1543164|Multisection & 3D reconstruction:Find:Pt:XXX:Doc:MRI
C1543164|Multisection & 3D reconstruction:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1543164|Deprecated XXX MRI +3DR
C1543164|Deprecated Unspecified body region MRI and 3D reconstruction
C1543180|UGI Flr W Air+Ba PO
C1543180|Gastrointestine upper Fluoroscopy W air and barium contrast PO
C1543180|Views^W air & barium contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1543180|Views^W air & barium contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1543193|Ankle XR AP+Lat+Obl
C1543193|Ankle X-ray AP and lateral and oblique
C1543193|Views AP & lateral & oblique:Find:Pt:Ankle:Doc:XR
C1543193|Views AP & lateral & oblique:Finding:Point in time:Ankle:Document:XR
C1543259|Fluoroscopic angiogram Guidance for vascular access of Vessel
C1543259|Guidance for vascular access:Finding:Point in time:Vessel:Document:XR.fluor.angio
C1543259|Guidance for vascular access:Find:Pt:Vessel:Doc:XR.fluor.angio
C1543259|Vesl XRA VA guid
C1543267|Breast duct - bilateral Mammogram W contrast intra multiple ducts
C1543267|Brst.duct-Bl Mam W contr intra Dcts
C1543267|Views^W contrast intra multiple ducts:Find:Pt:Breast.duct.bilateral:Doc:Mam
C1543267|Views^W contrast intra multiple ducts:Finding:Point in time:Breast.duct.bilateral:Document:Mam
C1543684|SPECT Abscess local guid WB W RNC IV
C1543684|SPECT Guidance for abscess localization whole body
C1543684|Guidance for abscess localization whole body^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543684|Guidance for abscess localization whole body^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1524259|Pelvis+Hip-R XR AP+Lat Xtable
C1524259|Pelvis and Hip - right X-ray AP and lateral crosstable
C1524259|Views AP & lateral crosstable:Find:Pt:Pelvis+Hip.right:Doc:XR
C1524259|Views AP & lateral crosstable:Finding:Point in time:Pelvis+Hip.right:Document:XR
C1526771|Foot - right X-ray AP standing
C1526771|Ft-R XR AP stand
C1526771|Views AP^standing:Finding:Point in time:Foot.right:Document:XR
C1526771|Views AP^standing:Find:Pt:Foot.right:Doc:XR
C1543706|Breast SPECT
C1543706|Brst SPECT W RNC IV
C1543706|Multisection^W radionuclide IV:Find:Pt:Breast:Doc:Radnuc.SPECT
C1543706|Multisection^W radionuclide Intravenous:Finding:Point in time:Breast:Document:Radnuc.SPECT
C1543707|Breast Scan limited
C1543707|Brst RI Ltd W RNC IV
C1543707|Views limited^W radionuclide Intravenous:Finding:Point in time:Breast:Document:Radnuc
C1543707|Views limited^W radionuclide IV:Find:Pt:Breast:Doc:Radnuc
C1526786|Should-L MRI W contr IV
C1526786|Shoulder - left MRI W contrast IV
C1526786|Multisection^W contrast Intravenous:Finding:Point in time:Shoulder.left:Document:MRI
C1526786|Multisection^W contrast IV:Find:Pt:Shoulder.left:Doc:MRI
C1526797|Ankle-L XR 2V stand
C1526797|Ankle - left X-ray 2 views standing
C1526797|Views 2^standing:Find:Pt:Ankle.left:Doc:XR
C1526797|Views 2^standing:Finding:Point in time:Ankle.left:Document:XR
C1526801|Femur-L XR stand
C1526801|Femur - left X-ray standing
C1526801|Views^standing:Find:Pt:Femur.left:Doc:XR
C1526801|Views^standing:Finding:Point in time:Femur.left:Document:XR
C1526804|Hand-L XR AP+Lat+Obl
C1526804|Hand - left X-ray AP and lateral and oblique
C1526804|Views AP & lateral & oblique:Finding:Point in time:Hand.left:Document:XR
C1526804|Views AP & lateral & oblique:Find:Pt:Hand.left:Doc:XR
C1524180|Should-R CT
C1524180|Shoulder - right CT
C1524180|Multisection:Finding:Point in time:Shoulder.right:Document:Computerized Tomography
C1524180|Multisection:Find:Pt:Shoulder.right:Doc:CT
C1524812|Ankle-L MRI WO contr
C1524812|Ankle - left MRI WO contrast
C1524812|Multisection^WO contrast:Find:Pt:Ankle.left:Doc:MRI
C1524812|Multisection^WO contrast:Finding:Point in time:Ankle.left:Document:MRI
C1524822|Brst-Bl MRI WO contr
C1524822|Breast - bilateral MRI WO contrast
C1524822|Multisection^WO contrast:Find:Pt:Breast.bilateral:Doc:MRI
C1524822|Multisection^WO contrast:Finding:Point in time:Breast.bilateral:Document:MRI
C1524829|Elbow-Bl CT WO contr
C1524829|Elbow - bilateral CT WO contrast
C1524829|Multisection^WO contrast:Finding:Point in time:Elbow.bilateral:Document:Computerized Tomography
C1524829|Multisection^WO contrast:Find:Pt:Elbow.bilateral:Doc:CT
C1524853|Foot - left CT WO contrast
C1524853|Ft-L CT WO contr
C1524853|Multisection^WO contrast:Find:Pt:Foot.left:Doc:CT
C1524853|Multisection^WO contrast:Finding:Point in time:Foot.left:Document:Computerized Tomography
C1525112|Upper extremity veins - left MRI angiogram
C1525112|UE vv-L MRI.Angio
C1525112|Multisection:Finding:Point in time:Upper extremity veins.left:Document:MRI.angio
C1525112|Multisection:Find:Pt:Upper extremity veins.left:Doc:MRI.angio
C1524462|Multisection^W contrast IS:Find:Pt:Elbow.left:Doc:MRI
C1524462|Multisection^W contrast Intrasynovial:Finding:Point in time:Elbow.left:Document:MRI
C1524462|Elbow - left MRI W contrast IS
C1524462|Elbow-L MRI W contr IS
C1525191|Temporal bone CT W contrast IV
C1525191|Temporal bone CT W contr IV
C1525191|Multisection^W contrast Intravenous:Finding:Point in time:Temporal bone:Document:Computerized Tomography
C1525191|Multisection^W contrast IV:Find:Pt:Temporal bone:Doc:CT
C1525210|Multisection^WO & W contrast IV:Find:Pt:Petrous part of temporal bone:Doc:CT
C1525210|Multisection^WO & W contrast Intravenous:Finding:Point in time:Petrous part of temporal bone:Document:Computerized Tomography
C1525210|Petr part temp bone CT WO+W contr IV
C1525210|Petrous part of temporal bone CT WO and W contrast IV
C1525280|Ft-L XR 3V stand
C1525280|Foot - left X-ray 3 views standing
C1525280|Views 3^standing:Find:Pt:Foot.left:Doc:XR
C1525280|Views 3^standing:Finding:Point in time:Foot.left:Document:XR
C1525346|Should-Bl XR Stryker Notch
C1525346|Shoulder - bilateral X-ray Stryker Notch
C1525346|View Stryker Notch:Find:Pt:Shoulder.bilateral:Doc:XR
C1525346|View Stryker Notch:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525469|Knee-L XR V1 Tunnel stand
C1525469|Knee - left X-ray tunnel standing
C1525469|View tunnel^standing:Finding:Point in time:Knee.left:Document:XR
C1525469|View tunnel^standing:Find:Pt:Knee.left:Doc:XR
C1525512|Knee XR AP+Lat+Tunnel
C1525512|Knee X-ray AP and lateral and tunnel
C1525512|Views AP & lateral & tunnel:Finding:Point in time:Knee:Document:XR
C1525512|Views AP & lateral & tunnel:Find:Pt:Knee:Doc:XR
C1525645|Circle of Willis MRI.Angio W contr IV
C1525645|Circle of Willis MRI angiogram W contrast IV
C1525645|Multisection^W contrast Intravenous:Finding:Point in time:Head+Neck>Circle of Willis:Document:MRI.angio
C1525645|Multisection^W contrast IV:Find:Pt:Head+Neck>Circle of Willis:Doc:MRI.angio
C1525665|TMJ CT WO contr
C1525665|Temporomandibular joint CT WO contrast
C1525665|Multisection^WO contrast:Find:Pt:Temporomandibular joint:Doc:CT
C1525665|Multisection^WO contrast:Finding:Point in time:Temporomandibular joint:Document:Computerized Tomography
C1525666|Temporomandibular joint MRI WO contrast
C1525666|TMJ MRI WO contr
C1525666|Multisection^WO contrast:Finding:Point in time:Temporomandibular joint:Document:MRI
C1525666|Multisection^WO contrast:Find:Pt:Temporomandibular joint:Doc:MRI
C1525688|Skull+Face+Mandible XR
C1525688|Skull and Facial bones and Mandible X-ray
C1525688|Views:Finding:Point in time:Skull+Facial bones+Mandible:Document:XR
C1525688|Views:Find:Pt:Skull+Facial bones+Mandible:Doc:XR
C1525718|Carot a+VA-Bl XRA W contr IA
C1525718|Carotid artery and Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA
C1525718|Views^W contrast IA:Find:Pt:Carotid artery+Vertebral artery.bilateral:Doc:XR.fluor.angio
C1525718|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Vertebral artery.bilateral:Document:XR.fluor.angio
C1525734|Temporomandibular joint - left Fluoroscopy W contrast IS
C1525734|Views^W contrast Intrasynovial:Finding:Point in time:Temporomandibular joint.left:Document:XR.fluor
C1525734|TMJ-L Flr W contr IS
C1525734|Views^W contrast IS:Find:Pt:Temporomandibular joint.left:Doc:XR.fluor
C1525764|Wrist CT WO+W contr IV
C1525764|Multisection^WO & W contrast IV:Find:Pt:Wrist:Doc:CT
C1525764|Wrist CT WO and W contrast IV
C1525764|Multisection^WO & W contrast Intravenous:Finding:Point in time:Wrist:Document:Computerized Tomography
C1525769|Wrist - bilateral MRI WO contrast
C1525769|Wrist-Bl MRI WO contr
C1525769|Multisection^WO contrast:Find:Pt:Wrist.bilateral:Doc:MRI
C1525769|Multisection^WO contrast:Finding:Point in time:Wrist.bilateral:Document:MRI
C1525781|Ankle-L XR Lat W Stress
C1525781|Ankle - left X-ray lateral W manual stress
C1525781|Views lateral^W manual stress:Finding:Point in time:Ankle.left:Document:XR
C1525781|Views lateral^W manual stress:Find:Pt:Ankle.left:Doc:XR
C1525853|Ankle-Bl XR W Stress
C1525853|Ankle - bilateral X-ray W manual stress
C1525853|Views^W manual stress:Find:Pt:Ankle.bilateral:Doc:XR
C1525853|Views^W manual stress:Finding:Point in time:Ankle.bilateral:Document:XR
C1525877|Acromioclavicular joint - left X-ray WO and W weight
C1525877|AC joint-L XR WO+W Wt
C1525877|Views^WO & W weight:Find:Pt:Acromioclavicular joint.left:Doc:XR
C1525877|Views^WO & W weight:Finding:Point in time:Acromioclavicular joint.left:Document:XR
C1525881|Jejunum Flr W contr
C1525881|Jejunum Fluoroscopy W contrast
C1525881|Views^W contrast:Find:Pt:Jejunum:Doc:XR.fluor
C1525881|Views^W contrast:Finding:Point in time:Jejunum:Document:XR.fluor
C1525884|Ac arch+Carot a.com-Bl XRA W contr IA
C1525884|Aortic arch and Carotid artery.common - bilateral Fluoroscopic angiogram W contrast IA
C1525884|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery.common.bilateral:Document:XR.fluor.angio
C1525884|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery.common.bilateral:Doc:XR.fluor.angio
C0881988|Views^W contrast Intravenous:Finding:Point in time:Kidney+Collecting system:Narrative:XR
C0881988|Kidney XR W contr IV
C0881988|Kidney X-ray W contrast IV
C0881988|Views^W contrast IV:Find:Pt:Kidney:Doc:XR
C0881988|Views^W contrast Intravenous:Finding:Point in time:Kidney:Document:XR
C1525896|Patella X-ray Single view
C1525896|Patella XR 1V
C1525896|View 1:Find:Pt:Patella:Doc:XR
C1525896|View 1:Finding:Point in time:Patella:Document:XR
C1525937|Pelvis XR AP+Judet
C1525937|Pelvis X-ray AP and Judet
C1525937|Views AP & Judet:Finding:Point in time:Pelvis:Document:XR
C1525937|Views AP & Judet:Find:Pt:Pelvis:Doc:XR
C1525840|Wrist - bilateral X-ray oblique
C1525840|Wrist-Bl XR Obl
C1525840|Views oblique:Find:Pt:Wrist.bilateral:Doc:XR
C1525840|Views oblique:Finding:Point in time:Wrist.bilateral:Document:XR
C1525956|Views:Finding:Point in time:Neck:Narrative:XR
C1525956|Neck X-ray
C1525956|Neck XR
C1525956|Views:Finding:Point in time:Neck:Document:XR
C1525956|Views:Find:Pt:Neck:Doc:XR
C1525983|Ankle-R XR AP+Lat
C1525983|Ankle - right X-ray AP and lateral
C1525983|Views AP & lateral:Find:Pt:Ankle.right:Doc:XR
C1525983|Views AP & lateral:Finding:Point in time:Ankle.right:Document:XR
C1526002|Elbow-R XR 2V Obl
C1526002|Elbow - right X-ray 2 views Oblique
C1526002|Views 2 oblique:Finding:Point in time:Elbow.right:Document:XR
C1526002|Views 2 oblique:Find:Pt:Elbow.right:Doc:XR
C1526050|Lower extremity - right X-ray standing
C1526050|LE-R XR stand
C1526050|View^standing:Finding:Point in time:Lower extremity.right:Document:XR
C1526050|View^standing:Find:Pt:Lower extremity.right:Doc:XR
C1526052|Humerus-R XR AP+Lat
C1526052|Humerus - right X-ray AP and lateral
C1526052|Views AP & lateral:Finding:Point in time:Humerus.right:Document:XR
C1526052|Views AP & lateral:Find:Pt:Humerus.right:Doc:XR
C1526053|Humerus - right X-ray oblique
C1526053|Humerus-R XR Obl
C1526053|Views oblique:Finding:Point in time:Humerus.right:Document:XR
C1526053|Views oblique:Find:Pt:Humerus.right:Doc:XR
C1526078|Knee-R XR 2V stand
C1526078|Knee - right X-ray 2 views standing
C1526078|Views 2^standing:Find:Pt:Knee.right:Doc:XR
C1526078|Views 2^standing:Finding:Point in time:Knee.right:Document:XR
C1525124|Brst-R Mam
C1525124|Breast - right Mammogram
C1525124|Views:Finding:Point in time:Breast.right:Document:Mam
C1525124|Views:Find:Pt:Breast.right:Doc:Mam
C1526137|Shoulder X-ray outlet
C1526137|Should XR Outlet
C1526137|View outlet:Find:Pt:Shoulder:Doc:XR
C1526137|View outlet:Finding:Point in time:Shoulder:Document:XR
C1526164|Skull X-ray lateral crosstable
C1526164|Skull XR Lat Xtable
C1526164|View lateral crosstable:Find:Pt:Skull:Doc:XR
C1526164|View lateral crosstable:Finding:Point in time:Skull:Document:XR
C1526179|Tib+Fib XR stand
C1526179|Tibia and Fibula X-ray standing
C1526179|Views^standing:Find:Pt:Tibia+Fibula:Doc:XR
C1526179|Views^standing:Finding:Point in time:Tibia+Fibula:Document:XR
C1524710|Wrist X-ray tomograph
C1524710|Wrist XRTomo
C1524710|Multisection:Find:Pt:Wrist:Doc:XR.tomo
C1524710|Multisection:Finding:Point in time:Wrist:Document:XR.tomo
C1526208|Ribs posterior X-ray
C1526208|Ribs post XR
C1526208|Views:Find:Pt:Ribs.posterior:Doc:XR
C1526208|Views:Finding:Point in time:Ribs.posterior:Document:XR
C1526232|UE aa-R XRA W contr IA
C1526232|Upper extremity arteries - right Fluoroscopic angiogram W contrast IA
C1526232|Upper extremity arteries - right Narrative Fluoroscopic angiogram W contrast IA
C1526232|Views^W contrast IA:Find:Pt:Upper extremity arteries.right:Doc:XR.fluor.angio
C1526232|Views^W contrast Intra-arterial:Finding:Point in time:Upper extremity arteries.right:Document:XR.fluor.angio
C1526238|Testicle ves Flr W contr
C1526238|Testicle vessels Fluoroscopy W contrast
C1526238|Views^W contrast:Find:Pt:Testicle vessels:Doc:XR.fluor
C1526238|Views^W contrast:Finding:Point in time:Testicle vessels:Document:XR.fluor
C1525145|Guidance for drainage:Find:Pt:Chest:Doc:US
C1525145|Guidance for drainage:Finding:Point in time:Chest:Document:Ultrasound
C1525145|Chest US Drain guid
C1525145|US Guidance for drainage of Chest
C1526344|Toe fifth - right X-ray
C1526344|Toe 5th-R XR
C1526344|Views:Find:Pt:Toe.fifth.right:Doc:XR
C1526344|Views:Finding:Point in time:Toe.fifth.right:Document:XR
C1524508|LE-L CT W contr IV
C1524508|Lower extremity - left CT W contrast IV
C1524508|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.left:Document:Computerized Tomography
C1524508|Multisection^W contrast IV:Find:Pt:Lower extremity.left:Doc:CT
C1524865|Hand - right CT WO contrast
C1524865|Hand-R CT WO contr
C1524865|Multisection^WO contrast:Finding:Point in time:Hand.right:Document:Computerized Tomography
C1524865|Multisection^WO contrast:Find:Pt:Hand.right:Doc:CT
C1524900|Pancreas MRI WO contrast
C1524900|Pancreas MRI WO contr
C1524900|Multisection^WO contrast:Finding:Point in time:Pancreas:Document:MRI
C1524900|Multisection^WO contrast:Find:Pt:Pancreas:Doc:MRI
C1524912|Thyroid MRI WO contr
C1524912|Thyroid MRI WO contrast
C1524912|Multisection^WO contrast:Finding:Point in time:Thyroid:Document:MRI
C1524912|Multisection^WO contrast:Find:Pt:Thyroid:Doc:MRI
C1524914|Lower leg-L CT WO contr
C1524914|Lower leg - left CT WO contrast
C1524914|Multisection^WO contrast:Finding:Point in time:Lower leg.left:Document:Computerized Tomography
C1524914|Multisection^WO contrast:Find:Pt:Lower leg.left:Doc:CT
C1524307|Thyroid CT Bx guid
C1524307|CT Guidance for biopsy of Thyroid
C1524307|Guidance for biopsy:Finding:Point in time:Thyroid:Document:Computerized Tomography
C1524307|Guidance for biopsy:Find:Pt:Thyroid:Doc:CT
C1524591|Sternum CT W contr IV
C1524591|Sternum CT W contrast IV
C1524591|Multisection^W contrast IV:Find:Pt:Sternum:Doc:CT
C1524591|Multisection^W contrast Intravenous:Finding:Point in time:Sternum:Document:Computerized Tomography
C1524616|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.left:Doc:CT
C1524616|LE-L CT WO+W contr IV
C1524616|Lower extremity - left CT WO and W contrast IV
C1524616|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.left:Document:Computerized Tomography
C1524976|Internal auditory canal X-ray
C1524976|IAC XR
C1524976|Views:Finding:Point in time:Internal auditory canal:Document:XR
C1524976|Views:Find:Pt:Internal auditory canal:Doc:XR
C1524339|Ankle - bilateral CT
C1524339|Ankle-Bl CT
C1524339|Multisection:Find:Pt:Ankle.bilateral:Doc:CT
C1524339|Multisection:Finding:Point in time:Ankle.bilateral:Document:Computerized Tomography
C1524638|Mandible XR 3V
C1524638|Mandible X-ray 3 views
C1524638|Views 3:Find:Pt:Mandible:Doc:XR
C1524638|Views 3:Finding:Point in time:Mandible:Document:XR
C1524652|Knee - left X-ray 4 views
C1524652|Knee-L XR 4V
C1524652|Views 4:Find:Pt:Knee.left:Doc:XR
C1524652|Views 4:Finding:Point in time:Knee.left:Document:XR
C1524353|IAC CT
C1524353|Internal auditory canal CT
C1524353|Multisection:Find:Pt:Internal auditory canal:Doc:CT
C1524353|Multisection:Finding:Point in time:Internal auditory canal:Document:Computerized Tomography
C1524361|Elbow - left X-ray tomograph
C1524361|Elbow-L XRTomo
C1524361|Multisection:Finding:Point in time:Elbow.left:Document:XR.tomo
C1524361|Multisection:Find:Pt:Elbow.left:Doc:XR.tomo
C1527031|Foot CT
C1527031|Ft CT
C1527031|Multisection:Find:Pt:Foot:Doc:CT
C1527031|Multisection:Finding:Point in time:Foot:Document:Computerized Tomography
C1524747|Hip-Bl MRI WO+W contr IV
C1524747|Multisection^WO & W contrast IV:Find:Pt:Hip.bilateral:Doc:MRI
C1524747|Hip - bilateral MRI WO and W contrast IV
C1524747|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip.bilateral:Document:MRI
C1525052|Patella-L XR AP+Lat
C1525052|Patella - left X-ray AP and lateral
C1525052|Views AP & lateral:Finding:Point in time:Patella.left:Document:XR
C1525052|Views AP & lateral:Find:Pt:Patella.left:Doc:XR
C1524790|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sternum:Document:Computerized Tomography
C1524790|Sternum CT WO+W contr IV
C1524790|Multisection^WO & W contrast IV:Find:Pt:Sternum:Doc:CT
C1524790|Sternum CT WO and W contrast IV
C1524806|Upper extremity Vessels CT angiogram WO and W contrast IV
C1524806|Multisection^WO & W contrast IV:Find:Pt:Upper extremity>Vessels:Doc:CT.angio
C1524806|EU ves CT.Angio WO+W contr IV
C1524806|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity>Vessels:Document:Computerized Tomography.angio
C1524678|Elbow - bilateral X-ray oblique
C1524678|Elbow-Bl XR Obl
C1524678|Views oblique:Find:Pt:Elbow.bilateral:Doc:XR
C1524678|Views oblique:Finding:Point in time:Elbow.bilateral:Document:XR
C1525072|Humerus - left X-ray oblique
C1525072|Humerus-L XR Obl
C1525072|Views oblique:Finding:Point in time:Humerus.left:Document:XR
C1525072|Views oblique:Find:Pt:Humerus.left:Doc:XR
C1525074|Knee-L XR Obl
C1525074|Knee - left X-ray oblique
C1525074|Views oblique:Find:Pt:Knee.left:Doc:XR
C1525074|Views oblique:Finding:Point in time:Knee.left:Document:XR
C1830217|Multisection^WO & W reduced contrast volume Intravenous:Finding:Point in time:Head:Document:Computerized Tomography
C1830217|Head CT WO+W red contr vol IV
C1830217|Multisection^WO & W reduced contrast volume IV:Find:Pt:Head:Doc:CT
C1830217|Head CT WO and W reduced contrast volume IV
C1830223|Kidney CT W contr IV
C1830223|Kidney CT W contrast IV
C1830223|Multisection^W contrast IV:Find:Pt:Kidney:Doc:CT
C1830223|Multisection^W contrast Intravenous:Finding:Point in time:Kidney:Document:Computerized Tomography
C1830240|Brst-UL Mam
C1830240|Breast - unilateral Mammogram
C1830240|Views:Find:Pt:Breast.unilateral:Doc:Mam
C1830240|Views:Finding:Point in time:Breast.unilateral:Document:Mam
C1830069|Chest CT Ltd WO contr
C1830069|Chest CT limited WO contrast
C1830069|Multisection limited^WO contrast:Finding:Point in time:Chest:Document:Computerized Tomography
C1830069|Multisection limited^WO contrast:Find:Pt:Chest:Doc:CT
C1715380|CT Guidance for fine needle aspiration of Adrenal gland
C1715380|Adrenal CT FNA Asp
C1715380|Guidance for aspiration.fine needle:Find:Pt:Abdomen>Adrenal gland:Doc:CT
C1715380|Guidance for aspiration.fine needle:Finding:Point in time:Abdomen>Adrenal gland:Document:Computerized Tomography
C1717311|Guidance for biopsy:Find:Pt:Abdomen>Retroperitoneum:Doc:CT
C1717311|Retroperitoneum CT Bx guid
C1717311|Guidance for biopsy:Finding:Point in time:Abdomen>Retroperitoneum:Document:Computerized Tomography
C1717311|CT Guidance for biopsy of Retroperitoneum
C1715396|Hrt MRI Cine for Flow VM W contr IV
C1715396|Heart MRI cine for blood flow velocity mapping W contrast IV
C1715396|Multisection cine for blood flow velocity mapping^W contrast Intravenous:Finding:Point in time:Heart:Document:MRI
C1715396|Multisection cine for blood flow velocity mapping^W contrast IV:Find:Pt:Heart:Doc:MRI
C1715404|Multisection^WO & W contrast Intravenous:Finding:Point in time:Renal vessels:Document:MRI.angio
C1715404|Multisection^WO & W contrast IV:Find:Pt:Renal vessels:Doc:MRI.angio
C1715404|Renal vessels MRI angiogram WO and W contrast IV
C1715404|Renal ves MRI.Angio WO+W contr IV
C1715405|Lower extremity vessels - bilateral MRI angiogram W contrast IV
C1715405|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity vessels.bilateral:Document:MRI.angio
C1715405|Multisection^W contrast IV:Find:Pt:Lower extremity vessels.bilateral:Doc:MRI.angio
C1715405|LE ves-Bl MRI.Angio W contr IV
C1715415|Thyroid RI +Uptake W Tc99mP IV
C1715415|Thyroid Scan and uptake W Tc-99m pertechnetate IV
C1715415|Views & uptake^W Tc-99m pertechnetate Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1715415|Views & uptake^W Tc-99m pertechnetate IV:Find:Pt:Thyroid:Doc:Radnuc
C1715458|Knee X-ray GE 5 views
C1715458|Knee XR GE 5V
C1715458|Views GE 5:Find:Pt:Knee:Doc:XR
C1715458|Views GE 5:Finding:Point in time:Knee:Document:XR
C1715491|Views^WO & W Tc-99m Mertiatide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1715491|Kdny-Bl RI WO+W Tc99mMertiatide IV
C1715491|Kidney - bilateral Scan WO and W Tc-99m Mertiatide IV
C1715491|Views^WO & W Tc-99m Mertiatide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1643599|UE a-L US
C1643599|Upper extremity artery - left US
C1643599|Multisection:Finding:Point in time:Upper extremity artery.left:Document:Ultrasound
C1643599|Multisection:Find:Pt:Upper extremity artery.left:Doc:US
C1632790|C-spine Flr Ltd W contr IT
C1632790|Views limited^W contrast IT:Find:Pt:Spine.cervical:Doc:XR.fluor
C1632790|Views limited^W contrast Intrathecal:Finding:Point in time:Spine.cervical:Document:XR.fluor
C1632790|Cervical spine Fluoroscopy limited W contrast IT
C1628565|Brain+Pituitary+ST MRI WO contr
C1628565|Brain and Pituitary and Sella turcica MRI WO contrast
C1628565|Multisection^WO contrast:Finding:Point in time:Brain+Pituitary+Sella turcica:Document:MRI
C1628565|Multisection^WO contrast:Find:Pt:Brain+Pituitary+Sella turcica:Doc:MRI
C1714806|XXX XR of FB
C1714806|Unspecified body region X-ray of foreign body
C1714806|Views of foreign body:Find:Pt:XXX:Doc:XR
C1714806|Views of foreign body:Finding:Point in time:To be specified in another part of the message:Document:XR
C1714807|Skull X-ray LE 3 views
C1714807|Skull XR LE 3V
C1714807|Views LE 3:Find:Pt:Skull:Doc:XR
C1714807|Views LE 3:Finding:Point in time:Skull:Document:XR
C1714911|Axilla-R MRI
C1714911|Axilla - right MRI
C1714911|Multisection:Find:Pt:Axilla.right:Doc:MRI
C1714911|Multisection:Finding:Point in time:Axilla.right:Document:MRI
C1714916|Wrist vessels - left MRI angiogram WO contrast
C1714916|Wrist Ves-L MRI.Angio WO contr
C1714916|Multisection^WO contrast:Find:Pt:Wrist vessels.left:Doc:MRI.angio
C1714916|Multisection^WO contrast:Finding:Point in time:Wrist vessels.left:Document:MRI.angio
C1714920|Mandible X-ray 1 or 2 views
C1714920|Mandible XR 1V or 2V
C1714920|Views 1 or 2:Find:Pt:Mandible:Doc:XR
C1714920|Views 1 or 2:Finding:Point in time:Mandible:Document:XR
C1715092|Vein-R XRA Thrombect guid W contr IV
C1715092|Fluoroscopic angiogram Guidance for thrombectomy of Vein - right-- W contrast IV
C1715092|Guidance for thrombectomy^W contrast Intravenous:Finding:Point in time:Vein.right:Document:XR.fluor.angio
C1715092|Guidance for thrombectomy^W contrast IV:Find:Pt:Vein.right:Doc:XR.fluor.angio
C1715120|Tibioperoneal arteries - bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C1715120|Angioplasty^W contrast IA:Find:Pt:Tibioperoneal arteries.bilateral:Doc:XR.fluor.angio
C1715120|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibioperoneal arteries.bilateral:Document:XR.fluor.angio
C1715120|Tibioperon aa-Bl XRA Angpsty W contr IA
C1635011|Sella turcica X-ray 2 views
C1635011|ST XR 2V
C1635011|Views 2:Find:Pt:Sella turcica:Doc:XR
C1635011|Views 2:Finding:Point in time:Sella turcica:Document:XR
C1639941|Abd Flr Replac of PCS guid
C1639941|Fluoroscopy Guidance for replacement of percutaneous cholecystostomy in Abdomen
C1639941|Guidance for replacement of percutaneous cholecystostomy:Find:Pt:Abdomen:Doc:XR.fluor
C1639941|Guidance for replacement of percutaneous cholecystostomy:Finding:Point in time:Abdomen:Document:XR.fluor
C1637286|Brst-R US Cyst Asp guid
C1637286|US Guidance for aspiration of cyst of Breast - right
C1637286|Guidance for aspiration of cyst:Find:Pt:Breast.right:Doc:US
C1637286|Guidance for aspiration of cyst:Finding:Point in time:Breast.right:Document:Ultrasound
C1626768|Shunt X-ray
C1626768|Shunt XR
C1626768|Views:Finding:Point in time:Shunt.To be specified in another part of the message:Document:XR
C1626768|Views:Find:Pt:Shunt.XXX:Doc:XR
C1632269|Ribs+Chest XR +PA Chst
C1632269|Ribs and Chest X-ray and PA chest
C1632269|Views & PA chest:Find:Pt:Ribs+Chest:Doc:XR
C1632269|Views & PA chest:Finding:Point in time:Ribs+Chest:Document:XR
C1642088|Elbow - right X-ray portable
C1642088|Elbow-R XR port
C1642088|Views portable:Finding:Point in time:Elbow.right:Document:XR
C1642088|Views portable:Find:Pt:Elbow.right:Doc:XR
C1635651|Colon Flr Ltd W Air+Ba PR
C1635651|Colon Fluoroscopy limited W air and barium contrast PR
C1635651|Views limited^W air & barium contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C1635651|Views limited^W air & barium contrast PR:Find:Pt:Colon:Doc:XR.fluor
C1630750|CT Guidance for biopsy of Kidney
C1630750|Kidney CT Bx guid
C1630750|Guidance for biopsy:Finding:Point in time:Kidney:Document:Computerized Tomography
C1630750|Guidance for biopsy:Find:Pt:Kidney:Doc:CT
C1630178|Guidance for drainage of abscess:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1630178|Guidance for drainage of abscess:Find:Pt:Pelvis:Doc:CT
C1630178|CT Guidance for drainage of abscess of Pelvis
C1630178|Pelvis CT Abscess drain guid
C1632955|Head vessels CT angiogram WO contrast
C1632955|Multisection^WO contrast:Finding:Point in time:Head>Vessels:Document:Computerized Tomography.angio
C1632955|Multisection^WO contrast:Find:Pt:Head>Vessels:Doc:CT.angio
C1632955|Head vess CT.Angio WO contr
C1632339|Orbit-L XR for FB
C1632339|Orbit - left X-ray for foreign body
C1632339|Views for foreign body:Finding:Point in time:Orbit.left:Document:XR
C1632339|Views for foreign body:Find:Pt:Orbit.left:Doc:XR
C1954363|Mammogram Guidance for localization of Breast
C1954363|Brst Mam Localization guid
C1954363|Guidance for localization:Find:Pt:Breast:Doc:Mam
C1954363|Guidance for localization:Finding:Point in time:Breast:Document:Mam
C1953327|Lower extremity arteries - left Fluoroscopic angiogram W contrast IA
C1953327|LE aa-L XRA W contr IA
C1953327|Views^W contrast Intra-arterial:Finding:Point in time:Lower extremity arteries.left:Document:XR.fluor.angio
C1953327|Views^W contrast IA:Find:Pt:Lower extremity arteries.left:Doc:XR.fluor.angio
C1953951|Larynx MRI WO contr
C1953951|Larynx MRI WO contrast
C1953951|Multisection^WO contrast:Find:Pt:Larynx:Doc:MRI
C1953951|Multisection^WO contrast:Finding:Point in time:Larynx:Document:MRI
C1953963|Clavicle-L MRI W contr IV
C1953963|Clavicle - left MRI W contrast IV
C1953963|Multisection^W contrast IV:Find:Pt:Clavicle.left:Doc:MRI
C1953963|Multisection^W contrast Intravenous:Finding:Point in time:Clavicle.left:Document:MRI
C3174151|Mammary artery.internal - left Fluoroscopic angiogram W contrast IA
C3174151|IMAl-L XRA W contr IA
C3174151|Views^W contrast Intra-arterial:Finding:Point in time:Mammary artery.internal.left:Document:XR.fluor.angio
C3174151|Views^W contrast IA:Find:Pt:Mammary artery.internal.left:Doc:XR.fluor.angio
C3174364|Fluoroscopic angiogram Guidance for placement of stent in Artery - left
C3174364|Artery-L XRA Stent plac guid
C3174364|Guidance for placement of stent:Finding:Point in time:Artery.left:Document:XR.fluor.angio
C3174364|Guidance for placement of stent:Find:Pt:Artery.left:Doc:XR.fluor.angio
C3533552|Guidance for repair of CVA catheter with port or pump:Find:Pt:Central vein:Doc:XR.fluor
C3533552|Centl v Flr CVA cath W pump repair guid
C3533552|Guidance for repair of CVA catheter with port or pump:Finding:Point in time:Central vein:Document:XR.fluor
C3533552|Fluoroscopy Guidance for repair of CVA catheter with port or pump of Central vein
C3533806|Toes-R MRI WO contr
C3533806|Multisection^WO contrast:Finding:Point in time:Toes.right:Document:MRI
C3533806|Multisection^WO contrast:Find:Pt:Toes.right:Doc:MRI
C3533806|Toes - right MRI WO contrast
C3262989|MRI Guidance for biopsy of Breast - bilateral
C3262989|Brst-Bl MRI Bx guid
C3262989|Guidance for biopsy:Find:Pt:Breast.bilateral:Doc:MRI
C3262989|Guidance for biopsy:Finding:Point in time:Breast.bilateral:Document:MRI
C3482441|C-spine US
C3482441|Multisection:Finding:Point in time:Spine.cervical:Document:Ultrasound
C3482441|Multisection:Find:Pt:Spine.cervical:Doc:US
C3482441|Cervical spine US
C3263015|Finger MRI W contrast IV
C3263015|Finger MRI W contr IV
C3263015|Multisection^W contrast IV:Find:Pt:Finger:Doc:MRI
C3263015|Multisection^W contrast Intravenous:Finding:Point in time:Finger:Document:MRI
C3263056|Lung Flr PC Abscess Drain guid
C3263056|Fluoroscopy Guidance for percutaneous drainage of abscess of Lung
C3263056|Guidance for percutaneous drainage of abscess:Finding:Point in time:Lung:Document:XR.fluor
C3263056|Guidance for percutaneous drainage of abscess:Find:Pt:Lung:Doc:XR.fluor
C3263080|Breast duct Mammogram Single view W contrast intra duct
C3263080|Brst.duct Mam 1V W contr intra Dct
C3263080|View 1^W contrast intra duct:Find:Pt:Breast.duct:Doc:Mam
C3263080|View 1^W contrast intra duct:Finding:Point in time:Breast.duct:Document:Mam
C3261471|Humerus - left X-ray Single view
C3261471|Humerus-L XR 1V
C3261471|View 1:Finding:Point in time:Humerus.left:Document:XR
C3261471|View 1:Find:Pt:Humerus.left:Doc:XR
C3262881|Hand - bilateral X-ray AP and lateral and oblique
C3262881|Hand-Bl XR AP+Lat+Obl
C3262881|Views AP & lateral & oblique:Finding:Point in time:Hand.bilateral:Document:XR
C3262881|Views AP & lateral & oblique:Find:Pt:Hand.bilateral:Doc:XR
C3262918|Bladder CT W contr IV
C3262918|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis>Urinary bladder:Document:Computerized Tomography
C3262918|Multisection^W contrast IV:Find:Pt:Abdomen+Pelvis>Urinary bladder:Doc:CT
C3262918|Urinary bladder CT W contrast IV
C2709260|Deprecated Multisection:Finding:Point in time:Thigh.bilateral:Narrative:MRI
C2709260|Multisection:Find:Pt:Thigh.bilateral:Nar:MRI
C2709260|Deprecated Thigh Bilateral MRI Multisection
C2709260|Deprecated Thigh-Bl MRI
C2709260|Multisection:Finding:Point in time:Thigh.bilateral:Narrative:MRI
C0942303|Brst-L Mam Needle local mass guid
C0942303|Mammogram Guidance for needle localization of mass of Breast - left
C0942303|Guidance for needle localization of mass:Find:Pt:Breast.left:Doc:Mam
C0942303|Guidance for needle localization of mass:Finding:Point in time:Breast.left:Document:Mam
C0942362|Shoulder - left X-ray 3 views
C0942362|Should-L XR 3V
C0942362|Views 3:Finding:Point in time:Shoulder.left:Document:XR
C0942362|Views 3:Find:Pt:Shoulder.left:Doc:XR
C0942377|Hip - right X-ray Single view
C0942377|Hip-R XR 1V
C0942377|View 1:Find:Pt:Hip.right:Doc:XR
C0942377|View 1:Finding:Point in time:Hip.right:Document:XR
C0882020|Lung Scan portable
C0882020|Lung RI port W RNC IV
C0882020|Views portable^W radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C0882020|Views portable^W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C0882213|Multisection:Finding:Point in time:To be specified in another part of the message:Narrative:ULTRASOUND
C0882213|Unspecified body region US
C0882213|XXX US
C0882213|Multisection:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C0882213|Multisection:Find:Pt:XXX:Doc:US
C0882227|Renal v-Bl XRA W contr IV+Renin Samp
C0882227|Renal vein - bilateral Fluoroscopic angiogram W contrast IV and W renin sampling
C0882227|Views^W contrast IV & W renin sampling:Find:Pt:Renal vein.bilateral:Doc:XR.fluor.angio
C0882227|Views^W contrast Intravenous & W renin sampling:Finding:Point in time:Renal vein.bilateral:Document:XR.fluor.angio
C0945308|Clavicle-L XR
C0945308|Clavicle - left X-ray
C0945308|Views:Finding:Point in time:Clavicle.left:Document:XR
C0945308|Views:Find:Pt:Clavicle.left:Doc:XR
C0881848|Carotid artery intracranial Fluoroscopic angiogram Angioplasty W contrast IA
C0881848|Carot a.IC XRA Angpsty W contr IA
C0881848|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Carotid artery.intracranial:Document:XR.fluor.angio
C0881848|Angioplasty^W contrast IA:Find:Pt:Carotid artery.intracranial:Doc:XR.fluor.angio
C0882524|Chest X-ray lordotic
C0882524|Chest XR Lordonic
C0882524|View lordotic:Finding:Point in time:Chest:Document:XR
C0882524|View lordotic:Find:Pt:Chest:Doc:XR
C0881950|Head US in Surg
C0881950|Head US during surgery
C0881950|Multisection^during surgery:Finding:Point in time:Head:Document:Ultrasound
C0881950|Multisection^during surgery:Find:Pt:Head:Doc:US
C0881966|Hip XR 1V
C0881966|Hip X-ray Single view
C0881966|View 1:Find:Pt:Hip:Doc:XR
C0881966|View 1:Finding:Point in time:Hip:Document:XR
C1114478|Brain MRI Local Str Guid W contr IV
C1114478|MRI Guidance.stereotactic for localization in Brain-- W contrast IV
C1114478|Guidance.stereotactic for localization^W contrast IV:Find:Pt:Brain:Doc:MRI
C1114478|Guidance.stereotactic for localization^W contrast Intravenous:Finding:Point in time:Brain:Document:MRI
C1114495|Pelvis MRI WO contrast
C1114495|Pelvis MRI WO contr
C1114495|Multisection^WO contrast:Find:Pt:Pelvis:Doc:MRI
C1114495|Multisection^WO contrast:Finding:Point in time:Pelvis:Document:MRI
C1114503|Forearm MRI WO contr
C1114503|Forearm MRI WO contrast
C1114503|Multisection^WO contrast:Finding:Point in time:Forearm:Document:MRI
C1114503|Multisection^WO contrast:Find:Pt:Forearm:Doc:MRI
C1114524|Upper extremity US
C1114524|UE US
C1114524|Multisection:Find:Pt:Upper extremity:Doc:US
C1114524|Multisection:Finding:Point in time:Upper extremity:Document:Ultrasound
C1114553|Chest XR R-or-L-Obl
C1114553|Chest X-ray right or-left oblique
C1114553|Views R-or-L-oblique:Finding:Point in time:Chest:Document:XR
C1114553|Views R-or-L-oblique:Find:Pt:Chest:Doc:XR
C1114598|Wrist XR AP+Lat
C1114598|Wrist X-ray AP and lateral
C1114598|Views AP & lateral:Find:Pt:Wrist:Doc:XR
C1114598|Views AP & lateral:Finding:Point in time:Wrist:Document:XR
C1114637|Aorta+Fem a-Bl XRA Runoff W contr IA
C1114637|Aorta and Femoral artery - bilateral Fluoroscopic angiogram runoff W contrast IA
C1114637|Views runoff^W contrast IA:Find:Pt:Aorta+Femoral artery.bilateral:Doc:XR.fluor.angio
C1114637|Views runoff^W contrast Intra-arterial:Finding:Point in time:Aorta+Femoral artery.bilateral:Document:XR.fluor.angio
C1114666|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower leg:Document:MRI
C1114666|Lower leg MRI WO+W contr IV
C1114666|Multisection^WO & W contrast IV:Find:Pt:Lower leg:Doc:MRI
C1114666|Lower leg MRI WO and W contrast IV
C1114667|Fem ves MRI.Angio
C1114667|Femoral vessels MRI angiogram
C1114667|Multisection:Find:Pt:Femoral vessels:Doc:MRI.angio
C1114667|Multisection:Finding:Point in time:Femoral vessels:Document:MRI.angio
C1114411|CT Guidance for injection of Spine facet joint
C1114411|Spine facet joint CT Inj guid
C1114411|Guidance for injection:Find:Pt:Spine facet joint:Doc:CT
C1114411|Guidance for injection:Finding:Point in time:Spine facet joint:Document:Computerized Tomography
C1114414|CT Guidance for radiation treatment of Unspecified body region-- WO contrast
C1114414|XXX CT RT guid WO contr
C1114414|Guidance for radiation treatment^WO contrast:Find:Pt:XXX:Doc:CT
C1114414|Guidance for radiation treatment^WO contrast:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1114470|Periph a XRA Angpsty W contr IA
C1114470|Peripheral artery Fluoroscopic angiogram Angioplasty W contrast IA
C1114470|Angioplasty^W contrast IA:Find:Pt:Peripheral artery:Doc:XR.fluor.angio
C1114470|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Peripheral artery:Document:XR.fluor.angio
C1114473|Brst US Bx CN guid
C1114473|US Guidance for core needle biopsy of Breast
C1114473|Guidance for biopsy.core needle:Find:Pt:Breast:Doc:US
C1114473|Guidance for biopsy.core needle:Finding:Point in time:Breast:Document:Ultrasound
C1526822|Ribs lower-L XR
C1526822|Ribs lower - left X-ray
C1526822|Views:Find:Pt:Ribs.lower.left:Doc:XR
C1526822|Views:Finding:Point in time:Ribs.lower.left:Document:XR
C1543751|Hrt RI PF Rest+W Tc99mMIBI IV
C1543751|Heart Scan perfusion at rest and W Tc-99m Sestamibi IV
C1543751|Views perfusion^at rest & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543751|Views perfusion^at rest & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543753|Hrt RI PF W ADE+RNC IV
C1543753|Heart Scan perfusion W adenosine and W radionuclide IV
C1543753|Views perfusion^W adenosine & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543753|Views perfusion^W adenosine & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543466|Knee-R XR 4V+Tunnel
C1543466|Knee - right X-ray 4 views and tunnel
C1543466|Views 4 & tunnel:Find:Pt:Knee.right:Doc:XR
C1543466|Views 4 & tunnel:Finding:Point in time:Knee.right:Document:XR
C2713300|Knee-R XR +Tunnel
C2713300|Knee - right X-ray and tunnel
C2713300|Views & tunnel:Find:Pt:Knee.right:Doc:XR
C2713300|Views & tunnel:Finding:Point in time:Knee.right:Document:XR
C1543486|T-spine XRTomo Lat
C1543486|Multisection lateral:Finding:Point in time:Spine.thoracic:Document:XR.tomo
C1543486|Multisection lateral:Find:Pt:Spine.thoracic:Doc:XR.tomo
C1543486|Thoracic spine X-ray tomograph lateral
C1543903|Bone SPECT 3 Phase WB W RNC IV
C1543903|Bone SPECT 3 phase whole body
C1543903|Multisection 3 phase whole body^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1543903|Multisection 3 phase whole body^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1543914|Hrt RI for Infarct+FP W RNC IV
C1543914|Heart Scan for infarct and first pass
C1543914|Views for infarct & first pass^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543914|Views for infarct & first pass^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543929|BM RI Mul Areas W RNC IV
C1543929|Bone marrow Scan multiple areas
C1543929|Views multiple areas^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc
C1543929|Views multiple areas^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc
C1543171|Ribs XR AP 1V
C1543171|Ribs X-ray AP single view
C1543171|View AP:Finding:Point in time:Ribs:Document:XR
C1543171|View AP:Find:Pt:Ribs:Doc:XR
C1543220|Ribs - bilateral and Chest X-ray 4 views and PA chest
C1543220|Views 4 & PA chest:Find:Pt:Ribs.bilateral+Chest:Doc:XR
C1543220|Views 4 & PA chest:Finding:Point in time:Ribs.bilateral+Chest:Document:XR
C1543220|Ribs-Bl+Chest XR 4V+PA Chst
C1543261|Hrt MRI Cine for Flow VM
C1543261|Heart MRI cine for blood flow velocity mapping
C1543261|Multisection cine for blood flow velocity mapping:Find:Pt:Heart:Doc:MRI
C1543261|Multisection cine for blood flow velocity mapping:Finding:Point in time:Heart:Document:MRI
C1524262|Should-R XR AP+West Point
C1524262|Shoulder - right X-ray AP and West Point
C1524262|Views AP & West Point:Find:Pt:Shoulder.right:Doc:XR
C1524262|Views AP & West Point:Finding:Point in time:Shoulder.right:Document:XR
C1526759|Clavicle-R XR 45 Deg Ceph Angle
C1526759|Clavicle - right X-ray 45 degree cephalic angle
C1526759|View 45 degree cephalic angle:Find:Pt:Clavicle.right:Doc:XR
C1526759|View 45 degree cephalic angle:Finding:Point in time:Clavicle.right:Document:XR
C1526775|Hip-R XR Lat in Surg
C1526775|Hip - right X-ray lateral during surgery
C1526775|View lateral^during surgery:Find:Pt:Hip.right:Doc:XR
C1526775|View lateral^during surgery:Finding:Point in time:Hip.right:Document:XR
C1543722|Hrt RI Rest+W DPY+RNC IV
C1543722|Heart Scan at rest and W dipyridamole and W radionuclide IV
C1543722|Views^at rest & W dipyridamole & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543722|Views^at rest & W dipyridamole & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543725|Hrt RI Rest+stress+W RNC IV
C1543725|Heart Scan at rest and W stress and W radionuclide IV
C1543725|Views^at rest & W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543725|Views^at rest & W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542971|RI Static for Inf W Ga-67 IV
C1542971|Views static for infection^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542971|Views static for infection^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1542971|Scan static for infection W Ga-67 IV
C1526781|Breast duct - right Mammogram W contrast intra duct
C1526781|Brst.duct-R Mam W contr intra Dct
C1526781|Views^W contrast intra duct:Find:Pt:Breast.duct.right:Doc:Mam
C1526781|Views^W contrast intra duct:Finding:Point in time:Breast.duct.right:Document:Mam
C1526818|Carot a+Cerebral a-L XRA W contr IA
C1526818|Carotid artery and Cerebral artery - left Fluoroscopic angiogram W contrast IA
C1526818|Views^W contrast IA:Find:Pt:Carotid artery+Cerebral artery.left:Doc:XR.fluor.angio
C1526818|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Cerebral artery.left:Document:XR.fluor.angio
C1543408|Spine CT W contrast intradisc
C1543408|Spine CT W contr ID
C1543408|Multisection^W contrast intradisc:Find:Pt:Spine:Doc:CT
C1543408|Multisection^W contrast intradisc:Finding:Point in time:Spine:Document:Computerized Tomography
C1543410|Wrist - left X-ray PA W clenched fist
C1543410|Wrist-L XR PA V1 W clenched fist
C1543410|View PA^W clenched fist:Finding:Point in time:Wrist.left:Document:XR
C1543410|View PA^W clenched fist:Find:Pt:Wrist.left:Doc:XR
C1525314|Hip - bilateral X-ray Judet
C1525314|Hip-Bl XR Judet
C1525314|View Judet:Finding:Point in time:Hip.bilateral:Document:XR
C1525314|View Judet:Find:Pt:Hip.bilateral:Doc:XR
C1525226|Upper extremity veins - right MRI angiogram WO and W contrast IV
C1525226|Multisection^WO & W contrast IV:Find:Pt:Upper extremity veins.right:Doc:MRI.angio
C1525226|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity veins.right:Document:MRI.angio
C1525226|UE vv-R MRI.Angio WO+W contr IV
C1525263|Head CT Bx Str Guid
C1525263|CT Guidance for stereotactic biopsy of Head
C1525263|Guidance for stereotactic biopsy:Find:Pt:Head:Doc:CT
C1525263|Guidance for stereotactic biopsy:Finding:Point in time:Head:Document:Computerized Tomography
C1525267|Multisection for calcium score^W contrast Intravenous:Finding:Point in time:Chest>Heart:Document:Computerized Tomography
C1525267|Multisection for calcium score^W contrast IV:Find:Pt:Chest>Heart:Doc:CT
C1525267|Hrt CT for Calcium Score W contr IV
C1525267|Heart CT for calcium scoring W contrast IV
C1525460|Humerus-L XR Transthoracic
C1525460|Humerus - left X-ray transthoracic
C1525460|View transthoracic:Find:Pt:Humerus.left:Doc:XR
C1525460|View transthoracic:Finding:Point in time:Humerus.left:Document:XR
C1525483|Wrist-L XR 5V
C1525483|Wrist - left X-ray 5 views
C1525483|Views 5:Finding:Point in time:Wrist.left:Document:XR
C1525483|Views 5:Find:Pt:Wrist.left:Doc:XR
C1525509|Patella-Bl XR AP+Lat+Sunrise
C1525509|Patella - bilateral X-ray AP and lateral and Sunrise
C1525509|Views AP & lateral & Sunrise:Find:Pt:Patella.bilateral:Doc:XR
C1525509|Views AP & lateral & Sunrise:Finding:Point in time:Patella.bilateral:Document:XR
C1525510|Patella-L XR AP+Lat+Sunrise
C1525510|Patella - left X-ray AP and lateral and Sunrise
C1525510|Views AP & lateral & Sunrise:Find:Pt:Patella.left:Doc:XR
C1525510|Views AP & lateral & Sunrise:Finding:Point in time:Patella.left:Document:XR
C1525523|Should-L XR AP+West Point
C1525523|Shoulder - left X-ray AP and West Point
C1525523|Views AP & West Point:Finding:Point in time:Shoulder.left:Document:XR
C1525523|Views AP & West Point:Find:Pt:Shoulder.left:Doc:XR
C1525562|Knee-Bl XR Sunrise+Tunnel
C1525562|Knee - bilateral X-ray Sunrise and tunnel
C1525562|Views Sunrise & tunnel:Find:Pt:Knee.bilateral:Doc:XR
C1525562|Views Sunrise & tunnel:Finding:Point in time:Knee.bilateral:Document:XR
C1525584|Views^W contrast IS:Find:Pt:Elbow.bilateral:Doc:XR.fluor
C1525584|Views^W contrast Intrasynovial:Finding:Point in time:Elbow.bilateral:Document:XR.fluor
C1525584|Elbow - bilateral Fluoroscopy W contrast IS
C1525584|Elbow-Bl Flr W contr IS
C1525648|L-spine+Sacrum XR 3V
C1525648|Spine Lumbar and Sacrum X-ray 3 views
C1525648|Views 3:Finding:Point in time:Spine.lumbar+Sacrum:Document:XR
C1525648|Views 3:Find:Pt:Spine.lumbar+Sacrum:Doc:XR
C1525671|Soft tissue MRI WO contrast
C1525671|Soft tissue MRI WO contr
C1525671|Multisection^WO contrast:Find:Pt:Soft tissue:Doc:MRI
C1525671|Multisection^WO contrast:Finding:Point in time:Soft tissue:Document:MRI
C1525689|L-spine+Sacrum XR
C1525689|Spine Lumbar and Sacrum X-ray
C1525689|Views:Find:Pt:Spine.lumbar+Sacrum:Doc:XR
C1525689|Views:Finding:Point in time:Spine.lumbar+Sacrum:Document:XR
C1525750|Wrist-L CT
C1525750|Wrist - left CT
C1525750|Multisection:Find:Pt:Wrist.left:Doc:CT
C1525750|Multisection:Finding:Point in time:Wrist.left:Document:Computerized Tomography
C1525754|Temporomandibular joint MRI cine
C1525754|TMJ MRI Cine
C1525754|Multisection cine:Finding:Point in time:Temporomandibular joint:Document:MRI
C1525754|Multisection cine:Find:Pt:Temporomandibular joint:Doc:MRI
C1525755|Brain MRI diffusion weighted
C1525755|Brain MRI Diff Wt
C1525755|Multisection diffusion weighted:Find:Pt:Brain:Doc:MRI
C1525755|Multisection diffusion weighted:Finding:Point in time:Brain:Document:MRI
C1524695|Wrist-Bl MRI W contr IV
C1524695|Wrist - bilateral MRI W contrast IV
C1524695|Multisection^W contrast IV:Find:Pt:Wrist.bilateral:Doc:MRI
C1524695|Multisection^W contrast Intravenous:Finding:Point in time:Wrist.bilateral:Document:MRI
C1525780|Shoulder - left X-ray Grashey
C1525780|Should-L XR Grashey
C1525780|View Grashey:Find:Pt:Shoulder.left:Doc:XR
C1525780|View Grashey:Finding:Point in time:Shoulder.left:Document:XR
C1525860|Thumb-L XR W Stress
C1525860|Thumb - left X-ray W manual stress
C1525860|Views^W manual stress:Finding:Point in time:Thumb.left:Document:XR
C1525860|Views^W manual stress:Find:Pt:Thumb.left:Doc:XR
C1525939|Pelvis XR AP+Obl
C1525939|Pelvis X-ray AP and oblique
C1525939|Views AP & oblique:Find:Pt:Pelvis:Doc:XR
C1525939|Views AP & oblique:Finding:Point in time:Pelvis:Document:XR
C1525820|Finger fifth - bilateral X-ray
C1525820|Finger.5th-Bl XR
C1525820|Views:Find:Pt:Finger.fifth.bilateral:Doc:XR
C1525820|Views:Finding:Point in time:Finger.fifth.bilateral:Document:XR
C1525951|Pelvis XR stand
C1525951|Pelvis X-ray standing
C1525951|View^standing:Finding:Point in time:Pelvis:Document:XR
C1525951|View^standing:Find:Pt:Pelvis:Doc:XR
C1525986|Ankle-R XR Lat+Mortise
C1525986|Ankle - right X-ray lateral and Mortise
C1525986|Views lateral & Mortise:Finding:Point in time:Ankle.right:Document:XR
C1525986|Views lateral & Mortise:Find:Pt:Ankle.right:Doc:XR
C1526130|Wrist-R XR 1V
C1526130|Wrist - right X-ray Single view
C1526130|View 1:Find:Pt:Wrist.right:Doc:XR
C1526130|View 1:Finding:Point in time:Wrist.right:Document:XR
C1526045|Hip-R XR Lat Frog
C1526045|Hip - right X-ray lateral frog
C1526045|View lateral frog:Find:Pt:Hip.right:Doc:XR
C1526045|View lateral frog:Finding:Point in time:Hip.right:Document:XR
C1526169|Spine X-ray AP single view
C1526169|Spine XR AP 1V
C1526169|View AP:Find:Pt:Spine:Doc:XR
C1526169|View AP:Finding:Point in time:Spine:Document:XR
C1524277|Thumb X-ray 3 views
C1524277|Thumb XR 3V
C1524277|Views 3:Find:Pt:Thumb:Doc:XR
C1524277|Views 3:Finding:Point in time:Thumb:Document:XR
C1526182|Toes X-ray 2 views
C1526182|Toes XR 2V
C1526182|Views 2:Find:Pt:Toes:Doc:XR
C1526182|Views 2:Finding:Point in time:Toes:Document:XR
C1524702|Wrist XR 1V
C1524702|Wrist X-ray Single view
C1524702|View 1:Finding:Point in time:Wrist:Document:XR
C1524702|View 1:Find:Pt:Wrist:Doc:XR
C1526244|Vertebral ves XRA W contr
C1526244|Vertebral vessels Fluoroscopic angiogram W contrast
C1526244|Views^W contrast:Find:Pt:Vertebral vessels:Doc:XR.fluor.angio
C1526244|Views^W contrast:Finding:Point in time:Vertebral vessels:Document:XR.fluor.angio
C1526259|US Guidance for fine needle aspiration of Unspecified body region
C1526259|XXX US FNA Asp
C1526259|Guidance for aspiration.fine needle:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1526259|Guidance for aspiration.fine needle:Find:Pt:XXX:Doc:US
C1526269|US Guidance for needle biopsy of Breast
C1526269|Brst US Bx needle guid
C1526269|Guidance for biopsy.needle:Finding:Point in time:Breast:Document:Ultrasound
C1526269|Guidance for biopsy.needle:Find:Pt:Breast:Doc:US
C1526333|Thoracic artery Fluoroscopic angiogram W contrast IA
C1526333|Thoracic a XRA W contr IA
C1526333|Views^W contrast Intra-arterial:Finding:Point in time:Thoracic artery:Document:XR.fluor.angio
C1526333|Views^W contrast IA:Find:Pt:Thoracic artery:Doc:XR.fluor.angio
C1526346|Submandibular gland Fluoroscopy W contrast intra salivary duct
C1526346|Submandib gland Flr W contr intra SD
C1526346|Views^W contrast intra salivary duct:Find:Pt:Submandibular gland:Doc:XR.fluor
C1526346|Views^W contrast intra salivary duct:Finding:Point in time:Submandibular gland:Document:XR.fluor
C1524483|Ankle-R CT W contr IV
C1524483|Ankle - right CT W contrast IV
C1524483|Multisection^W contrast IV:Find:Pt:Ankle.right:Doc:CT
C1524483|Multisection^W contrast Intravenous:Finding:Point in time:Ankle.right:Document:Computerized Tomography
C1524491|PA CT.Angio W contr IV
C1524491|Pulmonary artery CT angiogram W contrast IV
C1524491|Multisection^W contrast IV:Find:Pt:Pulmonary artery:Doc:CT.angio
C1524491|Multisection^W contrast Intravenous:Finding:Point in time:Pulmonary artery:Document:Computerized Tomography.angio
C1524503|Elbow-L CT W contr IV
C1524503|Elbow - left CT W contrast IV
C1524503|Multisection^W contrast IV:Find:Pt:Elbow.left:Doc:CT
C1524503|Multisection^W contrast Intravenous:Finding:Point in time:Elbow.left:Document:Computerized Tomography
C1524861|Forearm - right MRI WO contrast
C1524861|Forearm-R MRI WO contr
C1524861|Multisection^WO contrast:Finding:Point in time:Forearm.right:Document:MRI
C1524861|Multisection^WO contrast:Find:Pt:Forearm.right:Doc:MRI
C1524876|Upper arm CT WO contrast
C1524876|Upper arm CT WO contr
C1524876|Multisection^WO contrast:Find:Pt:Upper arm:Doc:CT
C1524876|Multisection^WO contrast:Finding:Point in time:Upper arm:Document:Computerized Tomography
C1524562|Knee-R MRI W contr IV
C1524562|Knee - right MRI W contrast IV
C1524562|Multisection^W contrast IV:Find:Pt:Knee.right:Doc:MRI
C1524562|Multisection^W contrast Intravenous:Finding:Point in time:Knee.right:Document:MRI
C1524566|Mandible CT W contr IV
C1524566|Mandible CT W contrast IV
C1524566|Multisection^W contrast Intravenous:Finding:Point in time:Mandible:Document:Computerized Tomography
C1524566|Multisection^W contrast IV:Find:Pt:Mandible:Doc:CT
C1524197|Knee - left X-ray Single view
C1524197|Knee-L XR 1V
C1524197|View 1:Find:Pt:Knee.left:Doc:XR
C1524197|View 1:Finding:Point in time:Knee.left:Document:XR
C1524216|Shoulder - bilateral X-ray AP single view
C1524216|Should-Bl XR AP 1V
C1524216|View AP:Finding:Point in time:Shoulder.bilateral:Document:XR
C1524216|View AP:Find:Pt:Shoulder.bilateral:Doc:XR
C1524282|Aorta Fluoroscopic angiogram Atherectomy W contrast IA
C1524282|Aorta XRA Atherect W contr IA
C1524282|Atherectomy^W contrast IA:Find:Pt:Aorta:Doc:XR.fluor.angio
C1524282|Atherectomy^W contrast Intra-arterial:Finding:Point in time:Aorta:Document:XR.fluor.angio
C1524290|Bone CT Bx guid
C1524290|CT Guidance for biopsy of Bone
C1524290|Guidance for biopsy:Finding:Point in time:Bone:Document:Computerized Tomography
C1524290|Guidance for biopsy:Find:Pt:Bone:Doc:CT
C1524608|Aorta thoracic MRI angiogram WO and W contrast IV
C1524608|Multisection^WO & W contrast IV:Find:Pt:Aorta.thoracic:Doc:MRI.angio
C1524608|Multisection^WO & W contrast Intravenous:Finding:Point in time:Aorta.thoracic:Document:MRI.angio
C1524608|TA MRI.Angio WO+W contr IV
C1524609|Multisection^WO & W contrast Intravenous:Finding:Point in time:Renal artery:Document:MRI.angio
C1524609|Renal artery MRI angiogram WO and W contrast IV
C1524609|Renal a MRI.Angio WO+W contr IV
C1524609|Multisection^WO & W contrast IV:Find:Pt:Renal artery:Doc:MRI.angio
C1524970|Hand - bilateral X-ray PA
C1524970|Hand-Bl XR PA V1
C1524970|View PA:Finding:Point in time:Hand.bilateral:Document:XR
C1524970|View PA:Find:Pt:Hand.bilateral:Doc:XR
C1524978|Hand-L XR
C1524978|Hand - left X-ray
C1524978|Views:Finding:Point in time:Hand.left:Document:XR
C1524978|Views:Find:Pt:Hand.left:Doc:XR
C1524347|Appendix CT
C1524347|Multisection:Finding:Point in time:Abdomen+Pelvis>Appendix:Document:Computerized Tomography
C1524347|Multisection:Find:Pt:Abdomen+Pelvis>Appendix:Doc:CT
C1525012|Toes - left X-ray 2 views
C1525012|Toes-L XR 2V
C1525012|Views 2:Find:Pt:Toes.left:Doc:XR
C1525012|Views 2:Finding:Point in time:Toes.left:Document:XR
C1524368|Lower extremity vessels - bilateral MRI angiogram
C1524368|Multisection:Finding:Point in time:Lower extremity vessels.bilateral:Document:MRI.angio
C1524368|Multisection:Find:Pt:Lower extremity vessels.bilateral:Doc:MRI.angio
C1524368|LE ves-Bl MRI.Angio
C1524372|Lower extremity - left MRI
C1524372|LE-L MRI
C1524372|Multisection:Finding:Point in time:Lower extremity.left:Document:MRI
C1524372|Multisection:Find:Pt:Lower extremity.left:Doc:MRI
C1524743|Multisection^WO & W contrast Intravenous:Finding:Point in time:Heart:Document:MRI
C1524743|Hrt MRI WO+W contr IV
C1524743|Heart MRI WO and W contrast IV
C1524743|Multisection^WO & W contrast IV:Find:Pt:Heart:Doc:MRI
C1524398|Hand-R CT
C1524398|Hand - right CT
C1524398|Multisection:Finding:Point in time:Hand.right:Document:Computerized Tomography
C1524398|Multisection:Find:Pt:Hand.right:Doc:CT
C1524404|Hip - bilateral X-ray tomograph
C1524404|Hip-Bl XRTomo
C1524404|Multisection:Finding:Point in time:Hip.bilateral:Document:XR.tomo
C1524404|Multisection:Find:Pt:Hip.bilateral:Doc:XR.tomo
C1524777|Sacrum+Coccyx MRI WO+W contr IV
C1524777|Sacrum and Coccyx MRI WO and W contrast IV
C1524777|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sacrum+Coccyx:Document:MRI
C1524777|Multisection^WO & W contrast IV:Find:Pt:Sacrum+Coccyx:Doc:MRI
C1524802|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity veins:Document:MRI.angio
C1524802|Upper extremity veins MRI angiogram WO and W contrast IV
C1524802|UE vv MRI.Angio WO+W contr IV
C1524802|Multisection^WO & W contrast IV:Find:Pt:Upper extremity veins:Doc:MRI.angio
C1524809|Abdomen CT WO contrast
C1524809|Abd CT WO contr
C1524809|Multisection^WO contrast:Find:Pt:Abdomen:Doc:CT
C1524809|Multisection^WO contrast:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524674|Thumb-L XR AP+Lat+Obl
C1524674|Thumb - left X-ray AP and lateral and oblique
C1524674|Views AP & lateral & oblique:Find:Pt:Thumb.left:Doc:XR
C1524674|Views AP & lateral & oblique:Finding:Point in time:Thumb.left:Document:XR
C1830200|Multisection:Finding:Point in time:Breast.unilateral:Narrative:MRI
C1830200|Brst-UL MRI
C1830200|Breast - unilateral MRI
C1830200|Multisection:Find:Pt:Breast.unilateral:Doc:MRI
C1830200|Multisection:Finding:Point in time:Breast.unilateral:Document:MRI
C1830262|Lung RI V W 133Xe IH
C1830262|Views ventilation^W Xe-133 IH:Find:Pt:Lung:Doc:Radnuc
C1830262|Lung Scan ventilation W Xe-133 IH
C1830262|Views ventilation^W Xe-133 Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1830278|Aorta US.doppler
C1830278|Aorta DOP
C1830278|Multisection:Find:Pt:Aorta:Doc:US.doppler
C1830278|Multisection:Finding:Point in time:Aorta:Document:Ultrasound.doppler
C1715399|Lower extremity vessels MRI angiogram WO contrast
C1715399|LE ves MRI.Angio WO contr
C1715399|Multisection^WO contrast:Find:Pt:Lower extremity vessels:Doc:MRI.angio
C1715399|Multisection^WO contrast:Finding:Point in time:Lower extremity vessels:Document:MRI.angio
C1715419|Hrt SPECT W Tc99mMIBI IV
C1715419|Heart SPECT W Tc-99m Sestamibi IV
C1715419|Multisection^W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1715419|Multisection^W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1715434|Guidance for drainage of abscess:Find:Pt:Pelvis:Doc:US
C1715434|Pelvis US Abscess drain guid
C1715434|US Guidance for drainage of abscess of Pelvis
C1715434|Guidance for drainage of abscess:Finding:Point in time:Pelvis:Document:Ultrasound
C1715441|Hip X-ray Single view portable
C1715441|Hip XR 1V port
C1715441|View 1 portable:Finding:Point in time:Hip:Document:XR
C1715441|View 1 portable:Find:Pt:Hip:Doc:XR
C1715455|Ribs+Chest XR GE 3V+PA Chst
C1715455|Ribs and Chest X-ray GE 3 and PA Chest views
C1715455|Views GE 3 & PA chest:Find:Pt:Ribs+Chest:Doc:XR
C1715455|Views GE 3 & PA chest:Finding:Point in time:Ribs+Chest:Document:XR
C1715465|Knee XR 1V or 2V Port
C1715465|Knee X-ray 1 or 2 views portable
C1715465|Views 1 or 2 portable:Find:Pt:Knee:Doc:XR
C1715465|Views 1 or 2 portable:Finding:Point in time:Knee:Document:XR
C1715483|Ovary Flr PC Abscess Drain guid
C1715483|Fluoroscopy Guidance for percutaneous drainage of abscess of Ovary
C1715483|Guidance for percutaneous drainage of abscess:Find:Pt:Ovary:Doc:XR.fluor
C1715483|Guidance for percutaneous drainage of abscess:Finding:Point in time:Ovary:Document:XR.fluor
C1715490|SM ves MRI.Angio WO contr
C1715490|Superior mesenteric vessels MRI angiogram WO contrast
C1715490|Multisection^WO contrast:Find:Pt:Superior mesenteric vessels:Doc:MRI.angio
C1715490|Multisection^WO contrast:Finding:Point in time:Superior mesenteric vessels:Document:MRI.angio
C1645319|Elbow-L XR Ltd
C1645319|Elbow - left X-ray limited
C1645319|Views limited:Find:Pt:Elbow.left:Doc:XR
C1645319|Views limited:Finding:Point in time:Elbow.left:Document:XR
C1648950|Bone RI Ltd W In-111 WBC IV
C1648950|Bone Scan limited W In-111 tagged WBC IV
C1648950|Views limited^W In-111 tagged WBC IV:Find:Pt:Bone:Doc:Radnuc
C1648950|Views limited^W In-111 tagged WBC Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1714803|Chest X-ray AP right lateral-decubitus
C1714803|Chest XR AP R-Lat Decub
C1714803|View AP R-lateral-decubitus:Find:Pt:Chest:Doc:XR
C1714803|View AP R-lateral-decubitus:Finding:Point in time:Chest:Document:XR
C1714808|Unspecified body region Fluoroscopy 2 hour
C1714808|XXX Flr 2h
C1714808|View:Finding:2 hours:To be specified in another part of the message:Document:XR.fluor
C1714808|View:Find:2H:XXX:Doc:XR.fluor
C1714810|BD+PDs Flr Endo guid 2h P contr retro
C1714810|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 2 hours post contrast retrograde
C1714810|Guidance for endoscopy^2H post contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1714810|Guidance for endoscopy^2 hours post contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1714908|Thymus gland MRI
C1714908|Thymus MRI
C1714908|Multisection:Finding:Point in time:Thymus gland:Document:MRI
C1714908|Multisection:Find:Pt:Thymus gland:Doc:MRI
C1714951|Skeletal Sys Periph RI BDM
C1714951|Skeletal system.peripheral Scan Bone density
C1714951|Bone density:Find:Pt:Skeletal system.peripheral:Doc:Radnuc
C1714951|Bone density:Finding:Point in time:Skeletal system.peripheral:Document:Radnuc
C1715033|Renal vessels Scan
C1715033|Renal ves RI W RNC IV
C1715033|Views^W radionuclide IV:Find:Pt:Renal vessels:Doc:Radnuc
C1715033|Views^W radionuclide Intravenous:Finding:Point in time:Renal vessels:Document:Radnuc
C1714508|Brst-R US Localization guid
C1714508|US Guidance for localization of Breast - right
C1714508|Guidance for localization:Find:Pt:Breast.right:Doc:US
C1714508|Guidance for localization:Finding:Point in time:Breast.right:Document:Ultrasound
C1715095|Kidney - bilateral CT
C1715095|Multisection:Find:Pt:Kidney.bilateral:Doc:CT
C1715095|Multisection:Finding:Point in time:Kidney.bilateral:Document:Computerized Tomography
C1715095|Kdny-Bl CT
C1631281|Knee-R XR Sunrise+(views Stand)
C1631281|Knee - right X-ray Sunrise and (views standing)
C1631281|View Sunrise & (views^standing):Finding:Point in time:Knee.right:Document:XR
C1631281|View Sunrise & (views^standing):Find:Pt:Knee.right:Doc:XR
C1637285|T-spine XR 3V stand
C1637285|Views 3^standing:Find:Pt:Spine.thoracic:Doc:XR
C1637285|Views 3^standing:Finding:Point in time:Spine.thoracic:Document:XR
C1637285|Thoracic spine X-ray 3 views standing
C1645333|T-spine XR AP W+WO R+L-bending
C1645333|Views AP^W R-bending & W L-bending & WO bending:Find:Pt:Spine.thoracic:Doc:XR
C1645333|Views AP^W R-bending & W L-bending & WO bending:Finding:Point in time:Spine.thoracic:Document:XR
C1645333|Thoracic spine X-ray AP W right bending and W left bending and WO bending
C1632361|Mastoid - bilateral X-ray limited
C1632361|Mastoid-Bl XR Ltd
C1632361|Views limited:Find:Pt:Mastoid.bilateral:Doc:XR
C1632361|Views limited:Finding:Point in time:Mastoid.bilateral:Document:XR
C1623576|Bladder+Urethra Flr W contr
C1623576|Urinary Bladder and Urethra Fluoroscopy W contrast
C1623576|Views^W contrast:Finding:Point in time:Urinary bladder+Urethra:Document:XR.fluor
C1623576|Views^W contrast:Find:Pt:Urinary bladder+Urethra:Doc:XR.fluor
C1637229|Guidance for superficial biopsy:Finding:Point in time:Bone:Document:Ultrasound
C1637229|US Guidance for superficial biopsy of Bone
C1637229|Bone US Bx super guid
C1637229|Guidance for superficial biopsy:Find:Pt:Bone:Doc:US
C1639909|Adrenal gland Scan
C1639909|Adrenal RI W RNC IV
C1639909|Views^W radionuclide Intravenous:Finding:Point in time:Adrenal gland:Narrative:Radnuc
C1639909|Views^W radionuclide Intravenous:Finding:Point in time:Adrenal gland:Document:Radnuc
C1639909|Views^W radionuclide IV:Find:Pt:Adrenal gland:Doc:Radnuc
C1630174|CT Guidance for superficial needle biopsy of Bone
C1630174|Guidance for superficial biopsy.needle:Find:Pt:Bone:Doc:CT
C1630174|Guidance for superficial biopsy.needle:Finding:Point in time:Bone:Document:Computerized Tomography
C1630174|Bone CT Bx super need guid
C1642085|GB RI W CCK+RNC IV
C1642085|Gallbladder Scan W cholecystokinin and W radionuclide IV
C1642085|Views^W cholecystokinin & W radionuclide IV:Find:Pt:Gallbladder:Doc:Radnuc
C1642085|Views^W cholecystokinin & W radionuclide Intravenous:Finding:Point in time:Gallbladder:Document:Radnuc
C1630179|Guidance for drainage:Finding:Point in time:Abdomen>Retroperitoneum:Document:Computerized Tomography
C1630179|CT Guidance for drainage of Retroperitoneum
C1630179|Retroperitoneum CT Drain guid
C1630179|Guidance for drainage:Find:Pt:Abdomen>Retroperitoneum:Doc:CT
C1632228|Guidance for placement of infusion port:Find:Pt:Hepatic artery:Nar:Radnuc
C1632228|Guidance for placement of infusion port:Finding:Point in time:Hepatic artery:Narrative:Radnuc
C1632228|Deprecated Scan Guidance for placement of infusion port in Hepatic artery
C1632228|Deprecated Hep a RI Infusion port plac g
C1632230|Orbit - right X-ray for foreign body
C1632230|Orbit-R XR for FB
C1632230|Views for foreign body:Finding:Point in time:Orbit.right:Document:XR
C1632230|Views for foreign body:Find:Pt:Orbit.right:Doc:XR
C1624697|Lower leg - bilateral MRI
C1624697|Lower leg-Bl MRI
C1624697|Multisection:Finding:Point in time:Lower leg.bilateral:Document:MRI
C1624697|Multisection:Find:Pt:Lower leg.bilateral:Doc:MRI
C1954314|TMJ-Ul XR Open+Closed Mouth
C1954314|Temporomandibular Joint - unilateral X-ray open and closed mouth
C1954314|Views open & closed mouth:Find:Pt:Temporomandibular joint.unilateral:Doc:XR
C1954314|Views open & closed mouth:Finding:Point in time:Temporomandibular joint.unilateral:Document:XR
C1953970|Views:Finding:Point in time:Trachea:Narrative:XR.fluor
C1953970|Trachea Fluoroscopy
C1953970|Trachea Flr
C1953970|Views:Find:Pt:Trachea:Doc:XR.fluor
C1953970|Views:Finding:Point in time:Trachea:Document:XR.fluor
C2598763|CT Cerebral atrophic index
C2598763|CT VFr Cerebral atrophic index
C2598763|Cerebral atrophic index:VFr:Pt:^Patient:Qn:CT
C2598763|Cerebral atrophic index:Volume Fraction:Point in time:^Patient:Quantitative:Computerized Tomography
C3174368|Kidney-R Flr View for cyst exam
C3174368|Kidney - right Fluoroscopy View for cyst examination
C3174368|View for cyst examination:Find:Pt:Kidney.right:Doc:XR.fluor
C3174368|View for cyst examination:Finding:Point in time:Kidney.right:Document:XR.fluor
C3533904|Multisection screening:Find:Pt:Breast.left:Doc:Mam.FFD.tomosynthesis
C3533904|Brst-L FFDM-DBT Screening
C3533904|Breast - left FFD mammogram-tomosynthesis screening
C3533904|Multisection screening:Finding:Point in time:Breast.left:Document:Mam.FFD.tomosynthesis
C3262991|Elbow - bilateral MRI WO contrast
C3262991|Elbow-Bl MRI WO contr
C3262991|Multisection^WO contrast:Finding:Point in time:Elbow.bilateral:Document:MRI
C3262991|Multisection^WO contrast:Find:Pt:Elbow.bilateral:Doc:MRI
C3263003|Upper arm - bilateral MRI WO contrast
C3263003|Upper arm-Bl MRI WO contr
C3263003|Multisection^WO contrast:Find:Pt:Upper arm.bilateral:Doc:MRI
C3263003|Multisection^WO contrast:Finding:Point in time:Upper arm.bilateral:Document:MRI
C3482439|L-spine Flr PC Vertebroplasty guid
C3482439|Guidance for percutaneous vertebroplasty:Find:Pt:Spine.lumbar:Doc:XR.fluor
C3482439|Guidance for percutaneous vertebroplasty:Finding:Point in time:Spine.lumbar:Document:XR.fluor
C3482439|Fluoroscopy Guidance for percutaneous vertebroplasty of Lumbar spine
C3263032|Wrist - right and Hand - right MRI
C3263032|Wrist+Hand-R MRI
C3263032|Multisection:Find:Pt:Wrist.right+Hand.right:Doc:MRI
C3263032|Multisection:Finding:Point in time:Wrist.right+Hand.right:Document:MRI
C3263085|Spine thoracolumbar junction XR 2V
C3263085|Spine Thoracolumbar Junction X-ray 2 views
C3263085|Views 2:Find:Pt:Spine.thoracolumbar junction:Doc:XR
C3263085|Views 2:Finding:Point in time:Spine.thoracolumbar junction:Document:XR
C3481961|Multisection^W contrast IV:Find:Pt:Abdomen+Pelvis>Vessels:Doc:CT.angio
C3481961|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis>Vessels:Document:Computerized Tomography.angio
C3481961|Abd+Pelvis>ves CT.Angio W contr IV
C3481961|Abdominal and Pelvic Vessels CT angiogram W contrast IV
C0800894|Thyroid Scan Study report
C0800894|Thyroid RI Study report
C0800894|Study report:Find:Pt:Thyroid:Doc:Radnuc
C0800894|Study report:Finding:Point in time:Thyroid:Document:Radnuc
C0944197|Liver US
C0944197|Multisection:Find:Pt:Liver:Doc:US
C0944197|Multisection:Finding:Point in time:Liver:Document:Ultrasound
C0944734|Chest CT WO contr
C0944734|Chest CT WO contrast
C0944734|Multisection^WO contrast:Find:Pt:Chest:Doc:CT
C0944734|Multisection^WO contrast:Finding:Point in time:Chest:Document:Computerized Tomography
C0942152|Mastoid - left X-ray
C0942152|Mastoid-L XR
C0942152|Views:Finding:Point in time:Mastoid.left:Document:XR
C0942152|Views:Find:Pt:Mastoid.left:Doc:XR
C0942269|Multisection:Finding:Point in time:Thigh.left:Narrative:MRI
C0942269|Thigh - left MRI
C0942269|Thigh-L MRI
C0942269|Multisection:Find:Pt:Thigh.left:Doc:MRI
C0942269|Multisection:Finding:Point in time:Thigh.left:Document:MRI
C0942273|Wrist - left MRI
C0942273|Wrist-L MRI
C0942273|Multisection:Finding:Point in time:Wrist.left:Document:MRI
C0942273|Multisection:Find:Pt:Wrist.left:Doc:MRI
C0942275|Wrist - right MRI
C0942275|Wrist-R MRI
C0942275|Multisection:Finding:Point in time:Wrist.right:Document:MRI
C0942275|Multisection:Find:Pt:Wrist.right:Doc:MRI
C0942287|Cent v-Bl XRA Cath repos W contr IV
C0942287|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - bilateral-- W contrast IV
C0942287|Guidance for reposition of catheter^W contrast IV:Find:Pt:Central vein.bilateral:Doc:XR.fluor.angio
C0942287|Guidance for reposition of catheter^W contrast Intravenous:Finding:Point in time:Central vein.bilateral:Document:XR.fluor.angio
C0945337|Cent v-Bl XRA Cath plac guid W contr IV
C0945337|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - bilateral-- W contrast IV
C0945337|Guidance for placement of catheter^W contrast IV:Find:Pt:Central vein.bilateral:Doc:XR.fluor.angio
C0945337|Guidance for placement of catheter^W contrast Intravenous:Finding:Point in time:Central vein.bilateral:Document:XR.fluor.angio
C0942352|Iliac a-R XRA Angpsty W contr IA
C0942352|Iliac artery - right Fluoroscopic angiogram Angioplasty W contrast IA
C0942352|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Iliac artery.right:Document:XR.fluor.angio
C0942352|Angioplasty^W contrast IA:Find:Pt:Iliac artery.right:Doc:XR.fluor.angio
C0942374|Patella - bilateral X-ray 2 views
C0942374|Patella-Bl XR 2V
C0942374|Views 2:Finding:Point in time:Patella.bilateral:Document:XR
C0942374|Views 2:Find:Pt:Patella.bilateral:Doc:XR
C0882031|Neck CT Asp guid
C0882031|CT Guidance for aspiration of Neck
C0882031|Guidance for aspiration:Finding:Point in time:Neck:Document:Computerized Tomography
C0882031|Guidance for aspiration:Find:Pt:Neck:Doc:CT
C0882050|Pancreas CT
C0882050|Multisection:Finding:Point in time:Pancreas:Narrative:Computerized Tomography
C0882050|Multisection:Find:Pt:Abdomen>Pancreas:Doc:CT
C0882050|Multisection:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C0882053|Panc a XRA W contr IA
C0882053|Pancreatic artery Fluoroscopic angiogram W contrast IA
C0882053|Views^W contrast IA:Find:Pt:Pancreatic artery:Doc:XR.fluor.angio
C0882053|Views^W contrast Intra-arterial:Finding:Point in time:Pancreatic artery:Document:XR.fluor.angio
C0882107|Spinal a XRA W contr IA
C0882107|Spinal artery Fluoroscopic angiogram W contrast IA
C0882107|Views^W contrast IA:Find:Pt:Spinal artery:Doc:XR.fluor.angio
C0882107|Views^W contrast Intra-arterial:Finding:Point in time:Spinal artery:Document:XR.fluor.angio
C0882115|Multisection:Finding:Point in time:Spine.cervical:Narrative:MRI
C0882115|C-spine MRI
C0882115|Multisection:Find:Pt:Spine.cervical:Doc:MRI
C0882115|Multisection:Finding:Point in time:Spine.cervical:Document:MRI
C0882115|Cervical spine MRI
C0882129|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.lumbar:Document:MRI
C0882129|Multisection^WO & W contrast IV:Find:Pt:Spine.lumbar:Doc:MRI
C0882129|L-spine MRI WO+W contr IV
C0882129|Lumbar spine MRI WO and W contrast IV
C0882146|Spine CT Bx guid
C0882146|CT Guidance for biopsy of Spine
C0882146|Guidance for biopsy:Finding:Point in time:Spine:Document:Computerized Tomography
C0882146|Guidance for biopsy:Find:Pt:Spine:Doc:CT
C0884114|Fluoroscopy Guidance for placement of stent in Intrahepatic portal system
C0884114|IHP Flr Stent plac guid
C0884114|Guidance for placement of stent:Find:Pt:Intrahepatic portal system:Doc:XR.fluor
C0884114|Guidance for placement of stent:Finding:Point in time:Intrahepatic portal system:Document:XR.fluor
C0942096|Knee - left Fluoroscopy W contrast IS
C0942096|Knee-L Flr W contr IS
C0942096|Views^W contrast Intrasynovial:Finding:Point in time:Knee.left:Document:XR.fluor
C0942096|Views^W contrast IS:Find:Pt:Knee.left:Doc:XR.fluor
C0942119|Ankle - right X-ray
C0942119|Ankle-R XR
C0942119|Views:Finding:Point in time:Ankle.right:Document:XR
C0942119|Views:Find:Pt:Ankle.right:Doc:XR
C0881786|Aorta US
C0881786|Multisection:Finding:Point in time:Aorta:Document:Ultrasound
C0881786|Multisection:Find:Pt:Aorta:Doc:US
C0881835|Brst US Needle local guid
C0881835|US Guidance for needle localization of Breast
C0881835|Guidance for needle localization:Finding:Point in time:Breast:Document:Ultrasound
C0881835|Guidance for needle localization:Find:Pt:Breast:Doc:US
C0881841|Breast Mammogram screening
C0881841|Brst Mam Screening
C0881841|Views screening:Find:Pt:Breast:Doc:Mam
C0881841|Views screening:Finding:Point in time:Breast:Document:Mam
C0881896|Fluoroscopy Guidance for aspiration of cyst of Unspecified body region
C0881896|XXX Flr Cyst Asp guid
C0881896|Guidance for aspiration of cyst:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C0881896|Guidance for aspiration of cyst:Find:Pt:XXX:Doc:XR.fluor
C0881899|Elbow MRI
C0881899|Multisection:Finding:Point in time:Elbow:Narrative:MRI
C0881899|Multisection:Find:Pt:Elbow:Doc:MRI
C0881899|Multisection:Finding:Point in time:Elbow:Document:MRI
C0881947|Multisection^WO & W contrast IV:Find:Pt:Head:Doc:CT.perfusion
C0881947|Head CT perfusion WO and W contrast IV
C0881947|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head:Document:Computerized Tomography.perfusion
C0881947|Head CT.perfusion WO+W contr IV
C0882539|Knee MRI
C0882539|Multisection:Finding:Point in time:Knee:Narrative:MRI
C0882539|Multisection:Finding:Point in time:Knee:Document:MRI
C0882539|Multisection:Find:Pt:Knee:Doc:MRI
C1114932|Prostate MRI
C1114932|Multisection:Finding:Point in time:Prostate:Document:MRI
C1114932|Multisection:Find:Pt:Prostate:Doc:MRI
C1114500|L-spine MRI WO contr
C1114500|Multisection^WO contrast:Find:Pt:Spine.lumbar:Doc:MRI
C1114500|Multisection^WO contrast:Finding:Point in time:Spine.lumbar:Document:MRI
C1114500|Lumbar spine MRI WO contrast
C1114505|Hand MRI WO contr
C1114505|Hand MRI WO contrast
C1114505|Multisection^WO contrast:Finding:Point in time:Hand:Document:MRI
C1114505|Multisection^WO contrast:Find:Pt:Hand:Doc:MRI
C1114535|Sinuses XR PA+Lat
C1114535|Sinuses X-ray PA and lateral
C1114535|Views PA & lateral:Finding:Point in time:Sinuses:Document:XR
C1114535|Views PA & lateral:Find:Pt:Sinuses:Doc:XR
C1114557|Views:Finding:Point in time:Chest:Narrative:XR
C1114557|Chest X-ray
C1114557|Chest XR
C1114557|Views:Find:Pt:Chest:Doc:XR
C1114557|Views:Finding:Point in time:Chest:Document:XR
C1114943|Abd XRTomo
C1114943|Abdomen X-ray tomograph
C1114943|Multisection:Finding:Point in time:Abdomen:Document:XR.tomo
C1114943|Multisection:Find:Pt:Abdomen:Doc:XR.tomo
C1114613|Posterior fossa Fluoroscopy W contrast IT
C1114613|Post fossa Flr W contr IT
C1114613|Views^W contrast Intrathecal:Finding:Point in time:Posterior fossa:Document:XR.fluor
C1114613|Views^W contrast IT:Find:Pt:Posterior fossa:Doc:XR.fluor
C1114635|Visceral artery Fluoroscopic angiogram Angioplasty W contrast IA
C1114635|Visceral a XRA Angpsty W contr IA
C1114635|Angioplasty^W contrast IA:Find:Pt:Visceral artery:Doc:XR.fluor.angio
C1114635|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Visceral artery:Document:XR.fluor.angio
C1114674|Guidance for drainage:Find:Pt:XXX:Nar:US
C1114674|Deprecated XXX US Drain guid
C1114674|Deprecated Unspecified system US Guidance for drainage
C1114674|Guidance for drainage:Finding:Point in time:To be specified in another part of the message:Narrative:Ultrasound
C1114674|Deprecated XXX US Guid for drain
C1114437|CT Guidance for biopsy of Spleen
C1114437|Spleen CT Bx guid
C1114437|Guidance for biopsy:Find:Pt:Abdomen>Spleen:Doc:CT
C1114437|Guidance for biopsy:Finding:Point in time:Abdomen>Spleen:Document:Computerized Tomography
C1114450|Spleen CT W contr IV
C1114450|Spleen CT W contrast IV
C1114450|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen>Spleen:Document:Computerized Tomography
C1114450|Multisection^W contrast IV:Find:Pt:Abdomen>Spleen:Doc:CT
C1114453|Lower extremity CT WO contrast
C1114453|LE CT WO contr
C1114453|Multisection^WO contrast:Finding:Point in time:Lower extremity:Document:Computerized Tomography
C1114453|Multisection^WO contrast:Find:Pt:Lower extremity:Doc:CT
C1114466|Vein XRA Add'l Angpsty W contr IV
C1114466|Vein Fluoroscopic angiogram Additional angioplasty W contrast IV
C1114466|Angioplasty.additional^W contrast IV:Find:Pt:Vein:Doc:XR.fluor.angio
C1114466|Angioplasty.additional^W contrast Intravenous:Finding:Point in time:Vein:Document:XR.fluor.angio
C1526821|Carot a+Cerebral a Int-L XRA W contr IA
C1526821|Carotid artery and Cerebral artery internal - left Fluoroscopic angiogram W contrast IA
C1526821|Views^W contrast IA:Find:Pt:Carotid artery+Cerebral artery internal.left:Doc:XR.fluor.angio
C1526821|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Cerebral artery internal.left:Document:XR.fluor.angio
C1526825|Ribs post-L XR
C1526825|Ribs posterior - left X-ray
C1526825|Views:Find:Pt:Ribs.posterior.left:Doc:XR
C1526825|Views:Finding:Point in time:Ribs.posterior.left:Document:XR
C1526830|Tib+Fib-L XR 2V Obl
C1526830|Tibia - left and Fibula - left X-ray 2 views Oblique
C1526830|Views 2 oblique:Finding:Point in time:Tibia.left+Fibula.left:Document:XR
C1526830|Views 2 oblique:Find:Pt:Tibia.left+Fibula.left:Doc:XR
C1543422|Should-Bl XR AP(w IR+ER)+Ax+Outlet
C1543422|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary and outlet
C1543422|Views AP (W internal rotation & W external rotation) & axillary & outlet:Find:Pt:Shoulder.bilateral:Doc:XR
C1543422|Views AP (W internal rotation & W external rotation) & axillary & outlet:Finding:Point in time:Shoulder.bilateral:Document:XR
C1543428|Should-Bl XR AP(w IR+ER)+Y
C1543428|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and Y
C1543428|Views AP (W internal rotation & W external rotation) & Y:Find:Pt:Shoulder.bilateral:Doc:XR
C1543428|Views AP (W internal rotation & W external rotation) & Y:Finding:Point in time:Shoulder.bilateral:Document:XR
C1543429|Should-Bl XR AP(w IR+ER)+Ax+Y
C1543429|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary and Y
C1543429|Views AP (W internal rotation & W external rotation) & axillary & Y:Find:Pt:Shoulder.bilateral:Doc:XR
C1543429|Views AP (W internal rotation & W external rotation) & axillary & Y:Finding:Point in time:Shoulder.bilateral:Document:XR
C1543740|RI Ltd W Ga-67 IV
C1543740|Views limited^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543740|Views limited^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543740|Scan limited W Ga-67 IV
C1543770|Hrt SPECT PF Rest+W RNC IV
C1543770|Heart SPECT perfusion at rest and W radionuclide IV
C1543770|Multisection perfusion^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543770|Multisection perfusion^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543476|Wrist-R XR 3V+Carpal Tunnel
C1543476|Wrist - right X-ray 3 views and carpal tunnel
C1543476|Views 3 & carpal tunnel:Find:Pt:Wrist.right:Doc:XR
C1543476|Views 3 & carpal tunnel:Finding:Point in time:Wrist.right:Document:XR
C1543480|Should XR Ax+Transcapular
C1543480|Shoulder X-ray axillary and transcapular
C1543480|Views axillary & transcapular:Finding:Point in time:Shoulder:Document:XR
C1543480|Views axillary & transcapular:Find:Pt:Shoulder:Doc:XR
C1543485|T-spine XRTomo AP
C1543485|Multisection AP:Finding:Point in time:Spine.thoracic:Document:XR.tomo
C1543485|Multisection AP:Find:Pt:Spine.thoracic:Doc:XR.tomo
C1543485|Thoracic spine X-ray tomograph AP
C1543884|Views static^W Tc-99m DMSA Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1543884|Views static^W Tc-99m DMSA IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1543884|Kidney - bilateral Scan static W Tc-99m DMSA IV
C1543884|Kdny-Bl RI Static W Tc99mDMCA IV
C1543926|Bone Scan multiple areas
C1543926|Bone RI Mul Areas W RNC IV
C1543926|Views multiple areas^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543926|Views multiple areas^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543933|Deprecated Heart Scan first pass & wall motion & ejection fraction single view
C1543933|Deprecated Hrt RI FP+WM+EF V1 W RNC IV
C1543933|View first pass & wall motion & ejection fraction^W radionuclide IV:Find:Pt:Heart:Nar:Radnuc
C1543933|View first pass & wall motion & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1543942|Hrt RI Gated Rest+W Tc99mMIBI IV
C1543942|Heart Scan gated at rest and W Tc-99m Sestamibi IV
C1543942|Views gated^at rest & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543942|Views gated^at rest & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543958|Views ventilation^W radionuclide gaseous IH single breath:Find:Pt:Lung:Doc:Radnuc
C1543958|Views ventilation^W radionuclide gaseous Inhalation single breath:Finding:Point in time:Lung:Document:Radnuc
C1543958|Lung RI V W RNC Gas IH SB
C1543958|Lung Scan ventilation W radionuclide gaseous IH single breath
C1543511|Renal a DOP
C1543511|Renal artery US.doppler
C1543511|Multisection:Find:Pt:Renal artery:Doc:US.doppler
C1543511|Multisection:Finding:Point in time:Renal artery:Document:Ultrasound.doppler
C1543156|Deprecated Multisection:Find:Pt:XXX:Nar:US
C1543156|Deprecated XXX US
C1543156|Multisection:Find:Pt:XXX:Nar:US
C1543156|Deprecated Unspecified system US Multisection
C1543156|Multisection:Finding:Point in time:To be specified in another part of the message:Narrative:Ultrasound
C1525163|Internal auditory canal - right CT
C1525163|IAC-R CT
C1525163|Multisection:Finding:Point in time:Internal auditory canal.right:Document:Computerized Tomography
C1525163|Multisection:Find:Pt:Internal auditory canal.right:Doc:CT
C1542862|Vas Deferens Flr W contr intra VD
C1542862|Vas deferens Fluoroscopy W contrast intra vas deferens
C1542862|Views^W contrast intra vas deferens:Find:Pt:Vas deferens:Doc:XR.fluor
C1542862|Views^W contrast intra vas deferens:Finding:Point in time:Vas deferens:Document:XR.fluor
C1543689|Bone Scan limited
C1543689|Bone RI Ltd W RNC IV
C1543689|Views limited^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543689|Views limited^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543700|Brain SPECT W I-123 IV
C1543700|Multisection^W I-123 IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1543700|Multisection^W I-123 Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1543727|Heart Scan for shunt detection
C1543727|Hrt RI for Shunt Det W RNC IV
C1543727|Views for shunt detection^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543727|Views for shunt detection^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1524430|Knee - right CT
C1524430|Knee-R CT
C1524430|Multisection:Finding:Point in time:Knee.right:Document:Computerized Tomography
C1524430|Multisection:Find:Pt:Knee.right:Doc:CT
C1527050|Liver MRI
C1527050|Multisection:Finding:Point in time:Liver:Narrative:MRI
C1527050|Multisection:Find:Pt:Liver:Doc:MRI
C1527050|Multisection:Finding:Point in time:Liver:Document:MRI
C1527071|Shoulder CT
C1527071|Should CT
C1527071|Multisection:Finding:Point in time:Shoulder:Document:Computerized Tomography
C1527071|Multisection:Find:Pt:Shoulder:Doc:CT
C1524187|Lower leg - left MRI
C1524187|Lower leg-L MRI
C1524187|Multisection:Find:Pt:Lower leg.left:Doc:MRI
C1524187|Multisection:Finding:Point in time:Lower leg.left:Document:MRI
C1524830|Elbow-L CT WO contr
C1524830|Elbow - left CT WO contrast
C1524830|Multisection^WO contrast:Find:Pt:Elbow.left:Doc:CT
C1524830|Multisection^WO contrast:Finding:Point in time:Elbow.left:Document:Computerized Tomography
C1524444|Chest CT Ltd
C1524444|Chest CT limited
C1524444|Multisection limited:Find:Pt:Chest:Doc:CT
C1524444|Multisection limited:Finding:Point in time:Chest:Document:Computerized Tomography
C1525295|Should-Bl XR Ax
C1525295|Shoulder - bilateral X-ray axillary
C1525295|View axillary:Find:Pt:Shoulder.bilateral:Doc:XR
C1525295|View axillary:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525196|Orbit-L MRI W contr IV
C1525196|Orbit - left MRI W contrast IV
C1525196|Multisection^W contrast IV:Find:Pt:Orbit.left:Doc:MRI
C1525196|Multisection^W contrast Intravenous:Finding:Point in time:Orbit.left:Document:MRI
C1525204|Carot ves MRI.Angio W contr IV
C1525204|Carotid vessel MRI angiogram W contrast IV
C1525204|Multisection^W contrast IV:Find:Pt:Carotid vessel:Doc:MRI.angio
C1525204|Multisection^W contrast Intravenous:Finding:Point in time:Carotid vessel:Document:MRI.angio
C1525229|Multisection^WO & W contrast IV:Find:Pt:Abdominal vessels:Doc:MRI.angio
C1525229|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdominal vessels:Document:MRI.angio
C1525229|Abd ves MRI.Angio WO+W contr IV
C1525229|Abdominal vessels MRI angiogram WO and W contrast IV
C1525232|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity vessels.left:Document:MRI.angio
C1525232|Lower extremity vessels - left MRI angiogram WO and W contrast IV
C1525232|Multisection^WO & W contrast IV:Find:Pt:Lower extremity vessels.left:Doc:MRI.angio
C1525232|LE ves-L MRI.Angio WO+W contr IV
C1525236|Knee vessels - right MRI angiogram WO and W contrast IV
C1525236|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee vessels.right:Document:MRI.angio
C1525236|Multisection^WO & W contrast IV:Find:Pt:Knee vessels.right:Doc:MRI.angio
C1525236|Knee ves-R MRI.Angio WO+W contr IV
C1525244|UE joint-R MRI WO contr
C1525244|Upper extremity joint - right MRI WO contrast
C1525244|Multisection^WO contrast:Finding:Point in time:Upper extremity.joint.right:Document:MRI
C1525244|Multisection^WO contrast:Find:Pt:Upper extremity.joint.right:Doc:MRI
C1525257|Orbit-L XR
C1525257|Orbit - left X-ray
C1525257|Views:Find:Pt:Orbit.left:Doc:XR
C1525257|Views:Finding:Point in time:Orbit.left:Document:XR
C1525270|Maxillofacial CT Ltd WO contr
C1525270|Maxillofacial region CT limited WO contrast
C1525270|Multisection limited^WO contrast:Find:Pt:Head>Maxillofacial region:Doc:CT
C1525270|Multisection limited^WO contrast:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1525499|Pelvis+Hip-L XR AP+Lat Xtable
C1525499|Pelvis and Hip - left X-ray AP and lateral crosstable
C1525499|Views AP & lateral crosstable:Finding:Point in time:Pelvis+Hip.left:Document:XR
C1525499|Views AP & lateral crosstable:Find:Pt:Pelvis+Hip.left:Doc:XR
C1525610|CT Guidance for superficial biopsy of Tissue
C1525610|tiss CT Bx super guid
C1525610|Guidance for superficial biopsy:Finding:Point in time:Tissue:Document:Computerized Tomography
C1525610|Guidance for superficial biopsy:Find:Pt:Tissue:Doc:CT
C1525619|Multisection:Finding:Point in time:Parotid gland:Narrative:MRI
C1525619|Parotid gland MRI
C1525619|Multisection:Find:Pt:Parotid gland:Doc:MRI
C1525619|Multisection:Finding:Point in time:Parotid gland:Document:MRI
C1525664|Sternoclavicular Joint CT WO contrast
C1525664|SC joint CT WO contr
C1525664|Multisection^WO contrast:Finding:Point in time:Sternoclavicular joint:Document:Computerized Tomography
C1525664|Multisection^WO contrast:Find:Pt:Sternoclavicular joint:Doc:CT
C1525676|Sternoclavicular joint - left X-ray Serendipity
C1525676|SC joint-L XR Serendipity
C1525676|View Serendipity:Finding:Point in time:Sternoclavicular joint.left:Document:XR
C1525676|View Serendipity:Find:Pt:Sternoclavicular joint.left:Doc:XR
C1525694|Pelvis+L-spine XR 5V
C1525694|Pelvis and Spine Lumbar X-ray 5 views
C1525694|Views 5:Find:Pt:Pelvis+Spine.lumbar:Doc:XR
C1525694|Views 5:Finding:Point in time:Pelvis+Spine.lumbar:Document:XR
C1525743|IM v XRA W contr IV
C1525743|Inferior mesenteric vein Fluoroscopic angiogram W contrast IV
C1525743|Views^W contrast Intravenous:Finding:Point in time:Inferior mesenteric vein:Document:XR.fluor.angio
C1525743|Views^W contrast IV:Find:Pt:Inferior mesenteric vein:Doc:XR.fluor.angio
C1525744|Orbit vv-L XRA W contr IV
C1525744|Orbit veins - left Fluoroscopic angiogram W contrast IV
C1525744|Views^W contrast Intravenous:Finding:Point in time:Orbit veins.left:Document:XR.fluor.angio
C1525744|Views^W contrast IV:Find:Pt:Orbit veins.left:Doc:XR.fluor.angio
C1525759|Lung parenchyma CT W contr IV
C1525759|Multisection^W contrast IV:Find:Pt:Chest>Lung parenchyma:Doc:CT
C1525759|Lung parenchyma CT W contrast IV
C1525759|Multisection^W contrast Intravenous:Finding:Point in time:Chest>Lung parenchyma:Document:Computerized Tomography
C1525775|Shoulder - bilateral X-ray 30 degree caudal angle
C1525775|Should-Bl XR 30 Deg Cau Angle
C1525775|View 30 degree caudal angle:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525775|View 30 degree caudal angle:Find:Pt:Shoulder.bilateral:Doc:XR
C1525787|Wrist - left X-ray 2 views
C1525787|Wrist-L XR 2V
C1525787|Views 2:Find:Pt:Wrist.left:Doc:XR
C1525787|Views 2:Finding:Point in time:Wrist.left:Document:XR
C1525788|Knee-L XR AP W Stress
C1525788|Knee - left X-ray AP W manual stress
C1525788|Views AP^W manual stress:Finding:Point in time:Knee.left:Document:XR
C1525788|Views AP^W manual stress:Find:Pt:Knee.left:Doc:XR
C1525872|Unspecified body region Fluoroscopy W gastrografin via fistula
C1525872|XXX Flr W Gastrografin via Fistula
C1525872|Views^W gastrografin via fistula:Find:Pt:XXX:Doc:XR.fluor
C1525872|Views^W gastrografin via fistula:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1524141|Lymph Abd+Pelvic-Bl Flr W contr IL
C1524141|Lymphatics abdominal and Lymphatics pelvic - bilateral Fluoroscopy W contrast intra lymphatic
C1524141|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.abdominal+Lymphatics.pelvic.bilateral:Doc:XR.fluor
C1524141|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.abdominal+Lymphatics.pelvic.bilateral:Document:XR.fluor
C1525893|Orbit-Bl XRTomo
C1525893|Orbit - bilateral X-ray tomograph
C1525893|Multisection:Find:Pt:Orbit.bilateral:Doc:XR.tomo
C1525893|Multisection:Finding:Point in time:Orbit.bilateral:Document:XR.tomo
C1525807|T-spine ves MRI.Angio W contr IV
C1525807|Thoracic Spine vessels MRI angiogram W contrast IV
C1525807|Multisection^W contrast Intravenous:Finding:Point in time:Spine.thoracic vessels:Document:MRI.angio
C1525807|Multisection^W contrast IV:Find:Pt:Spine.thoracic vessels:Doc:MRI.angio
C1525950|Pelvis X-ray tomograph
C1525950|Pelvis XRTomo
C1525950|Multisection:Find:Pt:Pelvis:Doc:XR.tomo
C1525950|Multisection:Finding:Point in time:Pelvis:Document:XR.tomo
C1525974|T+L-spine XR 2V Scoli
C1525974|Views 2 scoliosis:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1525974|Spine Thoracic and Lumbar X-ray 2 views scoliosis
C1525974|Views 2 scoliosis:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1526009|Femur - right X-ray standing
C1526009|Femur-R XR stand
C1526009|Views^standing:Finding:Point in time:Femur.right:Document:XR
C1526009|Views^standing:Find:Pt:Femur.right:Doc:XR
C1526041|Hip-R XR AP+Lat
C1526041|Hip - right X-ray AP and lateral
C1526041|Views AP & lateral:Finding:Point in time:Hip.right:Document:XR
C1526041|Views AP & lateral:Find:Pt:Hip.right:Doc:XR
C1526066|Knee-R XR Lat Hyperext
C1526066|Knee - right X-ray lateral hyperextension
C1526066|View lateral hyperextension:Finding:Point in time:Knee.right:Document:XR
C1526066|View lateral hyperextension:Find:Pt:Knee.right:Doc:XR
C1526138|SC joint XR Serendipity
C1526138|Sternoclavicular Joint X-ray Serendipity
C1526138|View Serendipity:Finding:Point in time:Sternoclavicular joint:Document:XR
C1526138|View Serendipity:Find:Pt:Sternoclavicular joint:Doc:XR
C1526143|Sinuses X-ray Single view
C1526143|Sinuses XR 1V
C1526143|View 1:Finding:Point in time:Sinuses:Document:XR
C1526143|View 1:Find:Pt:Sinuses:Doc:XR
C1524279|Thumb XR AP 1V
C1524279|Thumb X-ray AP single view
C1524279|View AP:Find:Pt:Thumb:Doc:XR
C1524279|View AP:Finding:Point in time:Thumb:Document:XR
C1526180|Tibial artery Fluoroscopic angiogram W contrast IA
C1526180|Tibl a XRA W contr IA
C1526180|Views^W contrast IA:Find:Pt:Tibial artery:Doc:XR.fluor.angio
C1526180|Views^W contrast Intra-arterial:Finding:Point in time:Tibial artery:Document:XR.fluor.angio
C1526215|Carotid artery.cervical - right Fluoroscopic angiogram W contrast IA
C1526215|Carot a.cervical-R XRA W contr IA
C1526215|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.cervical.right:Document:XR.fluor.angio
C1526215|Views^W contrast IA:Find:Pt:Carotid artery.cervical.right:Doc:XR.fluor.angio
C1526229|Ribs post-R XR
C1526229|Ribs posterior - right X-ray
C1526229|Views:Finding:Point in time:Ribs.posterior.right:Document:XR
C1526229|Views:Find:Pt:Ribs.posterior.right:Doc:XR
C1525133|Humerus-R XR Transthoracic
C1525133|Humerus - right X-ray transthoracic
C1525133|View transthoracic:Find:Pt:Humerus.right:Doc:XR
C1525133|View transthoracic:Finding:Point in time:Humerus.right:Document:XR
C1526291|Multisection:Find:Pt:Talus:Doc:CT
C1526291|Deprecated Talus CT
C1526291|Multisection:Finding:Point in time:Talus:Document:Computerized Tomography
C1526334|T-spine Flr Ltd W contr IT
C1526334|Views limited^W contrast IT:Find:Pt:Spine.thoracic:Doc:XR.fluor
C1526334|Views limited^W contrast Intrathecal:Finding:Point in time:Spine.thoracic:Document:XR.fluor
C1526334|Thoracic spine Fluoroscopy limited W contrast IT
C1526342|Toe 3rd-R XR
C1526342|Toe third - right X-ray
C1526342|Views:Find:Pt:Toe.third.right:Doc:XR
C1526342|Views:Finding:Point in time:Toe.third.right:Document:XR
C1526345|Great toe-R XR
C1526345|Great toe - right X-ray
C1526345|Views:Finding:Point in time:Great toe.right:Document:XR
C1526345|Views:Find:Pt:Great toe.right:Doc:XR
C1508088|Brst-L Mam W Air
C1508088|Breast - left Mammogram W air
C1508088|Views^W air:Finding:Point in time:Breast.left:Document:Mam
C1508088|Views^W air:Find:Pt:Breast.left:Doc:Mam
C1524860|Forearm-R CT WO contr
C1524860|Forearm - right CT WO contrast
C1524860|Multisection^WO contrast:Find:Pt:Forearm.right:Doc:CT
C1524860|Multisection^WO contrast:Finding:Point in time:Forearm.right:Document:Computerized Tomography
C1524881|Acromioclavicular Joint MRI WO contrast
C1524881|AC joint MRI WO contr
C1524881|Multisection^WO contrast:Find:Pt:Acromioclavicular joint:Doc:MRI
C1524881|Multisection^WO contrast:Finding:Point in time:Acromioclavicular joint:Document:MRI
C1524883|Lower extremity joint - left MRI WO contrast
C1524883|LE.joint-L MRI WO contr
C1524883|Multisection^WO contrast:Finding:Point in time:Lower extremity.joint.left:Document:MRI
C1524883|Multisection^WO contrast:Find:Pt:Lower extremity.joint.left:Doc:MRI
C1524888|Kidney - bilateral CT WO contrast
C1524888|Multisection^WO contrast:Find:Pt:Kidney.bilateral:Doc:CT
C1524888|Multisection^WO contrast:Finding:Point in time:Kidney.bilateral:Document:Computerized Tomography
C1524888|Kdny-Bl CT WO contr
C1524891|Knee - bilateral MRI WO contrast
C1524891|Knee-Bl MRI WO contr
C1524891|Multisection^WO contrast:Find:Pt:Knee.bilateral:Doc:MRI
C1524891|Multisection^WO contrast:Finding:Point in time:Knee.bilateral:Document:MRI
C1524516|Femur CT W contr IV
C1524516|Femur CT W contrast IV
C1524516|Multisection^W contrast IV:Find:Pt:Femur:Doc:CT
C1524516|Multisection^W contrast Intravenous:Finding:Point in time:Femur:Document:Computerized Tomography
C1524518|Femur-L CT W contr IV
C1524518|Femur - left CT W contrast IV
C1524518|Multisection^W contrast IV:Find:Pt:Femur.left:Doc:CT
C1524518|Multisection^W contrast Intravenous:Finding:Point in time:Femur.left:Document:Computerized Tomography
C1524521|Thigh-R MRI W contr IV
C1524521|Thigh - right MRI W contrast IV
C1524521|Multisection^W contrast IV:Find:Pt:Thigh.right:Doc:MRI
C1524521|Multisection^W contrast Intravenous:Finding:Point in time:Thigh.right:Document:MRI
C1524524|Ft-Bl MRI W contr IV
C1524524|Foot - bilateral MRI W contrast IV
C1524524|Multisection^W contrast IV:Find:Pt:Foot.bilateral:Doc:MRI
C1524524|Multisection^W contrast Intravenous:Finding:Point in time:Foot.bilateral:Document:MRI
C1524168|Hip-Bl MRI W contr IV
C1524168|Hip - bilateral MRI W contrast IV
C1524168|Multisection^W contrast Intravenous:Finding:Point in time:Hip.bilateral:Document:MRI
C1524168|Multisection^W contrast IV:Find:Pt:Hip.bilateral:Doc:MRI
C1524149|Shoulder - bilateral MRI WO contrast
C1524149|Should-Bl MRI WO contr
C1524149|Multisection^WO contrast:Finding:Point in time:Shoulder.bilateral:Document:MRI
C1524149|Multisection^WO contrast:Find:Pt:Shoulder.bilateral:Doc:MRI
C1524151|Should-R CT WO contr
C1524151|Shoulder - right CT WO contrast
C1524151|Multisection^WO contrast:Finding:Point in time:Shoulder.right:Document:Computerized Tomography
C1524151|Multisection^WO contrast:Find:Pt:Shoulder.right:Doc:CT
C1524926|Abdomen X-ray Single view
C1524926|Abd XR 1V
C1524926|View 1:Find:Pt:Abdomen:Doc:XR
C1524926|View 1:Finding:Point in time:Abdomen:Document:XR
C1524928|Chest XR 1V
C1524928|Chest X-ray Single view
C1524928|View 1:Find:Pt:Chest:Doc:XR
C1524928|View 1:Finding:Point in time:Chest:Document:XR
C1524552|SIJ MRI W contr IV
C1524552|Sacroiliac Joint MRI W contrast IV
C1524552|Multisection^W contrast IV:Find:Pt:Sacroiliac joint:Doc:MRI
C1524552|Multisection^W contrast Intravenous:Finding:Point in time:Sacroiliac joint:Document:MRI
C1524933|Femur X-ray Single view
C1524933|Femur XR 1V
C1524933|View 1:Finding:Point in time:Femur:Document:XR
C1524933|View 1:Find:Pt:Femur:Doc:XR
C1524304|L-spine CT Bx guid
C1524304|Guidance for biopsy:Find:Pt:Spine.lumbar:Doc:CT
C1524304|Guidance for biopsy:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1524304|CT Guidance for biopsy of Lumbar spine
C1524587|Should-R CT W contr IV
C1524587|Shoulder - right CT W contrast IV
C1524587|Multisection^W contrast IV:Find:Pt:Shoulder.right:Doc:CT
C1524587|Multisection^W contrast Intravenous:Finding:Point in time:Shoulder.right:Document:Computerized Tomography
C1524604|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ankle.right:Document:Computerized Tomography
C1524604|Ankle-R CT WO+W contr IV
C1524604|Multisection^WO & W contrast IV:Find:Pt:Ankle.right:Doc:CT
C1524604|Ankle - right CT WO and W contrast IV
C1524128|Multisection^WO & W contrast IV:Find:Pt:Calcaneus.left:Doc:CT
C1524128|Multisection^WO & W contrast Intravenous:Finding:Point in time:Calcaneus.left:Document:Computerized Tomography
C1524128|Deprecated Calcaneus - left CT WO and W contrast IV
C1524128|Deprecated Heel-L CT WO+W contr IV
C1524963|Ft-L XR Obl 1V
C1524963|Foot - left X-ray oblique single view
C1524963|View oblique:Finding:Point in time:Foot.left:Document:XR
C1524963|View oblique:Find:Pt:Foot.left:Doc:XR
C1524645|Brst Mam 4V
C1524645|Breast Mammogram 4 views
C1524645|Views 4:Finding:Point in time:Breast:Document:Mam
C1524645|Views 4:Find:Pt:Breast:Doc:Mam
C1525010|Tib+Fib-Bl XR 2V
C1525010|Tibia - bilateral and Fibula - bilateral X-ray 2 views
C1525010|Views 2:Find:Pt:Tibia.bilateral+Fibula.bilateral:Doc:XR
C1525010|Views 2:Finding:Point in time:Tibia.bilateral+Fibula.bilateral:Document:XR
C1524357|Elbow XRTomo
C1524357|Elbow X-ray tomograph
C1524357|Multisection:Finding:Point in time:Elbow:Document:XR.tomo
C1524357|Multisection:Find:Pt:Elbow:Doc:XR.tomo
C1524376|UE-L CT
C1524376|Upper extremity - left CT
C1524376|Multisection:Finding:Point in time:Upper extremity.left:Document:Computerized Tomography
C1524376|Multisection:Find:Pt:Upper extremity.left:Doc:CT
C1524736|Multisection^WO & W contrast IV:Find:Pt:Forearm.right:Doc:CT
C1524736|Forearm - right CT WO and W contrast IV
C1524736|Multisection^WO & W contrast Intravenous:Finding:Point in time:Forearm.right:Document:Computerized Tomography
C1524736|Forearm-R CT WO+W contr IV
C1525045|Humerus XR AP+Lat
C1525045|Humerus X-ray AP and lateral
C1525045|Views AP & lateral:Finding:Point in time:Humerus:Document:XR
C1525045|Views AP & lateral:Find:Pt:Humerus:Doc:XR
C1525059|Ankle-Bl XR AP+Lat+Obl
C1525059|Ankle - bilateral X-ray AP and lateral and oblique
C1525059|Views AP & lateral & oblique:Finding:Point in time:Ankle.bilateral:Document:XR
C1525059|Views AP & lateral & oblique:Find:Pt:Ankle.bilateral:Doc:XR
C1525065|Finger-Bl XR AP+Lat+Obl
C1525065|Finger - bilateral X-ray AP and lateral and oblique
C1525065|Views AP & lateral & oblique:Finding:Point in time:Finger.bilateral:Document:XR
C1525065|Views AP & lateral & oblique:Find:Pt:Finger.bilateral:Doc:XR
C1524408|Hip-L XRTomo
C1524408|Hip - left X-ray tomograph
C1524408|Multisection:Finding:Point in time:Hip.left:Document:XR.tomo
C1524408|Multisection:Find:Pt:Hip.left:Doc:XR.tomo
C1524770|Nasoph MRI WO+W contr IV
C1524770|Multisection^WO & W contrast IV:Find:Pt:Nasopharynx:Doc:MRI
C1524770|Nasopharynx MRI WO and W contrast IV
C1524770|Multisection^WO & W contrast Intravenous:Finding:Point in time:Nasopharynx:Document:MRI
C1525069|Ft-L XR AP+Lat+Obl
C1525069|Foot - left X-ray AP and lateral and oblique
C1525069|Views AP & lateral & oblique:Finding:Point in time:Foot.left:Document:XR
C1525069|Views AP & lateral & oblique:Find:Pt:Foot.left:Doc:XR
C1830272|Bone DXA Bone density
C1830272|Bone density:MAric:Pt:XXX bone:Qn:XR.DXA
C1830272|Bone density:Mass Aeric:Point in time:To be specified in another part of the message bone:Quantitative:XR.DXA
C1830272|Bone DXA BDM
C1831074|Knee - right X-ray GE 4 views
C1831074|Knee-R XR GE 4V
C1831074|Views GE 4:Find:Pt:Knee.right:Doc:XR
C1831074|Views GE 4:Finding:Point in time:Knee.right:Document:XR
C1830072|Liver SPECT blood pool
C1830072|Liver SPECT BP W RNC IV
C1830072|Multisection blood pool^W radionuclide IV:Find:Pt:Liver:Doc:Radnuc.SPECT
C1830072|Multisection blood pool^W radionuclide Intravenous:Finding:Point in time:Liver:Document:Radnuc.SPECT
C1715394|BD+PDs MRI WO contr
C1715394|Biliary ducts and Pancreatic duct MRI WO contrast
C1715394|Multisection^WO contrast:Find:Pt:Biliary ducts+Pancreatic duct:Doc:MRI
C1715394|Multisection^WO contrast:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:MRI
C2718313|Multisection:Finding:Point in time:Thoracic outlet:Narrative:ULTRASOUND
C2718313|Thoracic outlet US
C2718313|TO US
C2718313|Multisection:Finding:Point in time:Thoracic outlet:Document:Ultrasound
C2718313|Multisection:Find:Pt:Thoracic outlet:Doc:US
C1715449|Elbow X-ray 2 views portable
C1715449|Elbow XR 2V port
C1715449|Views 2 portable:Find:Pt:Elbow:Doc:XR
C1715449|Views 2 portable:Finding:Point in time:Elbow:Document:XR
C1717319|LE-Bl XR stand
C1717319|Lower extremity - bilateral X-ray standing
C1717319|View^standing:Finding:Point in time:Lower extremity.bilateral:Document:XR
C1717319|View^standing:Find:Pt:Lower extremity.bilateral:Doc:XR
C1635652|Fluoroscopy Guidance for drainage of Pharynx
C1635652|Pharynx Flr Drain guid
C1635652|Guidance for drainage:Finding:Point in time:Pharynx:Document:XR.fluor
C1635652|Guidance for drainage:Find:Pt:Pharynx:Doc:XR.fluor
C1627372|Wrist-Bl XR Scaphoid 1V
C1627372|Wrist - bilateral X-ray scaphoid single view
C1627372|View scaphoid:Find:Pt:Wrist.bilateral:Doc:XR
C1627372|View scaphoid:Finding:Point in time:Wrist.bilateral:Document:XR
C1626282|Wrist - left X-ray scaphoid single view
C1626282|Wrist-L XR Scaphoid 1V
C1626282|View scaphoid:Finding:Point in time:Wrist.left:Document:XR
C1626282|View scaphoid:Find:Pt:Wrist.left:Doc:XR
C1714802|Deprecated View AP L-lateral-decubitus:Finding:Point in time:Chest:Narrative:XR
C1714802|View AP L-lateral-decubitus:Find:Pt:Chest:Nar:XR
C1714802|Deprecated Chest X-ray AP L-lateral-decubitus
C1714802|Deprecated Chest XR AP L-Lat Decub
C1714802|View AP L-lateral-decubitus:Finding:Point in time:Chest:Narrative:XR
C1714938|Views perfusion^W stress:Finding:Point in time:Heart:Narrative:Radnuc
C1714938|Views perfusion^W stress:Find:Pt:Heart:Nar:Radnuc
C1714938|Deprecated Hrt RI PF W Stress
C1714938|Deprecated Heart Scan perfusion W stress
C1715029|Heart Scan perfusion quantitative
C1715029|Hrt RI PF Qn W RNC IV
C1715029|Views perfusion quantitative^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1715029|Views perfusion quantitative^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1715116|Should-R XR Grashey & Y
C1715116|Shoulder - right X-ray Grashey and Y
C1715116|Views Grashey & Y:Find:Pt:Shoulder.right:Doc:XR
C1715116|Views Grashey & Y:Finding:Point in time:Shoulder.right:Document:XR
C1640451|Extremity X-ray Single view
C1640451|Extr XR 1V
C1640451|View 1:Finding:Point in time:Extremity:Document:XR
C1640451|View 1:Find:Pt:Extremity:Doc:XR
C1626841|Deprecated View AP:Finding:Point in time:Abdomen:Narrative:XR
C1626841|Deprecated Abd XR AP 1V
C1626841|View AP:Find:Pt:Abdomen:Nar:XR
C1626841|Deprecated Abdomen X-ray AP
C1626841|View AP:Finding:Point in time:Abdomen:Narrative:XR
C1626175|UGI Flr +AP W H2O soluble contr PO
C1626175|Gastrointestine upper Fluoroscopy and AP W water soluble contrast PO
C1626175|Views & AP^W water soluble contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1626175|Views & AP^W water soluble contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1648359|Hand - right X-ray portable
C1648359|Hand-R XR port
C1648359|Views portable:Find:Pt:Hand.right:Doc:XR
C1648359|Views portable:Finding:Point in time:Hand.right:Document:XR
C1953990|SC joints XR GE 3V
C1953990|Sternoclavicular Joints X-ray GE 3 views
C1953990|Views GE 3:Finding:Point in time:Sternoclavicular joints:Document:XR
C1953990|Views GE 3:Find:Pt:Sternoclavicular joints:Doc:XR
C1953991|Wrist - bilateral X-ray GE 3 views
C1953991|Wrist-Bl XR GE 3V
C1953991|Views GE 3:Find:Pt:Wrist.bilateral:Doc:XR
C1953991|Views GE 3:Finding:Point in time:Wrist.bilateral:Document:XR
C3173521|Breast lymphatics - left Scan W radionuclide intra lymphatic
C3173521|Brst lymphr-L RI W RNC Intra Lymph
C3173521|Views^W radionuclide intra lymphatic:Finding:Point in time:Breast lymphatics.left:Document:Radnuc
C3173521|Views^W radionuclide intra lymphatic:Find:Pt:Breast lymphatics.left:Doc:Radnuc
C3533480|US Guidance for injection of sclerosing agent of Extremity veins - left
C3533480|Extr vv-L US Sclerosing agent inj guid
C3533480|Guidance for injection of sclerosing agent:Finding:Point in time:Extremity veins.left:Document:Ultrasound
C3533480|Guidance for injection of sclerosing agent:Find:Pt:Extremity veins.left:Doc:US
C3262946|Fluoroscopy Guidance for drainage of abscess of Pleural space
C3262946|Pl space Flr Abscess drain guid
C3262946|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space:Doc:XR.fluor
C3262946|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space:Document:XR.fluor
C3262952|Fluoroscopy Guidance for needle biopsy of Thyroid
C3262952|Thyroid Flr Bx needle guid
C3262952|Guidance for biopsy.needle:Find:Pt:Thyroid:Doc:XR.fluor
C3262952|Guidance for biopsy.needle:Finding:Point in time:Thyroid:Document:XR.fluor
C3262973|Should-L XR 3V+Ax
C3262973|Shoulder - left X-ray 3 views and axillary
C3262973|Views 3 & axillary:Find:Pt:Shoulder.left:Doc:XR
C3262973|Views 3 & axillary:Finding:Point in time:Shoulder.left:Document:XR
C3262988|Breast implant - bilateral MRI WO contrast
C3262988|Brst implant-Bl MRI WO contr
C3262988|Multisection^WO contrast:Find:Pt:Breast implant.bilateral:Doc:MRI
C3262988|Multisection^WO contrast:Finding:Point in time:Breast implant.bilateral:Document:MRI
C3482443|Deprecated Spine Lumbar CT stereotactic
C3482443|Multisection stereotactic:Find:Pt:Spine.lumbar:Doc:CT
C3482443|Deprecated L-spine CT Stereo
C3482443|Multisection stereotactic:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C3263018|MRI Guidance for needle biopsy of Muscle
C3263018|Muscle MRI Bx needle guid
C3263018|Guidance for biopsy.needle:Find:Pt:Muscle:Doc:MRI
C3263018|Guidance for biopsy.needle:Finding:Point in time:Muscle:Document:MRI
C3263028|Finger-R MRI W contr IV
C3263028|Finger - right MRI W contrast IV
C3263028|Multisection^W contrast IV:Find:Pt:Finger.right:Doc:MRI
C3263028|Multisection^W contrast Intravenous:Finding:Point in time:Finger.right:Document:MRI
C3263073|Patella - right X-ray 3 views
C3263073|Patella-R XR 3V
C3263073|Views 3:Finding:Point in time:Patella.right:Document:XR
C3263073|Views 3:Find:Pt:Patella.right:Doc:XR
C3263096|Brst-R US Asp guid
C3263096|US Guidance for aspiration of Breast - right
C3263096|Guidance for aspiration:Finding:Point in time:Breast.right:Document:Ultrasound
C3263096|Guidance for aspiration:Find:Pt:Breast.right:Doc:US
C3263216|Femoral vein and Popliteal vein US
C3263216|Fem v+Polliteal a US
C3263216|Multisection:Find:Pt:Femoral vein+Popliteal vein:Doc:US
C3263216|Multisection:Finding:Point in time:Femoral vein+Popliteal vein:Document:Ultrasound
C3484378|Elbow - bilateral X-ray and obliques
C3484378|Elbow-Bl XR +Obl
C3484378|Views & obliques:Find:Pt:Elbow.bilateral:Doc:XR
C3484378|Views & obliques:Finding:Point in time:Elbow.bilateral:Document:XR
C0942168|Should-L XR
C0942168|Shoulder - left X-ray
C0942168|Views:Find:Pt:Shoulder.left:Doc:XR
C0942168|Views:Finding:Point in time:Shoulder.left:Document:XR
C0942194|Multisection^WO & W contrast IV:Find:Pt:Ankle.right:Doc:MRI
C0942194|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ankle.right:Document:MRI
C0942194|Ankle - right MRI WO and W contrast IV
C0942194|Ankle-R MRI WO+W contr IV
C0942226|Extr-Bl CT
C0942226|Extremity - bilateral CT
C0942226|Multisection:Find:Pt:Extremity.bilateral:Doc:CT
C0942226|Multisection:Finding:Point in time:Extremity.bilateral:Document:Computerized Tomography
C0942232|Extr-R CT
C0942232|Extremity - right CT
C0942232|Multisection:Find:Pt:Extremity.right:Doc:CT
C0942232|Multisection:Finding:Point in time:Extremity.right:Document:Computerized Tomography
C0882019|CT Guidance for aspiration of Lung
C0882019|Lung CT Asp guid
C0882019|Guidance for aspiration:Find:Pt:Chest>Lung:Doc:CT
C0882019|Guidance for aspiration:Finding:Point in time:Chest>Lung:Document:Computerized Tomography
C0882032|CT Guidance for biopsy of Neck
C0882032|Neck CT Bx guid
C0882032|Guidance for biopsy:Find:Pt:Neck:Doc:CT
C0882032|Guidance for biopsy:Finding:Point in time:Neck:Document:Computerized Tomography
C0882546|Peritoneovenous shunt Scan for patency W Tc-99m DTPA IT
C0882546|PV shunt RI for Pat W Tc99mDTPA IT
C0882546|Views for shunt patency^W Tc-99m DTPA IT:Find:Pt:Peritoneovenous shunt:Doc:Radnuc
C0882546|Views for shunt patency^W Tc-99m DTPA Intrathecal:Finding:Point in time:Peritoneovenous shunt:Document:Radnuc
C0882067|Multisection^W contrast Intravenous:Finding:Point in time:Petrous part of temporal bone:Document:Computerized Tomography
C0882067|Multisection^W contrast IV:Find:Pt:Petrous part of temporal bone:Doc:CT
C0882067|Petr part temp bone CT W contr IV
C0882067|Petrous part of temporal bone CT W contrast IV
C0882105|Skull X-ray 5 views
C0882105|Skull XR 5V
C0882105|Views 5:Finding:Point in time:Skull:Document:XR
C0882105|Views 5:Find:Pt:Skull:Doc:XR
C0882551|Spine XR AP+Lat
C0882551|Spine X-ray AP and lateral
C0882551|Views AP & lateral:Find:Pt:Spine:Doc:XR
C0882551|Views AP & lateral:Finding:Point in time:Spine:Document:XR
C0882132|L-spine XR AP+Lat
C0882132|Views AP & lateral:Finding:Point in time:Spine.lumbar:Document:XR
C0882132|Views AP & lateral:Find:Pt:Spine.lumbar:Doc:XR
C0882132|Lumbar spine X-ray AP and lateral
C0882176|Bladder+Urethra Flr W contr RU
C0882176|Urinary Bladder and Urethra Fluoroscopy W contrast retrograde via urethra
C0882176|Views^W contrast retrograde via urethra:Find:Pt:Urinary bladder+Urethra:Doc:XR.fluor
C0882176|Views^W contrast retrograde via urethra:Finding:Point in time:Urinary bladder+Urethra:Document:XR.fluor
C0882197|XXX CT Asp or Bx guid W contr IV
C0882197|CT Guidance for aspiration or biopsy of Unspecified body region-- W contrast IV
C0882197|Guidance for aspiration or biopsy^W contrast IV:Find:Pt:XXX:Doc:CT
C0882197|Guidance for aspiration or biopsy^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882212|XXX US No charge
C0882212|Unspecified body region US No charge
C0882212|No charge:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C0882212|No charge:Find:Pt:XXX:Doc:US
C0942135|Deprecated Views:Finding:Point in time:Femur.bilateral:Narrative:XR.DEXA
C0942135|Deprecated Femur-Bl DEXA
C0942135|Views:Find:Pt:Femur.bilateral:Nar:XR.DEXA
C0942135|Views:Finding:Point in time:Femur.bilateral:Narrative:XR.DEXA
C0942135|Deprecated Femur - bilateral DEXA Bone density
C0942140|Views:Finding:Point in time:Finger.right:Narrative:XR
C0942140|Finger - right X-ray
C0942140|Finger-R XR
C0942140|Views:Find:Pt:Finger.right:Doc:XR
C0942140|Views:Finding:Point in time:Finger.right:Document:XR
C0942141|Foot - bilateral X-ray
C0942141|Ft-Bl XR
C0942141|Views:Finding:Point in time:Foot.bilateral:Document:XR
C0942141|Views:Find:Pt:Foot.bilateral:Doc:XR
C1114681|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity vessels:Narrative:MRI.angio
C1114681|UE ves MRI.Angio W contr IV
C1114681|Upper extremity vessels MRI angiogram W contrast IV
C1114681|Multisection^W contrast IV:Find:Pt:Upper extremity vessels:Doc:MRI.angio
C1114681|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity vessels:Document:MRI.angio
C0881795|Multisection:Finding:Point in time:Abdomen:Narrative:MRI
C0881795|Abdomen MRI
C0881795|Abd MRI
C0881795|Multisection:Find:Pt:Abdomen:Doc:MRI
C0881795|Multisection:Finding:Point in time:Abdomen:Document:MRI
C0881822|Head CT Bx Str Guid W contr IV
C0881822|Guidance for stereotactic biopsy^W contrast IV:Find:Pt:Head:Doc:CT
C0881822|CT Guidance for stereotactic biopsy of Head-- W contrast IV
C0881822|Guidance for stereotactic biopsy^W contrast Intravenous:Finding:Point in time:Head:Document:Computerized Tomography
C2607990|Views AP portable:Finding:Point in time:Chest:Narrative:XR
C2607990|Chest XR AP ports
C2607990|Chest X-ray AP portable
C2607990|Views AP portable:Finding:Point in time:Chest:Document:XR
C2607990|Views AP portable:Find:Pt:Chest:Doc:XR
C0881890|Sacrum+Coccyx XR
C0881890|Sacrum and Coccyx X-ray
C0881890|Views:Finding:Point in time:Sacrum+Coccyx:Narrative:XR
C0881890|Views:Find:Pt:Sacrum+Coccyx:Doc:XR
C0881890|Views:Finding:Point in time:Sacrum+Coccyx:Document:XR
C0882532|GB XR W contr PO
C0882532|Gallbladder X-ray W contrast PO
C0882532|Views^W contrast Oral:Finding:Point in time:Gallbladder:Document:XR
C0882532|Views^W contrast PO:Find:Pt:Gallbladder:Doc:XR
C0881956|Head.SS MRI
C0881956|Head Sagittal Sinus MRI
C0881956|Multisection:Finding:Point in time:Head.sagittal sinus:Document:MRI
C0881956|Multisection:Find:Pt:Head.sagittal sinus:Doc:MRI
C0881963|Vein VD admin into cath
C0881963|Administration of vasodilator into catheter of Vein
C0881963|Administration of vasodilator into catheter:Finding:Point in time:Vein:Document
C0881963|Administration of vasodilator into catheter:Find:Pt:Vein:Doc
C0881997|Abd XR AP+Obl Prone
C0881997|Abdomen X-ray AP and oblique prone
C0881997|Views AP & oblique prone:Finding:Point in time:Abdomen:Document:XR
C0881997|Views AP & oblique prone:Find:Pt:Abdomen:Doc:XR
C0882006|Knee XR AP 1V stand
C0882006|Knee X-ray AP single view standing
C0882006|View AP^standing:Find:Pt:Knee:Doc:XR
C0882006|View AP^standing:Finding:Point in time:Knee:Document:XR
C0882010|CT Guidance for biopsy of Liver
C0882010|Liver CT Bx guid
C0882010|Guidance for biopsy:Find:Pt:Abdomen>Liver:Doc:CT
C0882010|Guidance for biopsy:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C0882014|Liver SPECT W Tc99mIV
C0882014|Liver SPECT W Tc-99m IV
C0882014|Multisection^W Tc-99m IV:Find:Pt:Liver:Doc:Radnuc.SPECT
C0882014|Multisection^W Tc-99m Intravenous:Finding:Point in time:Liver:Document:Radnuc.SPECT
C1114529|T+L-spine XR Scoli AP+Lat
C1114529|Views scoliosis AP & lateral:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1114529|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral
C1114529|Views scoliosis AP & lateral:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1114559|Ribs XR port
C1114559|Ribs X-ray portable
C1114559|Views portable:Find:Pt:Ribs:Doc:XR
C1114559|Views portable:Finding:Point in time:Ribs:Document:XR
C1114560|Shoulder X-ray Single view
C1114560|Should XR 1V
C1114560|View 1:Find:Pt:Shoulder:Doc:XR
C1114560|View 1:Finding:Point in time:Shoulder:Document:XR
C1114573|Acetabulum XR port
C1114573|Acetabulum X-ray portable
C1114573|Views portable:Finding:Point in time:Acetabulum:Document:XR
C1114573|Views portable:Find:Pt:Acetabulum:Doc:XR
C1114574|Pelvis+Hip-Bl XR
C1114574|Pelvis and Hip - bilateral X-ray
C1114574|Views:Find:Pt:Pelvis+Hip.bilateral:Doc:XR
C1114574|Views:Finding:Point in time:Pelvis+Hip.bilateral:Document:XR
C1114609|Multisection^W & WO contrast IV:Find:Pt:Aorta+Femoral artery.bilateral:Doc:CT.angio
C1114609|Deprecated Aorta+Fem a-Bl CT.Angio W+WO
C1114609|Deprecated Aorta and Femoral artery - bilateral CT angiogram W and WO contrast IV
C1114609|Multisection^W & WO contrast Intravenous:Finding:Point in time:Aorta+Femoral artery.bilateral:Document:Computerized Tomography.angio
C2608012|Views^W contrast transhepatic:Finding:Point in time:Portal vein:Narrative:XR.fluor.angio
C2608012|Portal vein Fluoroscopic angiogram W contrast transhepatic
C2608012|Portal v XRA W contr TH
C2608012|Views^W contrast transhepatic:Finding:Point in time:Portal vein:Document:XR.fluor.angio
C2608012|Views^W contrast transhepatic:Find:Pt:Portal vein:Doc:XR.fluor.angio
C1114647|Extremity arteries Fluoroscopic angiogram W contrast IA
C1114647|Extr aa XRA W contr IA
C1114647|Views^W contrast IA:Find:Pt:Extremity arteries:Doc:XR.fluor.angio
C1114647|Views^W contrast Intra-arterial:Finding:Point in time:Extremity arteries:Document:XR.fluor.angio
C1114675|Head+Neck ves DOP
C1114675|Head vessels and Neck vessels US.doppler
C1114675|Multisection:Find:Pt:Head vessels+Neck vessels:Doc:US.doppler
C1114675|Multisection:Finding:Point in time:Head vessels+Neck vessels:Document:Ultrasound.doppler
C1114447|SIJ CT
C1114447|Sacroiliac Joint CT
C1114447|Multisection:Find:Pt:Sacroiliac joint:Doc:CT
C1114447|Multisection:Finding:Point in time:Sacroiliac joint:Document:Computerized Tomography
C1114448|L-spine CT WO contr
C1114448|Multisection^WO contrast:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1114448|Multisection^WO contrast:Find:Pt:Spine.lumbar:Doc:CT
C1114448|Lumbar spine CT WO contrast
C1543762|Hrt SPECT PF W Tc99mMIBI IV
C1543762|Heart SPECT perfusion W Tc-99m Sestamibi IV
C1543762|Multisection perfusion^W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543762|Multisection perfusion^W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543763|Hrt SPECT PF W Tl-201 IV
C1543763|Heart SPECT perfusion W Tl-201 IV
C1543763|Multisection perfusion^W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543763|Multisection perfusion^W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543767|Hrt RI PF W Stress+W Tl-201 IV
C1543767|Heart Scan perfusion W stress and W Tl-201 IV
C1543767|Views perfusion^W stress & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1543767|Views perfusion^W stress & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543768|Hrt RI PF W RNC IV
C1543768|Heart Scan perfusion
C1543768|Views perfusion^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543768|Views perfusion^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C2713299|Knee-R XR +Obl
C2713299|Knee - right X-ray and oblique
C2713299|Views & oblique:Finding:Point in time:Knee.right:Document:XR
C2713299|Views & oblique:Find:Pt:Knee.right:Doc:XR
C1543474|Should-R XR AP(w IR)+West Point
C1543474|Shoulder - right X-ray AP (W internal rotation) and West Point
C1543474|Views AP (W internal rotation) & West Point:Finding:Point in time:Shoulder.right:Document:XR
C1543474|Views AP (W internal rotation) & West Point:Find:Pt:Shoulder.right:Doc:XR
C1543781|Hrt SPECT PF Rest+W Tl201 IV
C1543781|Heart SPECT perfusion at rest and W Tl-201 IV
C1543781|Multisection perfusion^at rest & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543781|Multisection perfusion^at rest & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543853|SPECT for abscess
C1543853|SPECT for Abscess W RNC IV
C1543853|Multisection for abscess^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543853|Multisection for abscess^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543871|RI for Tumor WB W Ga-67 IV
C1543871|Views for tumor whole body^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543871|Views for tumor whole body^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543871|Scan for tumor whole body W Ga-67 IV
C1543887|Adrenal RI W I-131 mIBG IV
C1543887|Adrenal gland Scan W I-131 MIBG IV
C1543887|Views^W I-131 MIBG IV:Find:Pt:Adrenal gland:Doc:Radnuc
C1543887|Views^W I-131 MIBG Intravenous:Finding:Point in time:Adrenal gland:Document:Radnuc
C1543919|Liver+Lung RI W RNC IV
C1543919|Liver and Lung Scan
C1543919|Views^W radionuclide IV:Find:Pt:Liver+Lung:Doc:Radnuc
C1543919|Views^W radionuclide Intravenous:Finding:Point in time:Liver+Lung:Document:Radnuc
C1543924|Bone RI 3 Phase single W RNC IV
C1543924|Bone Scan 3 views phase single area
C1543924|Views 3 phase single area^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543924|Views 3 phase single area ^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543499|Upper extremity artery - bilateral US.doppler
C1543499|UE a-Bl DOP
C1543499|Multisection:Find:Pt:Upper extremity artery.bilateral:Doc:US.doppler
C1543499|Multisection:Finding:Point in time:Upper extremity artery.bilateral:Document:Ultrasound.doppler
C1543529|Multisection:Finding:Point in time:To be specified in another part of the message tendon:Narrative:ULTRASOUND
C1543529|Tendon US
C1543529|Multisection:Finding:Point in time:To be specified in another part of the message tendon:Document:Ultrasound
C1543529|Multisection:Find:Pt:XXX tendon:Doc:US
C1543191|Chest XR AP+Lat+Lordotic
C1543191|Chest X-ray AP and lateral and lordotic
C1543191|Views AP & lateral & lordotic:Finding:Point in time:Chest:Document:XR
C1543191|Views AP & lateral & lordotic:Find:Pt:Chest:Doc:XR
C1543598|Artery DOP
C1543598|Artery US.doppler
C1543598|Multisection:Finding:Point in time:To be specified in another part of the message artery:Document:Ultrasound.doppler
C1543598|Multisection:Find:Pt:XXX artery:Doc:US.doppler
C1543691|Meckels divertic RI W RNC IV
C1543691|Meckels diverticulum Scan
C1543691|Views^W radionuclide IV:Find:Pt:Meckels diverticulum:Doc:Radnuc
C1543691|Views^W radionuclide Intravenous:Finding:Point in time:Meckels diverticulum:Document:Radnuc
C1543692|Brain RI W Tc99mHMPAO IV
C1543692|Brain Scan W Tc-99m HMPAO IV
C1543692|Views^W Tc-99m HMPAO Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1543692|Views^W Tc-99m HMPAO IV:Find:Pt:Brain:Doc:Radnuc
C1524255|Shoulder - right X-ray Velpeau axillary
C1524255|Should-R XR Velpeau Ax
C1524255|View Velpeau axillary:Finding:Point in time:Shoulder.right:Document:XR
C1524255|View Velpeau axillary:Find:Pt:Shoulder.right:Doc:XR
C1526785|UE-L MRI W contr IV
C1526785|Upper extremity - left MRI W contrast IV
C1526785|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.left:Document:MRI
C1526785|Multisection^W contrast IV:Find:Pt:Upper extremity.left:Doc:MRI
C1526790|Shoulder - left MRI WO contrast
C1526790|Should-L MRI WO contr
C1526790|Multisection^WO contrast:Finding:Point in time:Shoulder.left:Document:MRI
C1526790|Multisection^WO contrast:Find:Pt:Shoulder.left:Doc:MRI
C1524842|UE-L CT WO contr
C1524842|Upper extremity - left CT WO contrast
C1524842|Multisection^WO contrast:Finding:Point in time:Upper extremity.left:Document:Computerized Tomography
C1524842|Multisection^WO contrast:Find:Pt:Upper extremity.left:Doc:CT
C1525116|IVC+LE vv MRI.Angio
C1525116|Vena cava.inferior and Lower extremity veins MRI angiogram
C1525116|Multisection:Finding:Point in time:Vena cava.inferior+Lower extremity veins:Document:MRI.angio
C1525116|Multisection:Find:Pt:Vena cava.inferior+Lower extremity veins:Doc:MRI.angio
C1525119|Carot ves MRI.Angio
C1525119|Carotid vessel MRI angiogram
C1525119|Multisection:Find:Pt:Carotid vessel:Doc:MRI.angio
C1525119|Multisection:Finding:Point in time:Carotid vessel:Document:MRI.angio
C1525171|Lower extremity vessels - left MRI angiogram
C1525171|LE ves-L MRI.Angio
C1525171|Multisection:Finding:Point in time:Lower extremity vessels.left:Document:MRI.angio
C1525171|Multisection:Find:Pt:Lower extremity vessels.left:Doc:MRI.angio
C1525181|Should ves MRI.Angio
C1525181|Shoulder vessels MRI angiogram
C1525181|Multisection:Find:Pt:Shoulder vessels:Doc:MRI.angio
C1525181|Multisection:Finding:Point in time:Shoulder vessels:Document:MRI.angio
C1525304|Wrist-L XR Lat W Flx
C1525304|Wrist - left X-ray lateral W flexion
C1525304|View lateral^W flexion:Find:Pt:Wrist.left:Doc:XR
C1525304|View lateral^W flexion:Finding:Point in time:Wrist.left:Document:XR
C1525306|Should-L XR Garth
C1525306|Shoulder - left X-ray Garth
C1525306|View Garth:Find:Pt:Shoulder.left:Doc:XR
C1525306|View Garth:Finding:Point in time:Shoulder.left:Document:XR
C1525209|Vessel CT angiogram W contrast IV
C1525209|Multisection^W contrast Intravenous:Finding:Point in time:Vessel:Document:Computerized Tomography.angio
C1525209|Multisection^W contrast IV:Find:Pt:Vessel:Doc:CT.angio
C1525209|Vesl CT.Angio W contr IV
C1525219|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ovary:Document:MRI
C1525219|Ovary MRI WO+W contr IV
C1525219|Ovary MRI WO and W contrast IV
C1525219|Multisection^WO & W contrast IV:Find:Pt:Ovary:Doc:MRI
C1525342|Chest XR R-Obl
C1525342|Chest X-ray right oblique
C1525342|View R-oblique:Finding:Point in time:Chest:Document:XR
C1525342|View R-oblique:Find:Pt:Chest:Doc:XR
C1525348|Skull XR SMV
C1525348|Skull X-ray submentovertex
C1525348|View submentovertex:Finding:Point in time:Skull:Document:XR
C1525348|View submentovertex:Find:Pt:Skull:Doc:XR
C1524228|Breast - left Mammogram XCCL
C1524228|Brst-L Mam XCCL
C1524228|View XCCL:Finding:Point in time:Breast.left:Document:Mam
C1524228|View XCCL:Find:Pt:Breast.left:Doc:Mam
C1525527|Should-Bl XR Ax+Y
C1525527|Shoulder - bilateral X-ray axillary and Y
C1525527|Views axillary & Y:Find:Pt:Shoulder.bilateral:Doc:XR
C1525527|Views axillary & Y:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525616|BD+PDs MRI
C1525616|Biliary ducts and Pancreatic duct MRI
C1525616|Multisection:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:MRI
C1525616|Multisection:Find:Pt:Biliary ducts+Pancreatic duct:Doc:MRI
C1525691|L-spine+Sacrum+SIJ+Coccyx XR
C1525691|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray
C1525691|Views:Finding:Point in time:Spine.lumbar+Sacrum+Sacroiliac joint+Coccyx:Document:XR
C1525691|Views:Find:Pt:Spine.lumbar+Sacrum+Sacroiliac joint+Coccyx:Doc:XR
C1525730|Subclavian a-Bl XRA W contr IA
C1525730|Subclavian artery - bilateral Fluoroscopic angiogram W contrast IA
C1525730|Views^W contrast IA:Find:Pt:Subclavian artery.bilateral:Doc:XR.fluor.angio
C1525730|Views^W contrast Intra-arterial:Finding:Point in time:Subclavian artery.bilateral:Document:XR.fluor.angio
C1525773|Wrist-R MRI WO contr
C1525773|Wrist - right MRI WO contrast
C1525773|Multisection^WO contrast:Find:Pt:Wrist.right:Doc:MRI
C1525773|Multisection^WO contrast:Finding:Point in time:Wrist.right:Document:MRI
C1525858|Knee - left X-ray W manual stress
C1525858|Knee-L XR W Stress
C1525858|Views^W manual stress:Finding:Point in time:Knee.left:Document:XR
C1525858|Views^W manual stress:Find:Pt:Knee.left:Doc:XR
C1525824|Finger second - bilateral X-ray
C1525824|Finger.2nd-Bl XR
C1525824|Views:Finding:Point in time:Finger.second.bilateral:Document:XR
C1525824|Views:Find:Pt:Finger.second.bilateral:Doc:XR
C1525954|Abdomen X-ray
C1525954|Abd XR
C1525954|Views:Finding:Point in time:Abdomen:Narrative:XR
C1525954|Views:Find:Pt:Abdomen:Doc:XR
C1525954|Views:Finding:Point in time:Abdomen:Document:XR
C1525996|Clavicle-R XR AP+Serendipity
C1525996|Clavicle - right X-ray AP and Serendipity
C1525996|Views AP & Serendipity:Find:Pt:Clavicle.right:Doc:XR
C1525996|Views AP & Serendipity:Finding:Point in time:Clavicle.right:Document:XR
C1526121|Tib+Fib-R XR AP+Lat
C1526121|Tibia - right and Fibula - right X-ray AP and lateral
C1526121|Views AP & lateral:Finding:Point in time:Tibia.right+Fibula.right:Document:XR
C1526121|Views AP & lateral:Find:Pt:Tibia.right+Fibula.right:Doc:XR
C1526082|LE-R XRTomo
C1526082|Lower extremity - right X-ray tomograph
C1526082|Multisection:Find:Pt:Lower extremity.right:Doc:XR.tomo
C1526082|Multisection:Finding:Point in time:Lower extremity.right:Document:XR.tomo
C1526090|Views^W contrast IS:Find:Pt:Sacroiliac joint.right:Doc:XR.fluor
C1526090|Sacroiliac joint - right Fluoroscopy W contrast IS
C1526090|SIJ-R Flr W contr IS
C1526090|Views^W contrast Intrasynovial:Finding:Point in time:Sacroiliac joint.right:Document:XR.fluor
C1524273|Sternum XR PA+Lat+Obl
C1524273|Sternum X-ray PA and lateral and oblique
C1524273|Views PA & lateral & oblique:Finding:Point in time:Sternum:Document:XR
C1524273|Views PA & lateral & oblique:Find:Pt:Sternum:Doc:XR
C1526184|T-spine XR 1V
C1526184|View 1:Finding:Point in time:Spine.thoracic:Document:XR
C1526184|View 1:Find:Pt:Spine.thoracic:Doc:XR
C1526184|Thoracic spine X-ray Single view
C1526250|Elbow XR Radial Head Capitellar
C1526250|Elbow X-ray radial head capitellar
C1526250|View radial head capitellar:Find:Pt:Elbow:Doc:XR
C1526250|View radial head capitellar:Finding:Point in time:Elbow:Document:XR
C1525135|T-spine XR AP+Lat+Swimmers
C1525135|Views AP & lateral & Swimmers:Finding:Point in time:Spine.thoracic:Document:XR
C1525135|Views AP & lateral & Swimmers:Find:Pt:Spine.thoracic:Doc:XR
C1525135|Thoracic spine X-ray AP and lateral and Swimmers
C1526261|Gallbladder US limited
C1526261|GB US Ltd
C1526261|Multisection limited:Find:Pt:Gallbladder:Doc:US
C1526261|Multisection limited:Finding:Point in time:Gallbladder:Document:Ultrasound
C1526263|GB US W CCK
C1526263|Gallbladder US W cholecystokinin
C1526263|Multisection^W cholecystokinin:Find:Pt:Gallbladder:Doc:US
C1526263|Multisection^W cholecystokinin:Finding:Point in time:Gallbladder:Document:Ultrasound
C1526271|US Guidance for needle biopsy of Spleen
C1526271|Spleen US Bx needle guid
C1526271|Guidance for biopsy.needle:Find:Pt:Spleen:Doc:US
C1526271|Guidance for biopsy.needle:Finding:Point in time:Spleen:Document:Ultrasound
C1526296|Hip - left X-ray lateral during surgery
C1526296|Hip-L XR Lat in Surg
C1526296|View lateral^during surgery:Find:Pt:Hip.left:Doc:XR
C1526296|View lateral^during surgery:Finding:Point in time:Hip.left:Document:XR
C1526335|T+L-spine XR 1V
C1526335|Spine Thoracic and Lumbar X-ray Single view
C1526335|View 1:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1526335|View 1:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1526337|T+L-spine XR stand
C1526337|Spine Thoracic and Lumbar X-ray standing
C1526337|Views^standing:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1526337|Views^standing:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1526307|Views magnification & spot^compression:Find:Pt:Breast.left:Nar:Mam
C1526307|Views magnification & spot^compression:Finding:Point in time:Breast.left:Narrative:Mam
C1526307|Deprecated Brst-L Mam Mag+Spot Compressi
C1526307|Deprecated Breast - left Mammogram magnification & spot compression
C1524527|Ft-R CT W contr IV
C1524527|Foot - right CT W contrast IV
C1524527|Multisection^W contrast IV:Find:Pt:Foot.right:Doc:CT
C1524527|Multisection^W contrast Intravenous:Finding:Point in time:Foot.right:Document:Computerized Tomography
C1524532|Forearm-L MRI W contr IV
C1524532|Forearm - left MRI W contrast IV
C1524532|Multisection^W contrast IV:Find:Pt:Forearm.left:Doc:MRI
C1524532|Multisection^W contrast Intravenous:Finding:Point in time:Forearm.left:Document:MRI
C1524165|Hip MRI W contr IV
C1524165|Hip MRI W contrast IV
C1524165|Multisection^W contrast IV:Find:Pt:Hip:Doc:MRI
C1524165|Multisection^W contrast Intravenous:Finding:Point in time:Hip:Document:MRI
C1524152|Shoulder - right MRI WO contrast
C1524152|Should-R MRI WO contr
C1524152|Multisection^WO contrast:Finding:Point in time:Shoulder.right:Document:MRI
C1524152|Multisection^WO contrast:Find:Pt:Shoulder.right:Doc:MRI
C1524555|Kidney-R MRI W contr IV
C1524555|Kidney - right MRI W contrast IV
C1524555|Multisection^W contrast IV:Find:Pt:Kidney.right:Doc:MRI
C1524555|Multisection^W contrast Intravenous:Finding:Point in time:Kidney.right:Document:MRI
C1524561|Knee-R CT W contr IV
C1524561|Knee - right CT W contrast IV
C1524561|Multisection^W contrast Intravenous:Finding:Point in time:Knee.right:Document:Computerized Tomography
C1524561|Multisection^W contrast IV:Find:Pt:Knee.right:Doc:CT
C1524291|Head CT Bx guid
C1524291|CT Guidance for biopsy of Head
C1524291|Guidance for biopsy:Find:Pt:Head:Doc:CT
C1524291|Guidance for biopsy:Finding:Point in time:Head:Document:Computerized Tomography
C1524303|C-spine CT Bx guid
C1524303|Guidance for biopsy:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C1524303|Guidance for biopsy:Find:Pt:Spine.cervical:Doc:CT
C1524303|CT Guidance for biopsy of Cervical spine
C1524620|Ankle X-ray 3 views
C1524620|Ankle XR 3V
C1524620|Views 3:Finding:Point in time:Ankle:Document:XR
C1524620|Views 3:Find:Pt:Ankle:Doc:XR
C1524960|Finger second X-ray oblique single view
C1524960|Finger.2nd XR Obl 1V
C1524960|View oblique:Find:Pt:Finger.second:Doc:XR
C1524960|View oblique:Finding:Point in time:Finger.second:Document:XR
C1524961|Finger.3rd XR Obl 1V
C1524961|Finger third X-ray oblique single view
C1524961|View oblique:Find:Pt:Finger.third:Doc:XR
C1524961|View oblique:Finding:Point in time:Finger.third:Document:XR
C1524318|CT Guidance for drainage of Liver
C1524318|Liver CT Drain guid
C1524318|Guidance for drainage:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1524318|Guidance for drainage:Find:Pt:Abdomen>Liver:Doc:CT
C1524629|Finger X-ray 3 views
C1524629|Finger XR 3V
C1524629|Views 3:Find:Pt:Finger:Doc:XR
C1524629|Views 3:Finding:Point in time:Finger:Document:XR
C1524647|Chest Fluoroscopy 4 views
C1524647|Chest Flr 4V
C1524647|Views 4:Finding:Point in time:Chest:Document:XR.fluor
C1524647|Views 4:Find:Pt:Chest:Doc:XR.fluor
C1524381|Femur - left CT
C1524381|Femur-L CT
C1524381|Multisection:Finding:Point in time:Femur.left:Document:Computerized Tomography
C1524381|Multisection:Find:Pt:Femur.left:Doc:CT
C1525025|Deprecated Calcaneus - bilateral X-ray AP and lateral
C1525025|Views AP & lateral:Finding:Point in time:Calcaneus.bilateral:Document:XR
C1525025|Deprecated Heel-Bl XR AP+Lat
C1525025|Views AP & lateral:Find:Pt:Calcaneus.bilateral:Doc:XR
C1525054|Scapula-L XR AP+Lat
C1525054|Scapula - left X-ray AP and lateral
C1525054|Views AP & lateral:Finding:Point in time:Scapula.left:Document:XR
C1525054|Views AP & lateral:Find:Pt:Scapula.left:Doc:XR
C1524420|Sacroiliac Joint MRI
C1524420|SIJ MRI
C1524420|Multisection:Finding:Point in time:Sacroiliac joint:Document:MRI
C1524420|Multisection:Find:Pt:Sacroiliac joint:Doc:MRI
C1527044|Knee CT
C1527044|Multisection:Find:Pt:Knee:Doc:CT
C1527044|Multisection:Finding:Point in time:Knee:Document:Computerized Tomography
C1525083|Hand XR PA+Lat+Obl
C1525083|Hand X-ray PA and lateral and oblique
C1525083|Views PA & lateral & oblique:Find:Pt:Hand:Doc:XR
C1525083|Views PA & lateral & oblique:Finding:Point in time:Hand:Document:XR
C1525088|AV shunt Fluoroscopic angiogram Angioplasty W contrast
C1525088|AV shunt XRA Angpsty W contr
C1525088|Angioplasty^W contrast:Find:Pt:AV shunt:Doc:XR.fluor.angio
C1525088|Angioplasty^W contrast:Finding:Point in time:AV shunt:Document:XR.fluor.angio
C1525090|Extremity vessel Fluoroscopic angiogram Angioplasty W contrast
C1525090|Extr ves XRA Angpsty W contr
C1525090|Angioplasty^W contrast:Find:Pt:Extremity vessel:Doc:XR.fluor.angio
C1525090|Angioplasty^W contrast:Finding:Point in time:Extremity vessel:Document:XR.fluor.angio
C1830197|Brst Mam Bx CN Str Guid
C1830197|Guidance for stereotactic biopsy.core needle:Finding:Point in time:Breast:Document:Mam
C1830197|Mammogram Guidance for stereotactic core needle biopsy of Breast
C1830197|Guidance for stereotactic biopsy.core needle:Find:Pt:Breast:Doc:Mam
C1830084|Pelvis US Bx needle guid
C1830084|US Guidance for needle biopsy of Pelvis
C1830084|Guidance for biopsy.needle:Find:Pt:Pelvis:Doc:US
C1830084|Guidance for biopsy.needle:Finding:Point in time:Pelvis:Document:Ultrasound
C1831068|Hand - left X-ray GE 3 views
C1831068|Hand-L XR GE 3V
C1831068|Views GE 3:Finding:Point in time:Hand.left:Document:XR
C1831068|Views GE 3:Find:Pt:Hand.left:Doc:XR
C1717312|Adrenal MRI W contr IV
C1717312|Adrenal gland MRI W contrast IV
C1717312|Multisection^W contrast IV:Find:Pt:Adrenal gland:Doc:MRI
C1717312|Multisection^W contrast Intravenous:Finding:Point in time:Adrenal gland:Document:MRI
C1717318|Spine X-ray GE 4 views W right bending and W left bending
C1717318|Spine XR GE 4V W R+L-bending
C1717318|Views GE 4^W R-Bending & W L-Bending:Find:Pt:Spine:Doc:XR
C1717318|Views GE 4^W R-Bending & W L-Bending:Finding:Point in time:Spine:Document:XR
C1643598|Ankle-L XR port
C1643598|Ankle - left X-ray portable
C1643598|Views portable:Find:Pt:Ankle.left:Doc:XR
C1643598|Views portable:Finding:Point in time:Ankle.left:Document:XR
C1714805|Views:Finding:Point in time:To be specified in another part of the message:Narrative:XR
C1714805|XXX XR
C1714805|Unspecified body region X-ray
C1714805|Views:Find:Pt:XXX:Doc:XR
C1714805|Views:Finding:Point in time:To be specified in another part of the message:Document:XR
C1714813|BD+PDs Flr Endo guid 45M p contr retro
C1714813|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 45 minutes post contrast retrograde
C1714813|Guidance for endoscopy^45M post contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1714813|Guidance for endoscopy^45M post contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1706622|Finger fourth - left X-ray GE 3 views
C1706622|Finger.4th-L XR GE 3V
C1706622|Finger fourth - left Narrative X-ray GE 3 views
C1706622|Views GE 3:Finding:Point in time:Finger.fourth.left:Document:XR
C1706622|Views GE 3:Find:Pt:Finger.fourth.left:Doc:XR
C1714918|Views survey limited:Finding:Point in time:To be specified in another part of the message bones:Narrative:XR
C1714918|Bones X-ray survey limited
C1714918|Bones XR Survey Ltd
C1714918|Views survey limited:Finding:Point in time:Bones:Document:XR
C1714918|Views survey limited:Find:Pt:Bones:Doc:XR
C1714927|Multisection^WO & W contrast IV:Find:Pt:Breast.unilateral:Doc:MRI
C1714927|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast.unilateral:Document:MRI
C1714927|Brst-UL MRI WO+W contr IV
C1714927|Breast - unilateral MRI WO and W contrast IV
C1706623|Deprecated Finger.4th-L XR GE 3V
C1706623|Deprecated Finger fourth Left X-ray GE 3 views
C1706623|Views GE 3:Find:Pt:Finger.fourth.left:Nar:XR
C1706623|Views GE 3:Finding:Point in time:Finger.fourth.left:Narrative:XR
C1706625|Deprecated Finger.4th-R XR GE 3V
C1706625|Views GE 3:Find:Pt:Finger.fourth.right:Nar:XR
C1706625|Deprecated Finger fourth Right X-ray GE 3 views
C1706625|Views GE 3:Finding:Point in time:Finger.fourth.right:Narrative:XR
C1714949|Views^W gastrografin PO & W barium contrast PR:Find:Pt:Colon:Nar:XR.fluor
C1714949|Views^W gastrografin Oral & W barium contrast Rectal:Finding:Point in time:Colon:Narrative:XR.fluor
C1714949|Deprecated Colon Fluoroscopy W gastrografin PO & W barium contrast PR
C1714949|Deprecated Colon Flr W Gastrografin PO+B
C1635016|US Guidance for biopsy of Breast - right
C1635016|Brst-R US Bx guid
C1635016|Guidance for biopsy:Find:Pt:Breast.right:Doc:US
C1635016|Guidance for biopsy:Finding:Point in time:Breast.right:Document:Ultrasound
C1638467|Gastrointestine upper Fluoroscopy W contrast PO
C1638467|UGI Flr W contr PO
C1638467|Views^W contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1638467|Views^W contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1634493|Pelvis+Hip-R XR 2V
C1634493|Pelvis and Hip - right X-ray 2 views
C1634493|Views 2:Find:Pt:Pelvis+Hip.right:Doc:XR
C1634493|Views 2:Finding:Point in time:Pelvis+Hip.right:Document:XR
C1644644|Abdomen X-ray during surgery
C1644644|Abd XR in Surg
C1644644|View^during surgery:Finding:Point in time:Abdomen:Document:XR
C1644644|View^during surgery:Find:Pt:Abdomen:Doc:XR
C1623598|Appendix US Abscess drain guid
C1623598|US Guidance for drainage of abscess of Appendix
C1623598|Guidance for drainage of abscess:Find:Pt:Appendix:Doc:US
C1623598|Guidance for drainage of abscess:Finding:Point in time:Appendix:Document:Ultrasound
C1977324|Hrt SPECT PF R+S+W Tl201+Tc99mMIBI IV
C1977324|Heart SPECT perfusion at rest and W stress and W Tl-201 IV and W Tc-99m Sestamibi IV
C1977324|Multisection perfusion^at rest & W stress & W Tl-201 IV & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1977324|Multisection perfusion^at rest & W stress & W Tl-201 Intravenous & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1954373|View 1:Find:Pt:Pelvis:Nar:XR (deprecated)
C1954373|View 1:Find:Pt:Pelvis:Nar:XR
C1954373|Deprecated Pelvis X-ray View
C1954373|Deprecated Pelvis XR 1V
C1954373|View 1:Finding:Point in time:Pelvis:Narrative:XR
C1953989|Elbow - bilateral X-ray GE 3 views
C1953989|Elbow-Bl XR GE 3V
C1953989|Views GE 3:Find:Pt:Elbow.bilateral:Doc:XR
C1953989|Views GE 3:Finding:Point in time:Elbow.bilateral:Document:XR
C3174365|Fluoroscopic angiogram Guidance for placement of stent in Artery - right
C3174365|Artery.-R XRA Stent plac guid
C3174365|Guidance for placement of stent:Finding:Point in time:Artery.right:Document:XR.fluor.angio
C3174365|Guidance for placement of stent:Find:Pt:Artery.right:Doc:XR.fluor.angio
C3533574|Axilla - right US
C3533574|Multisection:Find:Pt:Axilla.right:Doc:US
C3533574|Axilla-R US
C3533574|Multisection:Finding:Point in time:Axilla.right:Document:Ultrasound
C3533572|US Guidance for injection of Joint
C3533572|Joint US Inj guid
C3533572|Guidance for injection:Find:Pt:Joint:Doc:US
C3533572|Guidance for injection:Finding:Point in time:Joint:Document:Ultrasound
C3533569|Guidance for ambulatory phlebectomy:Finding:Point in time:Extremity vein.left:Document:Ultrasound
C3533569|Extr v-L US Amb phleb guid
C3533569|US Guidance for ambulatory phlebectomy of Extremity vein - left
C3533569|Guidance for ambulatory phlebectomy:Find:Pt:Extremity vein.left:Doc:US
C3262953|Hand XR AP+Lat
C3262953|Hand X-ray AP and lateral
C3262953|Views AP & lateral:Find:Pt:Hand:Doc:XR
C3262953|Views AP & lateral:Finding:Point in time:Hand:Document:XR
C3262965|Knee-L XR 4V+Tunnel
C3262965|Knee - left X-ray 4 views and tunnel
C3262965|Views 4 & tunnel:Finding:Point in time:Knee.left:Document:XR
C3262965|Views 4 & tunnel:Find:Pt:Knee.left:Doc:XR
C3262993|Femur - bilateral MRI WO contrast
C3262993|Femur-Bl MRI WO contr
C3262993|Multisection^WO contrast:Finding:Point in time:Femur.bilateral:Document:MRI
C3262993|Multisection^WO contrast:Find:Pt:Femur.bilateral:Doc:MRI
C3263041|Prostate Flr Bx needle guid
C3263041|Fluoroscopy Guidance for needle biopsy of Prostate
C3263041|Guidance for biopsy.needle:Find:Pt:Prostate:Doc:XR.fluor
C3263041|Guidance for biopsy.needle:Finding:Point in time:Prostate:Document:XR.fluor
C3261712|Adrenal gland US
C3261712|Adrenal US
C3261712|Multisection:Finding:Point in time:Adrenal gland:Document:Ultrasound
C3261712|Multisection:Find:Pt:Adrenal gland:Doc:US
C3484382|Extr vv-Bl DOP
C3484382|Extremity veins - bilateral US.doppler
C3484382|Multisection:Find:Pt:Extremity veins.bilateral:Doc:US.doppler
C3484382|Multisection:Finding:Point in time:Extremity veins.bilateral:Document:Ultrasound.doppler
C3262882|Hip - bilateral X-ray 2 views
C3262882|Hip-Bl XR 2V
C3262882|Views 2:Finding:Point in time:Hip.bilateral:Document:XR
C3262882|Views 2:Find:Pt:Hip.bilateral:Doc:XR
C3262892|Patella - bilateral X-ray Sunrise
C3262892|Patella-Bl XR Sunrise
C3262892|View Sunrise:Finding:Point in time:Patella.bilateral:Document:XR
C3262892|View Sunrise:Find:Pt:Patella.bilateral:Doc:XR
C3262912|Knee - bilateral CT WO contrast
C3262912|Knee-Bl CT WO contr
C3262912|Multisection^WO contrast:Find:Pt:Knee.bilateral:Doc:CT
C3262912|Multisection^WO contrast:Finding:Point in time:Knee.bilateral:Document:Computerized Tomography
C0942158|Views:Find:Pt:Radius+Ulna.left:Nar:XR.DEXA
C0942158|Deprecated DEXA
C0942158|Views:Finding:Point in time:Radius+Ulna.left:Narrative:XR.DEXA
C0942158|Deprecated Radius & Ulna left DEXA Bone density
C0942162|Ribs - left X-ray
C0942162|Ribs-L XR
C0942162|Views:Finding:Point in time:Ribs.left:Document:XR
C0942162|Views:Find:Pt:Ribs.left:Doc:XR
C0942199|Elbow-R MRI WO+W contr IV
C0942199|Multisection^WO & W contrast Intravenous:Finding:Point in time:Elbow.right:Document:MRI
C0942199|Multisection^WO & W contrast IV:Find:Pt:Elbow.right:Doc:MRI
C0942199|Elbow - right MRI WO and W contrast IV
C0942218|Brst-Bl US
C0942218|Breast - bilateral US
C0942218|Multisection:Find:Pt:Breast.bilateral:Doc:US
C0942218|Multisection:Finding:Point in time:Breast.bilateral:Document:Ultrasound
C0942243|Forearm-L MRI
C0942243|Forearm - left MRI
C0942243|Multisection:Find:Pt:Forearm.left:Doc:MRI
C0942243|Multisection:Finding:Point in time:Forearm.left:Document:MRI
C0942306|CT Guidance for injection of Sacroiliac joint - bilateral
C0942306|SIJ-Bl CT Inj guid
C0942306|Guidance for injection:Finding:Point in time:Sacroiliac joint.bilateral:Document:Computerized Tomography
C0942306|Guidance for injection:Find:Pt:Sacroiliac joint.bilateral:Doc:CT
C0942317|US Guidance for drainage of Kidney - right
C0942317|Kidney-R US Drain guid
C0942317|Guidance for drainage:Finding:Point in time:Kidney.right:Document:Ultrasound
C0942317|Guidance for drainage:Find:Pt:Kidney.right:Doc:US
C0945338|Cent v-R XRA CC change guid W contr IV
C0945338|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - right-- W contrast IV
C0945338|Guidance for change of central catheter^W contrast Intravenous:Finding:Point in time:Central vein.right:Document:XR.fluor.angio
C0945338|Guidance for change of central catheter^W contrast IV:Find:Pt:Central vein.right:Doc:XR.fluor.angio
C0942345|Knee-L XR AP+Lat stand
C0942345|Knee - left X-ray AP and lateral standing
C0942345|Views AP & lateral^standing:Find:Pt:Knee.left:Doc:XR
C0942345|Views AP & lateral^standing:Finding:Point in time:Knee.left:Document:XR
C0945347|Humerus-R XR 2V
C0945347|Humerus - right X-ray 2 views
C0945347|Views 2:Finding:Point in time:Humerus.right:Document:XR
C0945347|Views 2:Find:Pt:Humerus.right:Doc:XR
C0882047|Orbit - bilateral X-ray
C0882047|Orbit-Bl XR
C0882047|Views:Finding:Point in time:Orbit.bilateral:Document:XR
C0882047|Views:Find:Pt:Orbit.bilateral:Doc:XR
C0882068|Pituitary+ST MRI WO+W contr IV
C0882068|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pituitary+Sella turcica:Document:MRI
C0882068|Multisection^WO & W contrast IV:Find:Pt:Pituitary+Sella turcica:Doc:MRI
C0882068|Pituitary and Sella turcica MRI WO and W contrast IV
C0882072|Prostate US
C0882072|Multisection:Find:Pt:Prostate:Doc:US
C0882072|Multisection:Finding:Point in time:Prostate:Document:Ultrasound
C0882074|Pulmonary artery Fluoroscopic angiogram Embolectomy W contrast IA
C0882074|PA XRA Embolectomy W contr IA
C0882074|Embolectomy^W contrast Intra-arterial:Finding:Point in time:Pulmonary artery:Document:XR.fluor.angio
C0882074|Embolectomy^W contrast IA:Find:Pt:Pulmonary artery:Doc:XR.fluor.angio
C0882125|C-spine.odontoidaxis XR AP 1V
C0882125|Spine Cervical Odontoid and Cervical axis X-ray AP single view
C0882125|View AP:Find:Pt:Spine.cervical.odontoid+Spine.cervical.axis:Doc:XR
C0882125|View AP:Finding:Point in time:Spine.cervical.odontoid+Spine.cervical.axis:Document:XR
C0882139|T-spine CT
C0882139|Multisection:Find:Pt:Spine.thoracic:Doc:CT
C0882139|Multisection:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C0882139|Thoracic spine CT
C0882151|Splenic v+Portal v XRA W contr IA
C0882151|Splenic vein and Portal vein Fluoroscopic angiogram W contrast IA
C0882151|Views^W contrast Intra-arterial:Finding:Point in time:Splenic vein+Portal vein:Document:XR.fluor.angio
C0882151|Views^W contrast IA:Find:Pt:Splenic vein+Portal vein:Doc:XR.fluor.angio
C0882171|Two vessels Fluoroscopic angiogram W contrast
C0882171|2 vess XRA W contr
C0882171|Views^W contrast:Finding:Point in time:Two vessels:Document:XR.fluor.angio
C0882171|Views^W contrast:Find:Pt:Two vessels:Doc:XR.fluor.angio
C0882179|Vein XRA W contr IV
C0882179|Vein Fluoroscopic angiogram W contrast IV
C0882179|Views^W contrast IV:Find:Pt:Vein:Doc:XR.fluor.angio
C0882179|Views^W contrast Intravenous:Finding:Point in time:Vein:Document:XR.fluor.angio
C0882202|Unspecified body region CT W anesthesia
C0882202|XXX CT W anesthesia
C0882202|Multisection^W anesthesia:Find:Pt:XXX:Doc:CT
C0882202|Multisection^W anesthesia:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882204|Deprecated XXX CT.3D Sagittal & coronal
C0882204|Views multiple sagittal & coronal:Find:Pt:XXX:Nar:CT.3D
C0882204|Deprecated Unspecified body region CT 3D multiple sagittal & coronal
C0882204|Views multiple sagittal & coronal:Finding:Point in time:To be specified in another part of the message:Narrative:Computerized Tomography.3D
C0882228|Renal ves XRA Angpsty W contr IA
C0882228|Renal vessel Fluoroscopic angiogram Angioplasty W contrast IA
C0882228|Angioplasty^W contrast IA:Find:Pt:Renal vessel:Doc:XR.fluor.angio
C0882228|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Renal vessel:Document:XR.fluor.angio
C0942101|Carotid artery - left Fluoroscopic angiogram W contrast IA
C0942101|Carot a-L XRA W contr IA
C0942101|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.left:Document:XR.fluor.angio
C0942101|Views^W contrast IA:Find:Pt:Carotid artery.left:Doc:XR.fluor.angio
C0942105|Spinal artery - right Fluoroscopic angiogram W contrast IA
C0942105|Spinal a-R XRA W contr IA
C0942105|Views^W contrast Intra-arterial:Finding:Point in time:Spinal artery.right:Document:XR.fluor.angio
C0942105|Views^W contrast IA:Find:Pt:Spinal artery.right:Doc:XR.fluor.angio
C0881773|Abdomen retroperitoneum US
C0881773|Abd.reper US
C0881773|Multisection:Finding:Point in time:Abdomen.retroperitoneum:Document:Ultrasound
C0881773|Multisection:Find:Pt:Abdomen.retroperitoneum:Doc:US
C0881785|TA arch XRA W contr IA
C0881785|Aorta arch and Neck Fluoroscopic angiogram W contrast IA
C0881785|Views^W contrast Intra-arterial:Finding:Point in time:Aorta.thoracic.arch:Document:XR.fluor.angio
C0881785|Views^W contrast IA:Find:Pt:Aorta.thoracic.arch:Doc:XR.fluor.angio
C0881801|Abd XR AP (L+R Lat Decub)
C0881801|Abdomen X-ray AP (left lateral-decubitus and right lateral-decubitus)
C0881801|Views AP (L-lateral-decubitus & R-lateral-decubitus):Find:Pt:Abdomen:Doc:XR
C0881801|Views AP (L-lateral-decubitus & R-lateral-decubitus):Finding:Point in time:Abdomen:Document:XR
C0881927|Views:Finding:Point in time:Finger:Narrative:XR
C0881927|Finger XR
C0881927|Finger X-ray
C0881927|Views:Find:Pt:Finger:Doc:XR
C0881927|Views:Finding:Point in time:Finger:Document:XR
C0881964|Vein XRA Atherect guid W contr IV
C0881964|Fluoroscopic angiogram Guidance for atherectomy of Vein-- W contrast IV
C0881964|Guidance for atherectomy^W contrast Intravenous:Finding:Point in time:Vein:Document:XR.fluor.angio
C0881964|Guidance for atherectomy^W contrast IV:Find:Pt:Vein:Doc:XR.fluor.angio
C0881968|Humerus XR 2V
C0881968|Humerus X-ray 2 views
C0881968|Views 2:Finding:Point in time:Humerus:Document:XR
C0881968|Views 2:Find:Pt:Humerus:Doc:XR
C0882005|Knee X-ray 2 views
C0882005|Knee XR 2V
C0882005|Views 2:Find:Pt:Knee:Doc:XR
C0882005|Views 2:Finding:Point in time:Knee:Document:XR
C1114498|Deprecated Kidney - bilateral and Collecting system MRI W and WO contrast IV
C1114498|Deprecated KD-Bl+CS MRI W+WO contr IV
C1114498|Multisection^W & WO contrast IV:Find:Pt:Kidney.bilateral+Collecting system:Nar:MRI
C1114498|Multisection^W & WO contrast Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:MRI
C1114499|L-spine MRI W contr IV
C1114499|Multisection^W contrast Intravenous:Finding:Point in time:Spine.lumbar:Document:MRI
C1114499|Multisection^W contrast IV:Find:Pt:Spine.lumbar:Doc:MRI
C1114499|Lumbar spine MRI W contrast IV
C1114534|Orbit - bilateral X-ray for foreign body
C1114534|Orbit-Bl XR for FB
C1114534|Views for foreign body:Find:Pt:Orbit.bilateral:Doc:XR
C1114534|Views for foreign body:Finding:Point in time:Orbit.bilateral:Document:XR
C1114562|Shoulder X-ray West Point
C1114562|Should XR West Point
C1114562|View West Point:Find:Pt:Shoulder:Doc:XR
C1114562|View West Point:Finding:Point in time:Shoulder:Document:XR
C1114941|T-spine XR AP+Lat
C1114941|Views AP & lateral:Finding:Point in time:Spine.thoracic:Document:XR
C1114941|Views AP & lateral:Find:Pt:Spine.thoracic:Doc:XR
C1114941|Thoracic spine X-ray AP and lateral
C1114599|Multisection:Finding:Point in time:Breast:Narrative:MRI
C1114599|Breast MRI
C1114599|Brst MRI
C1114599|Multisection:Finding:Point in time:Breast:Document:MRI
C1114599|Multisection:Find:Pt:Breast:Doc:MRI
C1114618|Fluoroscopy Guidance for injection of Spine Lumbar Facet Joint
C1114618|L-spine facet joint Flr Inj guid
C1114618|Guidance for injection:Finding:Point in time:Spine.lumbar facet joint:Document:XR.fluor
C1114618|Guidance for injection:Find:Pt:Spine.lumbar facet joint:Doc:XR.fluor
C1114624|IC+Neck ves XRA W contr
C1114624|Intercranial vessel and Neck Vessel Fluoroscopic angiogram W contrast
C1114624|Views^W contrast:Find:Pt:Intracranial vessel+Neck vessel:Doc:XR.fluor.angio
C1114624|Views^W contrast:Finding:Point in time:Intracranial vessel+Neck vessel:Document:XR.fluor.angio
C1114632|Pelvis aa XRA W contr IA
C1114632|Pelvis arteries Fluoroscopic angiogram W contrast IA
C1114632|Views^W contrast IA:Find:Pt:Pelvis arteries:Doc:XR.fluor.angio
C1114632|Views^W contrast Intra-arterial:Finding:Point in time:Pelvis arteries:Document:XR.fluor.angio
C1114634|Deprecated Kidney arteries X-ray fluoroscopy angio W contrast IA
C1114634|Deprecated Flr
C1114634|View^W contrast.XXX IA:Find:Pt:Artery.renal:Nar:XR.fluor
C1114634|View^W contrast.XXX Intra-arterial:Finding:Point in time:Artery.renal:Narrative:XR.fluor
C1114658|Nasopharynx MRI
C1114658|Nasoph MRI
C1114658|Multisection:Find:Pt:Nasopharynx:Doc:MRI
C1114658|Multisection:Finding:Point in time:Nasopharynx:Document:MRI
C1114659|Ac arch+Neck ves MRI.Angio
C1114659|Aortic arch and Neck vessels MRI angiogram
C1114659|Multisection:Find:Pt:Aortic arch+Neck vessels:Doc:MRI.angio
C1114659|Multisection:Finding:Point in time:Aortic arch+Neck vessels:Document:MRI.angio
C1114474|Brst US Bx FN guid
C1114474|US Guidance for fine needle biopsy of Breast
C1114474|Guidance for biopsy.fine needle:Find:Pt:Breast:Doc:US
C1114474|Guidance for biopsy.fine needle:Finding:Point in time:Breast:Document:Ultrasound
C1526826|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast implant.left:Document:MRI
C1526826|Multisection^WO & W contrast IV:Find:Pt:Breast implant.left:Doc:MRI
C1526826|Brst implant-L MRI WO+W contr IV
C1526826|Breast implant - left MRI WO and W contrast IV
C1543749|Views perfusion^W radionuclide Intravenous:Finding:Point in time:Lung:Narrative:Radnuc
C1543749|Lung Scan perfusion
C1543749|Lung RI PF W RNC IV
C1543749|Views perfusion^W radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1543749|Views perfusion^W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1526122|Tib+Fib-R XR Obl
C1526122|Tib+Fib-R XR +Obl
C1526122|Tibia - right and Fibula - right X-ray oblique
C1526122|Tibia - right and Fibula - right X-ray and oblique
C1526122|Views & oblique:Find:Pt:Tibia.right+Fibula.right:Doc:XR
C1526122|Views oblique:Finding:Point in time:Tibia.right+Fibula.right:Document:XR
C1526122|Views oblique:Find:Pt:Tibia.right+Fibula.right:Doc:XR
C1526122|Views & oblique:Finding:Point in time:Tibia.right+Fibula.right:Document:XR
C1542974|RI for Tumor W Tc99mMIBI IV
C1542974|Scan for tumor W Tc-99m Sestamibi IV
C1542974|Views for tumor^W Tc-99m Sestamibi IV:Find:Pt:^Patient:Doc:Radnuc
C1542974|Views for tumor^W Tc-99m Sestamibi Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542979|Thyroid SPECT W I-131 IV
C1542979|Multisection^W I-131 Intravenous:Finding:Point in time:Thyroid:Document:Radnuc.SPECT
C1542979|Multisection^W I-131 IV:Find:Pt:Thyroid:Doc:Radnuc.SPECT
C1543866|Bone marrow Scan static
C1543866|BM RI Static W RNC IV
C1543866|Views static^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc
C1543866|Views static^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc
C1543867|Bone marrow SPECT whole body
C1543867|BM SPECT WB W RNC IV
C1543867|Multisection whole body^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc.SPECT
C1543867|Multisection whole body^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc.SPECT
C1543910|Hrt RI FP+WM W Stress+W RNC IV
C1543910|Heart Scan first pass and wall motion W stress and W radionuclide IV
C1543910|Views first pass & wall motion^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543910|Views first pass & wall motion^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543928|BM SPECT Mul Areas W RNC IV
C1543928|Bone marrow SPECT multiple areas
C1543928|Multisection multiple areas^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc.SPECT
C1543928|Multisection multiple areas^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc.SPECT
C1543941|Hrt RI Gated+FP W RNC IV
C1543941|Heart Scan gated and first pass
C1543941|Views gated & first pass^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543941|Views gated & first pass^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542854|RI for Inf Mul Areas W Ga-67 IV
C1542854|Views for infection multiple areas^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542854|Views for infection multiple areas^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1542854|Scan for infection multiple areas W Ga-67 IV
C1543966|RI Tum local guid Mul Areas W RNC IV
C1543966|Scan Guidance for localization of tumor multiple areas
C1543966|Guidance for localization of tumor multiple areas^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543966|Guidance for localization of tumor multiple areas^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C1543506|Lower extremity vessels - left US.doppler limited
C1543506|LE ves-L DOP Ltd
C1543506|Multisection limited:Find:Pt:Lower extremity vessels.left:Doc:US.doppler
C1543506|Multisection limited:Finding:Point in time:Lower extremity vessels.left:Document:Ultrasound.doppler
C1543150|Multisection^WO & W contrast Intravenous:Finding:Point in time:Orbit+Face:Document:MRI
C1543150|Orbit+Face MRI WO+W contr IV
C1543150|Multisection^WO & W contrast IV:Find:Pt:Orbit+Face:Doc:MRI
C1543150|Orbit and Face MRI WO and W contrast IV
C1543179|Views:Finding:Point in time:Salivary gland:Narrative:XR
C1543179|Salivary gland X-ray
C1543179|Salivary gland XR
C1543179|Views:Find:Pt:Salivary gland:Doc:XR
C1543179|Views:Finding:Point in time:Salivary gland:Document:XR
C1543195|Chest XR AP+Lat+R-Obl+L-Obl
C1543195|Chest X-ray AP and lateral and right oblique and left oblique
C1543195|Views AP & lateral & R-oblique & L-oblique:Find:Pt:Chest:Doc:XR
C1543195|Views AP & lateral & R-oblique & L-oblique:Finding:Point in time:Chest:Document:XR
C1543690|Meckels divertic SPECT W RNC IV
C1543690|Meckels diverticulum SPECT
C1543690|Multisection^W radionuclide IV:Find:Pt:Meckels diverticulum:Doc:Radnuc.SPECT
C1543690|Multisection^W radionuclide Intravenous:Finding:Point in time:Meckels diverticulum:Document:Radnuc.SPECT
C1543711|Hrt SPECT W RNC IV
C1543711|Heart SPECT
C1543711|Multisection^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543711|Multisection^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543714|Hrt RI W DBM+ Tl-201 IV
C1543714|Heart Scan W dobutamine and W Tl-201 IV
C1543714|Views^W dobutamine & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543714|Views^W dobutamine & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1543719|Hrt RI for Infarct W Tc99mPyp IV
C1543719|Heart Scan for infarct W Tc-99m PYP IV
C1543719|Views for infarct^W Tc-99m PYP IV:Find:Pt:Heart:Doc:Radnuc
C1543719|Views for infarct^W Tc-99m PYP Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543729|Hrt RI W Stress+W RNC IV
C1543729|Heart Scan W stress and W radionuclide IV
C1543729|Views^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543729|Views^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543732|RI for Tumor W Ga-67 IV
C1543732|Views for tumor^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543732|Views for tumor^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543732|Scan for tumor W Ga-67 IV
C1526780|Knee-R XR Sunrise 20+40+60 Deg
C1526780|Knee - right X-ray Sunrise 20 and 40 and 60 degrees
C1526780|Views Sunrise 20 & 40 & 60 degrees:Finding:Point in time:Knee.right:Document:XR
C1526780|Views Sunrise 20 & 40 & 60 degrees:Find:Pt:Knee.right:Doc:XR
C1527072|Spine MRI
C1527072|Multisection:Finding:Point in time:Spine:Narrative:MRI
C1527072|Multisection:Finding:Point in time:Spine:Document:MRI
C1527072|Multisection:Find:Pt:Spine:Doc:MRI
C1524815|Multisection^WO contrast:Finding:Point in time:Chest+Abdomen>Aorta:Document:Computerized Tomography
C1524815|Multisection^WO contrast:Find:Pt:Chest+Abdomen>Aorta:Doc:CT
C1524815|Chest+Abd Aorta CT WO contr
C1524815|Chest and Abdomen Aorta CT WO contrast
C1524852|Ft-Bl MRI WO contr
C1524852|Foot - bilateral MRI WO contrast
C1524852|Multisection^WO contrast:Finding:Point in time:Foot.bilateral:Document:MRI
C1524852|Multisection^WO contrast:Find:Pt:Foot.bilateral:Doc:MRI
C1525182|Should ves-L MRI.Angio
C1525182|Shoulder vessels - left MRI angiogram
C1525182|Multisection:Finding:Point in time:Shoulder vessels.left:Document:MRI.angio
C1525182|Multisection:Find:Pt:Shoulder vessels.left:Doc:MRI.angio
C1524237|Pelvis CT limited WO contrast
C1524237|Pelvis CT Ltd WO contr
C1524237|Multisection limited^WO contrast:Find:Pt:Pelvis:Doc:CT
C1524237|Multisection limited^WO contrast:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1524468|Knee CT W contrast IS
C1524468|Multisection^W contrast Intrasynovial:Finding:Point in time:Knee:Document:Computerized Tomography
C1524468|Multisection^W contrast IS:Find:Pt:Knee:Doc:CT
C1524468|Knee CT W contr IS
C1525282|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Adrenal gland:Doc:CT
C1525282|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Adrenal gland:Document:Computerized Tomography
C1525282|Adrenal gland CT WO and W contrast IV
C1525282|Adrenal CT WO+W contr IV
C1525199|LE.L-Veins CT W contr IV
C1525199|Lower extremity - left Veins CT W contrast IV
C1525199|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.left>Veins:Document:Computerized Tomography
C1525199|Multisection^W contrast IV:Find:Pt:Lower extremity.left>Veins:Doc:CT
C1525330|C-spine XR Lat W Flx
C1525330|View lateral^W flexion:Find:Pt:Spine.cervical:Doc:XR
C1525330|View lateral^W flexion:Finding:Point in time:Spine.cervical:Document:XR
C1525330|Cervical spine X-ray lateral W flexion
C1525482|Wrist - left X-ray 4 views
C1525482|Wrist-L XR 4V
C1525482|Views 4:Finding:Point in time:Wrist.left:Document:XR
C1525482|Views 4:Find:Pt:Wrist.left:Doc:XR
C1525532|C-spine XR Lat W FE
C1525532|Views lateral^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C1525532|Views lateral^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C1525532|Cervical spine X-ray lateral W flexion and W extension
C1525577|Superior mesenteric artery Fluoroscopic angiogram W contrast IA
C1525577|SM a XRA W contr IA
C1525577|Views^W contrast IA:Find:Pt:Superior mesenteric artery:Doc:XR.fluor.angio
C1525577|Views^W contrast Intra-arterial:Finding:Point in time:Superior mesenteric artery:Document:XR.fluor.angio
C1525708|Ac arch+Subclavian a XRA W contr IA
C1525708|Aortic arch and Subclavian artery Fluoroscopic angiogram W contrast IA
C1525708|Views^W contrast IA:Find:Pt:Aortic arch+Subclavian artery:Doc:XR.fluor.angio
C1525708|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Subclavian artery:Document:XR.fluor.angio
C1525731|Subclavian a-L XRA W contr IA
C1525731|Subclavian artery - left Fluoroscopic angiogram W contrast IA
C1525731|Views^W contrast IA:Find:Pt:Subclavian artery.left:Doc:XR.fluor.angio
C1525731|Views^W contrast Intra-arterial:Finding:Point in time:Subclavian artery.left:Document:XR.fluor.angio
C1525761|Brain MRI spectroscopy
C1525761|Brain MRI Spectro
C1525761|Multisection spectroscopy:Finding:Point in time:Brain:Document:MRI
C1525761|Multisection spectroscopy:Find:Pt:Brain:Doc:MRI
C1525777|Clavicle - left X-ray 45 degree cephalic angle
C1525777|Clavicle-L XR 45 Deg Ceph Angle
C1525777|View 45 degree cephalic angle:Find:Pt:Clavicle.left:Doc:XR
C1525777|View 45 degree cephalic angle:Finding:Point in time:Clavicle.left:Document:XR
C1525895|Orbit-Bl XR Waters
C1525895|Orbit - bilateral X-ray Waters
C1525895|View Waters:Finding:Point in time:Orbit.bilateral:Document:XR
C1525895|View Waters:Find:Pt:Orbit.bilateral:Doc:XR
C1525971|Scapula X-ray Single view
C1525971|Scapula XR 1V
C1525971|View 1:Finding:Point in time:Scapula:Document:XR
C1525971|View 1:Find:Pt:Scapula:Doc:XR
C1526001|Elbow-R XR AP+Lat+Obl
C1526001|Elbow - right X-ray AP and lateral and oblique
C1526001|Views AP & lateral & oblique:Finding:Point in time:Elbow.right:Document:XR
C1526001|Views AP & lateral & oblique:Find:Pt:Elbow.right:Doc:XR
C1526012|Finger-R XR AP+Lat+Obl
C1526012|Finger - right X-ray AP and lateral and oblique
C1526012|Views AP & lateral & oblique:Finding:Point in time:Finger.right:Document:XR
C1526012|Views AP & lateral & oblique:Find:Pt:Finger.right:Doc:XR
C1526017|Ft-R XR AP+Lat
C1526017|Foot - right X-ray AP and lateral
C1526017|Views AP & lateral:Find:Pt:Foot.right:Doc:XR
C1526017|Views AP & lateral:Finding:Point in time:Foot.right:Document:XR
C1526117|Thumb - right X-ray 3 views
C1526117|Thumb-R XR 3V
C1526117|Views 3:Find:Pt:Thumb.right:Doc:XR
C1526117|Views 3:Finding:Point in time:Thumb.right:Document:XR
C1526147|Sinuses X-ray 4 views
C1526147|Sinuses XR 4V
C1526147|Views 4:Finding:Point in time:Sinuses:Document:XR
C1526147|Views 4:Find:Pt:Sinuses:Doc:XR
C1526149|Sinuses XR Caldwell
C1526149|Sinuses X-ray Caldwell
C1526149|View Caldwell:Find:Pt:Sinuses:Doc:XR
C1526149|View Caldwell:Finding:Point in time:Sinuses:Document:XR
C1526192|Brst-Bl US Bx guid
C1526192|US Guidance for biopsy of Breast - bilateral
C1526192|Guidance for biopsy:Finding:Point in time:Breast.bilateral:Document:Ultrasound
C1526192|Guidance for biopsy:Find:Pt:Breast.bilateral:Doc:US
C1526199|US Guidance for biopsy of Pancreas
C1526199|Pancreas US Bx guid
C1526199|Guidance for biopsy:Find:Pt:Pancreas:Doc:US
C1526199|Guidance for biopsy:Finding:Point in time:Pancreas:Document:Ultrasound
C1526247|Deprecated Calcaneus - bilateral X-ray Broden
C1526247|Views Broden:Find:Pt:Calcaneus.bilateral:Doc:XR
C1526247|Deprecated Heel-Bl XR Broden
C1526247|Views Broden:Finding:Point in time:Calcaneus.bilateral:Document:XR
C1525139|LE-Bl US
C1525139|Lower extremity - bilateral US
C1525139|Multisection:Finding:Point in time:Lower extremity.bilateral:Document:Ultrasound
C1525139|Multisection:Find:Pt:Lower extremity.bilateral:Doc:US
C1524714|Kidney-L US
C1524714|Kidney - left US
C1524714|Multisection:Finding:Point in time:Kidney.left:Document:Ultrasound
C1524714|Multisection:Find:Pt:Kidney.left:Doc:US
C1524715|LE-L US Ltd
C1524715|Lower extremity - left US limited
C1524715|Multisection limited:Finding:Point in time:Lower extremity.left:Document:Ultrasound
C1524715|Multisection limited:Find:Pt:Lower extremity.left:Doc:US
C1526280|Abdomen retroperitoneum US limited
C1526280|Abd.reper US Ltd
C1526280|Multisection limited:Finding:Point in time:Abdomen.retroperitoneum:Document:Ultrasound
C1526280|Multisection limited:Find:Pt:Abdomen.retroperitoneum:Doc:US
C1526288|Multisection^W contrast:Find:Pt:XXX:Doc:US
C1526288|Deprecated Unspecified body region US W contrast
C1526288|Multisection^W contrast:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1526288|Deprecated XXX US W contr
C1525916|Subclavian ves-Bl US
C1525916|Subclavian vessels - bilateral US
C1525916|Multisection:Find:Pt:Subclavian vessels.bilateral:Doc:US
C1525916|Multisection:Finding:Point in time:Subclavian vessels.bilateral:Document:Ultrasound
C1526340|Parotid gland US
C1526340|Multisection:Find:Pt:Parotid gland:Doc:US
C1526340|Multisection:Finding:Point in time:Parotid gland:Document:Ultrasound
C1525147|Finger.2nd-R XR
C1525147|Finger second - right X-ray
C1525147|Views:Finding:Point in time:Finger.second.right:Document:XR
C1525147|Views:Find:Pt:Finger.second.right:Doc:XR
C1526299|Brst implant-Bl Mam
C1526299|Breast implant - bilateral Mammogram
C1526299|Views:Find:Pt:Breast implant.bilateral:Doc:Mam
C1526299|Views:Finding:Point in time:Breast implant.bilateral:Document:Mam
C1526319|Kidney XR W contr Ante
C1526319|Views^W contrast antegrade:Finding:Point in time:Kidney:Document:XR
C1526319|Kidney X-ray W contrast antegrade
C1526319|Views^W contrast antegrade:Find:Pt:Kidney:Doc:XR
C1526330|Parotid gland Flr W contr intra SD
C1526330|Parotid gland Fluoroscopy W contrast intra salivary duct
C1526330|Views^W contrast intra salivary duct:Find:Pt:Parotid gland:Doc:XR.fluor
C1526330|Views^W contrast intra salivary duct:Finding:Point in time:Parotid gland:Document:XR.fluor
C1524473|Multisection^W contrast IS:Find:Pt:Shoulder:Doc:MRI
C1524473|Multisection^W contrast Intrasynovial:Finding:Point in time:Shoulder:Document:MRI
C1524473|Shoulder MRI W contrast IS
C1524473|Should MRI W contr IS
C1524866|Hand-R MRI WO contr
C1524866|Hand - right MRI WO contrast
C1524866|Multisection^WO contrast:Find:Pt:Hand.right:Doc:MRI
C1524866|Multisection^WO contrast:Finding:Point in time:Hand.right:Document:MRI
C1524172|Hip-R MRI W contr IV
C1524172|Hip - right MRI W contrast IV
C1524172|Multisection^W contrast IV:Find:Pt:Hip.right:Doc:MRI
C1524172|Multisection^W contrast Intravenous:Finding:Point in time:Hip.right:Document:MRI
C1524925|Neck vessels MRI angiogram WO contrast
C1524925|Neck ves MRI.Angio WO contr
C1524925|Multisection^WO contrast:Finding:Point in time:Neck vessels:Document:MRI.angio
C1524925|Multisection^WO contrast:Find:Pt:Neck vessels:Doc:MRI.angio
C1524553|Kidney - bilateral MRI W contrast IV
C1524553|Multisection^W contrast IV:Find:Pt:Kidney.bilateral:Doc:MRI
C1524553|Multisection^W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:MRI
C1524553|Kdny-Bl MRI W contr IV
C1524577|Post fossa MRI W contr IV
C1524577|Posterior fossa MRI W contrast IV
C1524577|Multisection^W contrast IV:Find:Pt:Posterior fossa:Doc:MRI
C1524577|Multisection^W contrast Intravenous:Finding:Point in time:Posterior fossa:Document:MRI
C1524931|Lower extremity - bilateral X-ray Single view
C1524931|LE-Bl XR 1V
C1524931|View 1:Find:Pt:Lower extremity.bilateral:Doc:XR
C1524931|View 1:Finding:Point in time:Lower extremity.bilateral:Document:XR
C1524209|Ft XR AP 1V
C1524209|Foot X-ray AP single view
C1524209|View AP:Finding:Point in time:Foot:Document:XR
C1524209|View AP:Find:Pt:Foot:Doc:XR
C1524602|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ankle:Document:Computerized Tomography
C1524602|Ankle CT WO and W contrast IV
C1524602|Ankle CT WO+W contr IV
C1524602|Multisection^WO & W contrast IV:Find:Pt:Ankle:Doc:CT
C1524958|Finger.5th XR Obl 1V
C1524958|Finger fifth X-ray oblique single view
C1524958|View oblique:Find:Pt:Finger.fifth:Doc:XR
C1524958|View oblique:Finding:Point in time:Finger.fifth:Document:XR
C1524984|Knee-L XR
C1524984|Knee - left X-ray
C1524984|Views:Find:Pt:Knee.left:Doc:XR
C1524984|Views:Finding:Point in time:Knee.left:Document:XR
C1524321|CT Guidance for drainage of Unspecified body region
C1524321|XXX CT Drain guid
C1524321|Guidance for drainage:Find:Pt:XXX:Doc:CT
C1524321|Guidance for drainage:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1524331|L-spine CT Nerve Block guid
C1524331|Guidance for nerve block:Find:Pt:Spine.lumbar:Doc:CT
C1524331|Guidance for nerve block:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1524331|CT Guidance for nerve block of Lumbar spine
C1524154|Finger - left X-ray 2 views
C1524154|Finger-L XR 2V
C1524154|Views 2:Finding:Point in time:Finger.left:Document:XR
C1524154|Views 2:Find:Pt:Finger.left:Doc:XR
C1527018|Elbow CT
C1527018|Multisection:Finding:Point in time:Elbow:Document:Computerized Tomography
C1527018|Multisection:Find:Pt:Elbow:Doc:CT
C1524388|Foot - left X-ray tomograph
C1524388|Ft-L XRTomo
C1524388|Multisection:Finding:Point in time:Foot.left:Document:XR.tomo
C1524388|Multisection:Find:Pt:Foot.left:Doc:XR.tomo
C1524748|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip.left:Document:Computerized Tomography
C1524748|Multisection^WO & W contrast IV:Find:Pt:Hip.left:Doc:CT
C1524748|Hip - left CT WO and W contrast IV
C1524748|Hip-L CT WO+W contr IV
C1524765|Knee CT WO and W contrast IV
C1524765|Knee CT WO+W contr IV
C1524765|Multisection^WO & W contrast IV:Find:Pt:Knee:Doc:CT
C1524765|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee:Document:Computerized Tomography
C1525063|Elbow-L XR AP+Lat+Obl
C1525063|Elbow - left X-ray AP and lateral and oblique
C1525063|Views AP & lateral & oblique:Find:Pt:Elbow.left:Doc:XR
C1525063|Views AP & lateral & oblique:Finding:Point in time:Elbow.left:Document:XR
C1525064|Finger XR AP+Lat+Obl
C1525064|Finger X-ray AP and lateral and oblique
C1525064|Views AP & lateral & oblique:Find:Pt:Finger:Doc:XR
C1525064|Views AP & lateral & oblique:Finding:Point in time:Finger:Document:XR
C1524415|Upper arm - bilateral CT
C1524415|Upper arm-Bl CT
C1524415|Multisection:Find:Pt:Upper arm.bilateral:Doc:CT
C1524415|Multisection:Finding:Point in time:Upper arm.bilateral:Document:Computerized Tomography
C1524774|Prostate MRI WO and W contrast IV
C1524774|Prostate MRI WO+W contr IV
C1524774|Multisection^WO & W contrast Intravenous:Finding:Point in time:Prostate:Document:MRI
C1524774|Multisection^WO & W contrast IV:Find:Pt:Prostate:Doc:MRI
C1830234|Breast - unilateral MRI WO contrast
C1830234|Brst-UL MRI WO contr
C1830234|Multisection^WO contrast:Find:Pt:Breast.unilateral:Doc:MRI
C1830234|Multisection^WO contrast:Finding:Point in time:Breast.unilateral:Document:MRI
C1830264|Lower extremity vein US
C1830264|LE v US
C1830264|Multisection:Find:Pt:Lower extremity vein:Doc:US
C1830264|Multisection:Finding:Point in time:Lower extremity vein:Document:Ultrasound
C1830269|CT Guidance for needle biopsy of Breast
C1830269|Brst CT Bx needle guid
C1830269|Guidance for biopsy.needle:Find:Pt:Breast:Doc:CT
C1830269|Guidance for biopsy.needle:Finding:Point in time:Breast:Document:Computerized Tomography
C1830093|Upper extremity vessels - bilateral US.doppler
C1830093|UE ves-Bl DOP
C1830093|Multisection:Find:Pt:Upper extremity vessels.bilateral:Doc:US.doppler
C1830093|Multisection:Finding:Point in time:Upper extremity vessels.bilateral:Document:Ultrasound.doppler
C1715375|CT Guidance for fine needle aspiration of Lymph node
C1715375|LN CT FNA Asp
C1715375|Guidance for aspiration.fine needle:Finding:Point in time:Lymph node:Document:Computerized Tomography
C1715375|Guidance for aspiration.fine needle:Find:Pt:Lymph node:Doc:CT
C1715383|Multisection^WO & W contrast Intravenous:Finding:Point in time:Skull.base:Document:Computerized Tomography
C1715383|Skull.base CT WO+W contr IV
C1715383|Skull.base CT WO and W contrast IV
C1715383|Multisection^WO & W contrast IV:Find:Pt:Skull.base:Doc:CT
C1717316|Liver US Bx needle guid
C1717316|US Guidance for needle biopsy of Liver
C1717316|Guidance for biopsy.needle:Find:Pt:Liver:Doc:US
C1717316|Guidance for biopsy.needle:Finding:Point in time:Liver:Document:Ultrasound
C1715444|Sacrum+Coccyx XR 2V
C1715444|Sacrum and Coccyx X-ray 2 views
C1715444|Views 2:Find:Pt:Sacrum+Coccyx:Doc:XR
C1715444|Views 2:Finding:Point in time:Sacrum+Coccyx:Document:XR
C1715459|L-spine XR GE 5V W R+L-bending
C1715459|Views GE 5^W R-Bending & W L-Bending:Find:Pt:Spine.lumbar:Doc:XR
C1715459|Views GE 5^W R-Bending & W L-Bending:Finding:Point in time:Spine.lumbar:Document:XR
C1715459|Lumbar spine X-ray GE 5 views W right bending and W left bending
C2729168|Orbit CT
C2729168|Multisection:Finding:Point in time:Head>Orbit:Document:Computerized Tomography
C2729168|Multisection:Find:Pt:Head>Orbit:Doc:CT
C1649482|Elbow - left X-ray portable
C1649482|Elbow-L XR port
C1649482|Views portable:Finding:Point in time:Elbow.left:Document:XR
C1649482|Views portable:Find:Pt:Elbow.left:Doc:XR
C1632798|L-spine XR AP 1V W R-bending
C1632798|View AP^W R-bending:Find:Pt:Spine.lumbar:Doc:XR
C1632798|View AP^W R-bending:Finding:Point in time:Spine.lumbar:Document:XR
C1632798|Lumbar spine X-ray AP single view W right bending
C1714815|BD+PDs Flr Endo guid 1.5h p contr retro
C1714815|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 1.5 hours post contrast retrograde
C1714815|Guidance for endoscopy^1 1/2 hour post contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1714815|Guidance for endoscopy^1.5H post contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1705862|Finger.2nd-R XR GE 3V
C1705862|Finger second - right X-ray GE 3 views
C1705862|Finger second - right Narrative X-ray GE 3 views
C1705862|Views GE 3:Finding:Point in time:Finger.second.right:Document:XR
C1705862|Views GE 3:Find:Pt:Finger.second.right:Doc:XR
C1717267|Brain RI Flow W Tc99mDTPA IV
C1717267|Brain Scan flow W Tc-99m DTPA IV
C1717267|Views flow^W Tc-99m DTPA IV:Find:Pt:Brain:Doc:Radnuc
C1717267|Views flow^W Tc-99m DTPA Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1715023|Liver+BDs+GB RI W Sinc+RNC IV
C1715023|Liver and Biliary ducts and Gallbladder Scan W sincalide and W radionuclide IV
C1715023|Views^W sincalide & W radionuclide IV:Find:Pt:Liver+Biliary ducts+Gallbladder:Doc:Radnuc
C1715023|Views^W sincalide & W radionuclide Intravenous:Finding:Point in time:Liver+Biliary ducts+Gallbladder:Document:Radnuc
C1714500|KD-Bl+Renal ves RI Flow W Tc99mGHA IV
C1714500|Views flow^W Tc-99m glucoheptonate IV:Find:Pt:Kidney.bilateral+Renal vessels:Doc:Radnuc
C1714500|Kidney - bilateral and Renal vessels Scan flow W Tc-99m glucoheptonate IV
C1714500|Views flow^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Kidney.bilateral+Renal vessels:Document:Radnuc
C1715096|Multisection^WO & W contrast Intravenous:Finding:Point in time:Kidney:Document:Computerized Tomography
C1715096|Kidney CT WO+W contr IV
C1715096|Multisection^WO & W contrast IV:Find:Pt:Kidney:Doc:CT
C1715096|Kidney CT WO and W contrast IV
C1715106|Knee XR Sunrise
C1715106|Knee X-ray Sunrise
C1715106|View Sunrise:Find:Pt:Knee:Doc:XR
C1715106|View Sunrise:Finding:Point in time:Knee:Document:XR
C1640449|Carot a DOP
C1640449|Carotid artery US.doppler
C1640449|Multisection:Finding:Point in time:Carotid artery:Document:Ultrasound.doppler
C1640449|Multisection:Find:Pt:Carotid artery:Doc:US.doppler
C1627297|L-spine XR +Obl
C1627297|Views & oblique:Finding:Point in time:Spine.lumbar:Document:XR
C1627297|Views & oblique:Find:Pt:Spine.lumbar:Doc:XR
C1627297|Lumbar spine X-ray and oblique
C1626176|RI for Tumor WB W RNC IV
C1626176|Scan for tumor whole body
C1626176|Views for tumor whole body^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1626176|Views for tumor whole body^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C2361224|CT Guidance for replacement of percutaneous drainage tube in Pelvis
C2361224|Pelvis CT Replac of PC drain tube guid
C2361224|Guidance for replacement of percutaneous drainage tube:Finding:Point in time:Pelvis:Document:Computerized Tomography
C2361224|Guidance for replacement of percutaneous drainage tube:Find:Pt:Pelvis:Doc:CT
C3261217|XXX Image ID
C3261217|Image ID:ID:Pt:XXX:Nom
C3261217|Unspecified body region Image ID
C3261217|Image ID:Identifier:Point in time:To be specified in another part of the message:Nominal
C3533568|US Guidance for laser ablation of vein(s) of Extremity vein - right
C3533568|Guidance for laser ablation of vein(s):Find:Pt:Extremity vein.right:Doc:US
C3533568|Guidance for laser ablation of vein(s):Finding:Point in time:Extremity vein.right:Document:Ultrasound
C3533568|Extr v-R US Laser ablation guid
C3262977|Breast implant X-ray diagnostic
C3262977|Brst implant XR Dx
C3262977|Views diagnostic:Finding:Point in time:Breast implant:Document:XR
C3262977|Views diagnostic:Find:Pt:Breast implant:Doc:XR
C3483133|C-spine US CSF asp guid
C3483133|Guidance for CSF aspiration:Finding:Point in time:Spine.cervical:Document:Ultrasound
C3483133|Guidance for CSF aspiration:Find:Pt:Spine.cervical:Doc:US
C3483133|US Guidance for CSF aspiration of Cervical spine
C3263017|MRI Guidance for needle biopsy of Liver
C3263017|Liver MRI Bx needle guid
C3263017|Guidance for biopsy.needle:Find:Pt:Liver:Doc:MRI
C3263017|Guidance for biopsy.needle:Finding:Point in time:Liver:Document:MRI
C3263033|Skull.base MRI WO+W contr IV
C3263033|Multisection^WO & W contrast Intravenous:Finding:Point in time:Skull.base:Document:MRI
C3263033|Multisection^WO & W contrast IV:Find:Pt:Skull.base:Doc:MRI
C3263033|Skull.base MRI WO and W contrast IV
C3263050|SPECT for Tumor WB W RNC IV
C3263050|SPECT for tumor whole body
C3263050|Multisection for tumor whole body^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C3263050|Multisection for tumor whole body^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C3261720|Eye US limited
C3261720|Eye US Ltd
C3261720|Multisection limited:Find:Pt:Eye:Doc:US
C3261720|Multisection limited:Finding:Point in time:Eye:Document:Ultrasound
C3262887|Knee-Bl XR Sunrise+(views Stand)
C3262887|Knee - bilateral X-ray Sunrise and (views standing)
C3262887|View Sunrise & (views^standing):Finding:Point in time:Knee.bilateral:Document:XR
C3262887|View Sunrise & (views^standing):Find:Pt:Knee.bilateral:Doc:XR
C3262893|Ribs - bilateral X-ray anterior and lateral
C3262893|Ribs-Bl XR Ant+Lat
C3262893|Views anterior & lateral:Find:Pt:Ribs.bilateral:Doc:XR
C3262893|Views anterior & lateral:Finding:Point in time:Ribs.bilateral:Document:XR
C0942239|Finger - right MRI
C0942239|Finger-R MRI
C0942239|Multisection:Finding:Point in time:Finger.right:Document:MRI
C0942239|Multisection:Find:Pt:Finger.right:Doc:MRI
C0942249|IAC-L XRTomo
C0942249|Internal auditory canal - left X-ray tomograph
C0942249|Multisection:Finding:Point in time:Internal auditory canal.left:Document:XR.tomo
C0942249|Multisection:Find:Pt:Internal auditory canal.left:Doc:XR.tomo
C0942265|Shoulder - right MRI
C0942265|Should-R MRI
C0942265|Multisection:Finding:Point in time:Shoulder.right:Document:MRI
C0942265|Multisection:Find:Pt:Shoulder.right:Doc:MRI
C0942305|Brst-R US Needle local guid
C0942305|US Guidance for needle localization of Breast - right
C0942305|Guidance for needle localization:Find:Pt:Breast.right:Doc:US
C0942305|Guidance for needle localization:Finding:Point in time:Breast.right:Document:Ultrasound
C0942313|US Guidance for drainage of Extremity - left
C0942313|Extr-L US Drain guid
C0942313|Guidance for drainage:Finding:Point in time:Extremity.left:Document:Ultrasound
C0942313|Guidance for drainage:Find:Pt:Extremity.left:Doc:US
C0945343|Hand - right X-ray arthritis
C0945343|Hand-R XR Arthritis
C0945343|View arthritis:Find:Pt:Hand.right:Doc:XR
C0945343|View arthritis:Finding:Point in time:Hand.right:Document:XR
C0942363|Should-R XR 3V
C0942363|Shoulder - right X-ray 3 views
C0942363|Views 3:Find:Pt:Shoulder.right:Doc:XR
C0942363|Views 3:Finding:Point in time:Shoulder.right:Document:XR
C0942367|Hand - bilateral X-ray 2 views
C0942367|Hand-Bl XR 2V
C0942367|Views 2:Finding:Point in time:Hand.bilateral:Document:XR
C0942367|Views 2:Find:Pt:Hand.bilateral:Doc:XR
C0882034|Multisection^WO & W contrast IV:Find:Pt:Neck:Doc:MRI
C0882034|Neck MRI WO+W contr IV
C0882034|Neck MRI WO and W contrast IV
C0882034|Multisection^WO & W contrast Intravenous:Finding:Point in time:Neck:Document:MRI
C0882042|Orbit - bilateral CT WO and W contrast IV
C0882042|Orbit-Bl CT WO+W contr IV
C0882042|Multisection^WO & W contrast IV:Find:Pt:Head>Orbit.bilateral:Doc:CT
C0882042|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head>Orbit.bilateral:Document:Computerized Tomography
C0882061|Pelvis vessels US.doppler
C0882061|Pelvis ves DOP
C0882061|Multisection:Finding:Point in time:Pelvis vessels:Document:Ultrasound.doppler
C0882061|Multisection:Find:Pt:Pelvis vessels:Doc:US.doppler
C0882064|Periph aa XRA W contr IA
C0882064|Peripheral arteries Fluoroscopic angiogram W contrast IA
C0882064|Views^W contrast IA:Find:Pt:Peripheral arteries:Doc:XR.fluor.angio
C0882064|Views^W contrast Intra-arterial:Finding:Point in time:Peripheral arteries:Document:XR.fluor.angio
C0882547|Popliteal space US
C0882547|Multisection:Find:Pt:Popliteal space:Doc:US
C0882547|Multisection:Finding:Point in time:Popliteal space:Document:Ultrasound
C0882548|Deprecated Pulmonary artery Bilateral X-ray fluoroscopy angio W contrast IA
C0882548|Deprecated PAA XRA
C0882548|Views^W contrast in pulmonary artery:Find:Pt:Pulmonary arteries:Nar:XR.fluor.angio
C0882548|Views^W contrast in pulmonary artery:Finding:Point in time:Pulmonary arteries:Narrative:XR.fluor.angio
C0882549|Rectum US
C0882549|Multisection:Find:Pt:Rectum:Doc:US
C0882549|Multisection:Finding:Point in time:Rectum:Document:Ultrasound
C0882094|Shunt Flr
C0882094|Shunt Fluoroscopy
C0882094|Views:Finding:Point in time:Shunt.To be specified in another part of the message:Document:XR.fluor
C0882094|Views:Find:Pt:Shunt.XXX:Doc:XR.fluor
C0882154|Views:Finding:Point in time:Sternum:Narrative:XR
C0882154|Sternum X-ray
C0882154|Sternum XR
C0882154|Views:Find:Pt:Sternum:Doc:XR
C0882154|Views:Finding:Point in time:Sternum:Document:XR
C0882168|Thyroid US
C0882168|Multisection:Find:Pt:Thyroid:Doc:US
C0882168|Multisection:Finding:Point in time:Thyroid:Document:Ultrasound
C0882561|Urinary Bladder and Urethra Fluoroscopy W contrast intra bladder
C0882561|Views^W contrast intra bladder:Finding:Point in time:Urinary bladder+Urethra:Document:XR.fluor
C0882561|Views^W contrast intra bladder:Find:Pt:Urinary bladder+Urethra:Doc:XR.fluor
C0882561|Bladder+Urethra Flr W contr IUB
C0942097|Views^W contrast IS:Find:Pt:Knee.right:Doc:XR.fluor
C0942097|Knee - right Fluoroscopy W contrast IS
C0942097|Knee-R Flr W contr IS
C0942097|Views^W contrast Intrasynovial:Finding:Point in time:Knee.right:Document:XR.fluor
C0942106|Knee - bilateral X-ray standing
C0942106|Knee-Bl XR stand
C0942106|Views^standing:Find:Pt:Knee.bilateral:Doc:XR
C0942106|Views^standing:Finding:Point in time:Knee.bilateral:Document:XR
C0942108|Knee - right X-ray standing
C0942108|Knee-R XR stand
C0942108|Views^standing:Find:Pt:Knee.right:Doc:XR
C0942108|Views^standing:Finding:Point in time:Knee.right:Document:XR
C0942129|Elbow-R XR
C0942129|Elbow - right X-ray
C0942129|Views:Finding:Point in time:Elbow.right:Document:XR
C0942129|Views:Find:Pt:Elbow.right:Doc:XR
C0945312|Finger - bilateral X-ray
C0945312|Finger-Bl XR
C0945312|Views:Finding:Point in time:Finger.bilateral:Document:XR
C0945312|Views:Find:Pt:Finger.bilateral:Doc:XR
C0942147|Acetabulum - right X-ray
C0942147|Acetabulum-R XR
C0942147|Views:Finding:Point in time:Acetabulum.right:Document:XR
C0942147|Views:Find:Pt:Acetabulum.right:Doc:XR
C0881823|Brain MRI W anesthesia
C0881823|Multisection^W anesthesia:Find:Pt:Brain:Doc:MRI
C0881823|Multisection^W anesthesia:Finding:Point in time:Brain:Document:MRI
C0881830|Brst Mam Cyst Asp guid
C0881830|Mammogram Guidance for aspiration of cyst of Breast
C0881830|Guidance for aspiration of cyst:Find:Pt:Breast:Doc:Mam
C0881830|Guidance for aspiration of cyst:Finding:Point in time:Breast:Document:Mam
C0881833|Breast specimen Mammogram
C0881833|Brst specimen Mam
C0881833|Views:Finding:Point in time:Breast specimen:Document:Mam
C0881833|Views:Find:Pt:Breast specimen:Doc:Mam
C0881836|Brst US
C0881836|Breast US
C0881836|Multisection:Finding:Point in time:Breast:Document:Ultrasound
C0881836|Multisection:Find:Pt:Breast:Doc:US
C0881864|Chest XR port W insp+exp
C0881864|Chest X-ray portable W inspiration and expiration
C0881864|Views portable^W inspiration & expiration:Finding:Point in time:Chest:Document:XR
C0881864|Views portable ^W inspiration & expiration:Find:Pt:Chest:Doc:XR
C0881867|Chest XR L-Lat Upr port
C0881867|Chest X-ray left lateral upright portable
C0881867|View L-lateral upright portable:Finding:Point in time:Chest:Document:XR
C0881867|View L-lateral upright portable:Find:Pt:Chest:Doc:XR
C0881941|Hand X-ray arthritis
C0881941|Hand XR Arthritis
C0881941|View arthritis:Finding:Point in time:Hand:Document:XR
C0881941|View arthritis:Find:Pt:Hand:Doc:XR
C0882535|Multisection:Finding:Point in time:Coronary arteries:Document:Computerized Tomography.fast
C0882535|Deprecated Coronary arteries CT fast
C0882535|Multisection:Find:Pt:Coronary arteries:Doc:CT.fast
C0882535|Deprecated Coronary aa CT.Fast
C0881979|Fluoroscopy Guidance for placement of percutaneous nephrostomy in Kidney - bilateral-- W contrast via tube
C0881979|Guidance for placement of percutaneous nephrostomy^W contrast via tube:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C0881979|Guidance for placement of percutaneous nephrostomy^W contrast via tube:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C0881979|Kdny-Bl Flr PN guid W contr via tb
C0881986|Deprecated Kidney Bilateral & Collecting system X-ray tomograph Multisection W & WO contrast IV
C0881986|Deprecated KD-Bl+CS XR.Tomo W+WO contr I
C0881986|Multisection^W & WO contrast IV:Find:Pt:Kidney.bilateral+Collecting system:Nar:XR.tomo
C0881986|Multisection^W & WO contrast Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:XR.tomo
C0881986|Deprecated KDs+CS XR.Tomo W+WO contr IV
C1114526|Hip US WO developmental joint assessment
C1114526|Hip US WO devel joint assess
C1114526|Multisection^WO developmental joint assessment:Find:Pt:Hip:Doc:US
C1114526|Multisection^WO developmental joint assessment:Finding:Point in time:Hip:Document:Ultrasound
C1114542|Views^flexion & extension:Find:Pt:Spine.cervical:Nar:XR
C1114542|Deprecated C-spine XR
C1114542|Deprecated Spine Cervical X-ray W flexion & W extension
C1114542|Views^flexion & extension:Finding:Point in time:Spine.cervical:Narrative:XR
C1114607|Multisection^WO & W contrast IV:Find:Pt:Chest>Vessels:Doc:CT.angio
C1114607|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest>Vessels:Document:Computerized Tomography.angio
C1114607|Chest Ves CT.Angio WO+W contr IV
C1114607|Chest vessels CT angiogram WO and W contrast IV
C1114616|BD+PDs Flr Endo guid W contr retro
C1114616|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- W contrast retrograde
C1114616|Guidance for endoscopy^W contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1114616|Guidance for endoscopy^W contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1114630|PA-Bl XRA W contr IA
C1114630|Pulmonary artery - bilateral Fluoroscopic angiogram W contrast IA
C1114630|Views^W contrast Intra-arterial:Finding:Point in time:Pulmonary artery.bilateral:Document:XR.fluor.angio
C1114630|Views^W contrast IA:Find:Pt:Pulmonary artery.bilateral:Doc:XR.fluor.angio
C1114644|IVC XRA W contr IV
C1114644|Inferior vena cava Fluoroscopic angiogram W contrast IV
C1114644|Views^W contrast IV:Find:Pt:Vena cava.inferior:Doc:XR.fluor.angio
C1114644|Views^W contrast Intravenous:Finding:Point in time:Vena cava.inferior:Document:XR.fluor.angio
C1114648|Extr aa-Bl XRA W contr IA
C1114648|Extremity arteries - bilateral Fluoroscopic angiogram W contrast IA
C1114648|Views^W contrast Intra-arterial:Finding:Point in time:Extremity arteries.bilateral:Document:XR.fluor.angio
C1114648|Views^W contrast IA:Find:Pt:Extremity arteries.bilateral:Doc:XR.fluor.angio
C1114661|Abd vv+IVC MRI.Angio
C1114661|Abdominal veins and IVC MRI angiogram
C1114661|Multisection:Find:Pt:Abdominal veins+Vena cava.inferior:Doc:MRI.angio
C1114661|Multisection:Finding:Point in time:Abdominal veins+Vena cava.inferior:Document:MRI.angio
C1114923|Petrous part of temporal bone CT WO contrast
C1114923|Multisection^WO contrast:Finding:Point in time:Petrous part of temporal bone:Document:Computerized Tomography
C1114923|Multisection^WO contrast:Find:Pt:Petrous part of temporal bone:Doc:CT
C1114923|Petr part temp bone CT WO contr
C1114925|Multisection^W positive contrast via enteroclysis tube:Find:Pt:Small bowel:Doc:CT
C1114925|Small bowel CT W positive contrast via enteroclysis tube
C1114925|Multisection^W positive contrast via enteroclysis tube:Finding:Point in time:Small bowel:Document:Computerized Tomography
C1114925|SB CT W Pos Cntrst Enteroclysis Tube
C1114456|Fluoroscopy Guidance for procedure of Unspecified body region
C1114456|XXX Flr Procedure guid
C1114456|Guidance for procedure:Find:Pt:XXX:Doc:XR.fluor
C1114456|Guidance for procedure:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1114462|Colon Fluoroscopy Reduction W views W contrast PR
C1114462|Colon Flr Reduction W views W contr PR
C1114462|Reduction W views^W contrast PR:Find:Pt:Colon:Doc:XR.fluor
C1114462|Reduction W views^W contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C1114464|Vessel Fluoroscopic angiogram W contrast
C1114464|View^W contrast:Find:Pt:Vessel:Doc:XR.fluor.angio
C1114464|View^W contrast:Finding:Point in time:Vessel:Document:XR.fluor.angio
C1114464|Vesl XRA W contr
C1526827|Knee-L XR 2V Obl
C1526827|Knee - left X-ray 2 views Oblique
C1526827|Views 2 oblique:Finding:Point in time:Knee.left:Document:XR
C1526827|Views 2 oblique:Find:Pt:Knee.left:Doc:XR
C1114946|Pelvis XR +Inlet+Outlet
C1114946|Pelvis XR Inlet+Outlet
C1114946|Pelvis X-ray inlet and outlet
C1114946|Pelvis X-ray and inlet and outlet
C1114946|Views inlet & outlet:Find:Pt:Pelvis:Doc:XR
C1114946|Views inlet & outlet:Finding:Point in time:Pelvis:Document:XR
C1114946|Views & inlet & outlet:Find:Pt:Pelvis:Doc:XR
C1114946|Views & inlet & outlet:Finding:Point in time:Pelvis:Document:XR
C1543764|Heart SPECT perfusion
C1543764|Hrt SPECT PF W RNC IV
C1543764|Multisection perfusion^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543764|Multisection perfusion^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543775|Hrt SPECT PF Rest+stress+W Tl201 IV
C1543775|Heart SPECT perfusion at rest and W stress and W Tl-201 IV
C1543775|Multisection perfusion^at rest & W stress & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543775|Multisection perfusion^at rest & W stress & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1955478|T-spine XR +Obl
C1955478|Views & oblique:Finding:Point in time:Spine.thoracic:Document:XR
C1955478|Views & oblique:Find:Pt:Spine.thoracic:Doc:XR
C1955478|Thoracic spine X-ray and oblique
C1543494|Extremity vein - bilateral US.doppler
C1543494|Extr v-Bl DOP
C1543494|Multisection:Find:Pt:Extremity vein.bilateral:Doc:US.doppler
C1543494|Multisection:Finding:Point in time:Extremity vein.bilateral:Document:Ultrasound.doppler
C1542978|Thyroid RI Ltd W I-131 IV
C1542978|Thyroid Scan limited W I-131 IV
C1542978|Views limited^W I-131 IV:Find:Pt:Thyroid:Doc:Radnuc
C1542978|Views limited^W I-131 Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1542897|Lung Scan ventilation W radionuclide aerosol IH
C1542897|Views ventilation^W radionuclide aerosol Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1542897|Lung RI V W RNC Aero IH
C1542897|Views ventilation^W radionuclide aerosol IH:Find:Pt:Lung:Doc:Radnuc
C1542921|Hrt RI FP Rest+W Tc99mMIBI IV
C1542921|Heart Scan first pass at rest and W Tc-99m Sestamibi IV
C1542921|Views first pass^at rest & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542921|Views first pass^at rest & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543899|Liver+Spleen RI W RNC IV
C1543899|Liver and Spleen Scan
C1543899|Views^W radionuclide IV:Find:Pt:Liver+Spleen:Doc:Radnuc
C1543899|Views^W radionuclide Intravenous:Finding:Point in time:Liver+Spleen:Document:Radnuc
C1543900|Liver+Spleen RI Static W RNC IV
C1543900|Liver and Spleen Scan static
C1543900|Views static^W radionuclide IV:Find:Pt:Liver+Spleen:Doc:Radnuc
C1543900|Views static^W radionuclide Intravenous:Finding:Point in time:Liver+Spleen:Document:Radnuc
C1543907|Hrt RI FP+VV W RNC IV
C1543907|Heart Scan first pass and ventricular volume
C1543907|Views first pass & ventricular volume^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543907|Views first pass & ventricular volume^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543944|Hrt RI Gated Rest+W Tc-99mP IV
C1543944|Heart Scan gated at rest and W Tc-99m pertechnetate IV
C1543944|Views gated^at rest & W Tc-99m pertechnetate IV:Find:Pt:Heart:Doc:Radnuc
C1543944|Views gated^at rest & W Tc-99m pertechnetate Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542851|Hrt SPECT Gated W Stress+W RNC IV
C1542851|Heart SPECT gated W stress and W radionuclide IV
C1542851|Multisection gated^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1542851|Multisection gated^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543952|Joint RI W RNC IV
C1543952|Joint Scan
C1543952|Views^W radionuclide IV:Find:Pt:Joint:Doc:Radnuc
C1543952|Views^W radionuclide Intravenous:Finding:Point in time:Joint:Document:Radnuc
C1543956|Lung RI VP W RNC IH+Particulate IV
C1543956|Views ventilation & perfusion^W radionuclide IH & W particulate radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1543956|Lung Scan ventilation and perfusion W radionuclide IH and W particulate radionuclide IV
C1543956|Views ventilation & perfusion^W radionuclide Inhalation & W particulate radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1524718|Chest X-ray Diameter.lateral
C1524718|Diameter.lateral:Len:Pt:Chest:Qn:XR
C1524718|Chest XR Diam Lat
C1524718|Diameter.lateral:Length:Point in time:Chest:Quantitative:XR
C1543497|LE a-Bl DOP
C1543497|Lower extremity artery - bilateral US.doppler
C1543497|Multisection:Finding:Point in time:Lower extremity artery.bilateral:Document:Ultrasound.doppler
C1543497|Multisection:Find:Pt:Lower extremity artery.bilateral:Doc:US.doppler
C1543505|Extr v-L DOP
C1543505|Extremity vein - left US.doppler
C1543505|Multisection:Find:Pt:Extremity vein.left:Doc:US.doppler
C1543505|Multisection:Finding:Point in time:Extremity vein.left:Document:Ultrasound.doppler
C1543527|Guidance for drainage of abscess:Find:Pt:XXX:Doc:US
C1543527|Guidance for drainage of abscess:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1543527|XXX US Abscess drain guid
C1543527|US Guidance for drainage of abscess of Unspecified body region
C1543573|Iliac ves DOP
C1543573|Iliac vessels US.doppler
C1543573|Multisection:Finding:Point in time:Iliac vessels:Document:Ultrasound.doppler
C1543573|Multisection:Find:Pt:Iliac vessels:Doc:US.doppler
C1543589|Hip-R XR Danelius Miller
C1543589|Hip - right X-ray Danelius Miller
C1543589|View Danelius Miller:Find:Pt:Hip.right:Doc:XR
C1543589|View Danelius Miller:Finding:Point in time:Hip.right:Document:XR
C1525161|US Guidance for biopsy of Liver transplant
C1525161|Liver Transplant US Bx guid
C1525161|Guidance for biopsy:Find:Pt:Liver transplant:Doc:US
C1525161|Guidance for biopsy:Finding:Point in time:Liver transplant:Document:Ultrasound
C1543726|Hrt RI for Shunt Det W Tc99mMAA IV
C1543726|Heart Scan for shunt detection W Tc-99m MAA IV
C1543726|Views for shunt detection^W Tc-99m MAA Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543726|Views for shunt detection^W Tc-99m MAA IV:Find:Pt:Heart:Doc:Radnuc
C1526779|Views magnification & spot^compression:Find:Pt:Breast.right:Nar:Mam
C1526779|Views magnification & spot^compression:Finding:Point in time:Breast.right:Narrative:Mam
C1526779|Deprecated Breast - right Mammogram magnification & spot compression
C1526779|Deprecated Brst-R Mam Mag+Spot Compressi
C1526806|LE-L XR stand
C1526806|Lower extremity - left X-ray standing
C1526806|View^standing:Find:Pt:Lower extremity.left:Doc:XR
C1526806|View^standing:Finding:Point in time:Lower extremity.left:Document:XR
C1526807|Knee - left X-ray 2 views standing
C1526807|Knee-L XR 2V stand
C1526807|Views 2^standing:Find:Pt:Knee.left:Doc:XR
C1526807|Views 2^standing:Finding:Point in time:Knee.left:Document:XR
C1526812|Ribs-L XR Ant+Lat
C1526812|Ribs - left X-ray anterior and lateral
C1526812|Views anterior & lateral:Find:Pt:Ribs.left:Doc:XR
C1526812|Views anterior & lateral:Finding:Point in time:Ribs.left:Document:XR
C1543378|Lower extremity MRI WO contrast
C1543378|LE MRI WO contr
C1543378|Multisection^WO contrast:Finding:Point in time:Lower extremity:Document:MRI
C1543378|Multisection^WO contrast:Find:Pt:Lower extremity:Doc:MRI
C1524840|LE-R MRI WO contr
C1524840|Lower extremity - right MRI WO contrast
C1524840|Multisection^WO contrast:Finding:Point in time:Lower extremity.right:Document:MRI
C1524840|Multisection^WO contrast:Find:Pt:Lower extremity.right:Doc:MRI
C1524233|Head CT limited WO contrast
C1524233|Head CT Ltd WO contr
C1524233|Multisection limited^WO contrast:Finding:Point in time:Head:Document:Computerized Tomography
C1524233|Multisection limited^WO contrast:Find:Pt:Head:Doc:CT
C1525285|Adrenal gland CT WO contrast
C1525285|Adrenal CT WO contr
C1525285|Multisection^WO contrast:Find:Pt:Abdomen>Adrenal gland:Doc:CT
C1525285|Multisection^WO contrast:Finding:Point in time:Abdomen>Adrenal gland:Document:Computerized Tomography
C1525194|UE joint-L MRI W contr IV
C1525194|Upper extremity joint - left MRI W contrast IV
C1525194|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.joint.left:Document:MRI
C1525194|Multisection^W contrast IV:Find:Pt:Upper extremity.joint.left:Doc:MRI
C1525218|Multisection^WO & W contrast Intravenous:Finding:Point in time:Orbit.right:Document:MRI
C1525218|Orbit - right MRI WO and W contrast IV
C1525218|Orbit-R MRI WO+W contr IV
C1525218|Multisection^WO & W contrast IV:Find:Pt:Orbit.right:Doc:MRI
C1527093|Views:Finding:Point in time:Orbit:Narrative:XR
C1527093|Orbit X-ray
C1527093|Orbit XR
C1527093|Views:Finding:Point in time:Orbit:Document:XR
C1527093|Views:Find:Pt:Orbit:Doc:XR
C1525264|Head CT Bx Str Guid WO contr
C1525264|Guidance for stereotactic biopsy^WO contrast:Finding:Point in time:Head:Document:Computerized Tomography
C1525264|Guidance for stereotactic biopsy^WO contrast:Find:Pt:Head:Doc:CT
C1525264|CT Guidance for stereotactic biopsy of Head-- WO contrast
C1525281|L-spine XR 3V stand
C1525281|Views 3^standing:Finding:Point in time:Spine.lumbar:Document:XR
C1525281|Views 3^standing:Find:Pt:Spine.lumbar:Doc:XR
C1525281|Lumbar spine X-ray 3 views standing
C1524231|Acromioclavicular joint - bilateral X-ray Zanca
C1524231|AC joint-Bl XR Zanca
C1524231|View Zanca:Finding:Point in time:Acromioclavicular joint.bilateral:Document:XR
C1524231|View Zanca:Find:Pt:Acromioclavicular joint.bilateral:Doc:XR
C1525517|Knee-L XR AP+Lat+Sunrise+Tunnel
C1525517|Knee - left X-ray AP and lateral and Sunrise and tunnel
C1525517|Views AP & lateral & Sunrise & tunnel:Find:Pt:Knee.left:Doc:XR
C1525517|Views AP & lateral & Sunrise & tunnel:Finding:Point in time:Knee.left:Document:XR
C1525753|Hrt MRI Cine for Function
C1525753|Heart MRI cine for function
C1525753|Multisection cine for function:Finding:Point in time:Heart:Document:MRI
C1525753|Multisection cine for function:Find:Pt:Heart:Doc:MRI
C1525852|Ankle XR W Stress
C1525852|Ankle X-ray W manual stress
C1525852|Views^W manual stress:Finding:Point in time:Ankle:Document:XR
C1525852|Views^W manual stress:Find:Pt:Ankle:Doc:XR
C1525863|Colon Flr W contr via Colostomy
C1525863|Colon Fluoroscopy W contrast via colostomy
C1525863|Views^W contrast via colostomy:Finding:Point in time:Colon:Document:XR.fluor
C1525863|Views^W contrast via colostomy:Find:Pt:Colon:Doc:XR.fluor
C1525865|Bladder Flr W contr via SP tb
C1525865|Urinary bladder Fluoroscopy W contrast via suprapubic tube
C1525865|Views^W contrast via suprapubic tube:Find:Pt:Urinary bladder:Doc:XR.fluor
C1525865|Views^W contrast via suprapubic tube:Finding:Point in time:Urinary bladder:Document:XR.fluor
C1525867|Wrist - left Fluoroscopy W contrast IS
C1525867|Views^W contrast IS:Find:Pt:Wrist.left:Doc:XR.fluor
C1525867|Views^W contrast Intrasynovial:Finding:Point in time:Wrist.left:Document:XR.fluor
C1525867|Wrist-L Flr W contr IS
C1524138|Coronary graft XRA W contr IA
C1524138|Coronary graft Fluoroscopic angiogram W contrast IA
C1524138|Views^W contrast IA:Find:Pt:Coronary graft:Doc:XR.fluor.angio
C1524138|Views^W contrast Intra-arterial:Finding:Point in time:Coronary graft:Document:XR.fluor.angio
C1525995|Clavicle - right X-ray 2 views
C1525995|Clavicle-R XR 2V
C1525995|Views 2:Find:Pt:Clavicle.right:Doc:XR
C1525995|Views 2:Finding:Point in time:Clavicle.right:Document:XR
C1526016|Foot - right X-ray 3 views standing
C1526016|Ft-R XR 3V stand
C1526016|Views 3^standing:Finding:Point in time:Foot.right:Document:XR
C1526016|Views 3^standing:Find:Pt:Foot.right:Doc:XR
C1526028|Hand-R XR Lat
C1526028|Hand - right X-ray lateral
C1526028|View lateral:Find:Pt:Hand.right:Doc:XR
C1526028|View lateral:Finding:Point in time:Hand.right:Document:XR
C1525902|Wrist-R XR AP+Lat
C1525902|Wrist - right X-ray AP and lateral
C1525902|Views AP & lateral:Find:Pt:Wrist.right:Doc:XR
C1525902|Views AP & lateral:Finding:Point in time:Wrist.right:Document:XR
C1526063|Knee-R XR AP+Lat+Tunnel
C1526063|Knee - right X-ray AP and lateral and tunnel
C1526063|Views AP & lateral & tunnel:Find:Pt:Knee.right:Doc:XR
C1526063|Views AP & lateral & tunnel:Finding:Point in time:Knee.right:Document:XR
C1526077|Knee - right X-ray tunnel
C1526077|Knee-R XR V1 Tunnel
C1526077|View tunnel:Finding:Point in time:Knee.right:Document:XR
C1526077|View tunnel:Find:Pt:Knee.right:Doc:XR
C1526086|Breast - right Mammogram tangential
C1526086|Brst-R Mam Tangential
C1526086|View tangential:Find:Pt:Breast.right:Doc:Mam
C1526086|View tangential:Finding:Point in time:Breast.right:Document:Mam
C1526157|Deprecated View 1 limited:Find:Pt:Sinuses:Nar:XR
C1526157|Deprecated Sinuses XR 1V Ltd
C1526157|Deprecated Sinuses X-ray View
C1526157|View 1 limited:Find:Pt:Sinuses:Nar:XR
C1526157|View 1 limited:Finding:Point in time:Sinuses:Narrative:XR
C1526170|Spine XR Lat Xtable
C1526170|Spine X-ray lateral crosstable
C1526170|View lateral crosstable:Find:Pt:Spine:Doc:XR
C1526170|View lateral crosstable:Finding:Point in time:Spine:Document:XR
C1526178|Tib+Fib XRTomo
C1526178|Tibia and Fibula X-ray tomograph
C1526178|Multisection:Finding:Point in time:Tibia+Fibula:Document:XR.tomo
C1526178|Multisection:Find:Pt:Tibia+Fibula:Doc:XR.tomo
C1526197|Muscle US Bx guid
C1526197|US Guidance for biopsy of Muscle
C1526197|Guidance for biopsy:Finding:Point in time:Muscle:Document:Ultrasound
C1526197|Guidance for biopsy:Find:Pt:Muscle:Doc:US
C1526226|Ribs upper-R XR
C1526226|Ribs upper - right X-ray
C1526226|Views:Find:Pt:Ribs.upper.right:Doc:XR
C1526226|Views:Finding:Point in time:Ribs.upper.right:Document:XR
C1526233|Vertebral artery - right Fluoroscopic angiogram W contrast IA
C1526233|VA-R XRA W contr IA
C1526233|Views^W contrast Intra-arterial:Finding:Point in time:Vertebral artery.right:Document:XR.fluor.angio
C1526233|Views^W contrast IA:Find:Pt:Vertebral artery.right:Doc:XR.fluor.angio
C1525142|Penis ves US
C1525142|Penis vessels US
C1525142|Multisection:Finding:Point in time:Penis vessels:Document:Ultrasound
C1525142|Multisection:Find:Pt:Penis vessels:Doc:US
C1508086|Knee-Bl XR Sunrise 20+40+60 Deg
C1508086|Knee - bilateral X-ray Sunrise 20 and 40 and 60 degrees
C1508086|Views Sunrise 20 & 40 & 60 degrees:Find:Pt:Knee.bilateral:Doc:XR
C1508086|Views Sunrise 20 & 40 & 60 degrees:Finding:Point in time:Knee.bilateral:Document:XR
C1524476|Multisection^W contrast IS:Find:Pt:Shoulder.right:Doc:MRI
C1524476|Shoulder - right MRI W contrast IS
C1524476|Multisection^W contrast Intrasynovial:Finding:Point in time:Shoulder.right:Document:MRI
C1524476|Should-R MRI W contr IS
C1524497|Deprecated Calcaneus - left CT W contrast IV
C1524497|Multisection^W contrast IV:Find:Pt:Calcaneus.left:Doc:CT
C1524497|Deprecated Heel-L CT W contr IV
C1524497|Multisection^W contrast Intravenous:Finding:Point in time:Calcaneus.left:Document:Computerized Tomography
C1524868|Multisection^WO contrast:Find:Pt:Calcaneus:Doc:CT
C1524868|Multisection^WO contrast:Finding:Point in time:Calcaneus:Document:Computerized Tomography
C1524868|Deprecated Heel CT WO contr
C1524868|Deprecated Calcaneus CT WO contrast
C1524894|Knee - right CT WO contrast
C1524894|Knee-R CT WO contr
C1524894|Multisection^WO contrast:Find:Pt:Knee.right:Doc:CT
C1524894|Multisection^WO contrast:Finding:Point in time:Knee.right:Document:Computerized Tomography
C1524909|Spleen MRI WO contr
C1524909|Spleen MRI WO contrast
C1524909|Multisection^WO contrast:Finding:Point in time:Spleen:Document:MRI
C1524909|Multisection^WO contrast:Find:Pt:Spleen:Doc:MRI
C1524916|Lower leg-R CT WO contr
C1524916|Lower leg - right CT WO contrast
C1524916|Multisection^WO contrast:Find:Pt:Lower leg.right:Doc:CT
C1524916|Multisection^WO contrast:Finding:Point in time:Lower leg.right:Document:Computerized Tomography
C1524554|Kidney-L MRI W contr IV
C1524554|Kidney - left MRI W contrast IV
C1524554|Multisection^W contrast IV:Find:Pt:Kidney.left:Doc:MRI
C1524554|Multisection^W contrast Intravenous:Finding:Point in time:Kidney.left:Document:MRI
C1524565|Liver MRI W contr IV
C1524565|Liver MRI W contrast IV
C1524565|Multisection^W contrast IV:Find:Pt:Liver:Doc:MRI
C1524565|Multisection^W contrast Intravenous:Finding:Point in time:Liver:Document:MRI
C1524936|Hand XR 1V
C1524936|Hand X-ray Single view
C1524936|View 1:Find:Pt:Hand:Doc:XR
C1524936|View 1:Finding:Point in time:Hand:Document:XR
C1524201|Ankle XR AP 1V
C1524201|Ankle X-ray AP single view
C1524201|View AP:Find:Pt:Ankle:Doc:XR
C1524201|View AP:Finding:Point in time:Ankle:Document:XR
C1524205|Femur X-ray AP single view
C1524205|Femur XR AP 1V
C1524205|View AP:Find:Pt:Femur:Doc:XR
C1524205|View AP:Finding:Point in time:Femur:Document:XR
C1524299|Fluoroscopy Guidance for biopsy of Liver
C1524299|Liver Flr Bx guid
C1524299|Guidance for biopsy:Finding:Point in time:Liver:Document:XR.fluor
C1524299|Guidance for biopsy:Find:Pt:Liver:Doc:XR.fluor
C1524301|Pancreas Flr Bx guid
C1524301|Fluoroscopy Guidance for biopsy of Pancreas
C1524301|Guidance for biopsy:Finding:Point in time:Pancreas:Document:XR.fluor
C1524301|Guidance for biopsy:Find:Pt:Pancreas:Doc:XR.fluor
C1524971|Hand-L XR PA V1
C1524971|Hand - left X-ray PA
C1524971|View PA:Find:Pt:Hand.left:Doc:XR
C1524971|View PA:Finding:Point in time:Hand.left:Document:XR
C1524334|T-spine CT PC Vertebroplasty guid
C1524334|Guidance for percutaneous vertebroplasty:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C1524334|Guidance for percutaneous vertebroplasty:Find:Pt:Spine.thoracic:Doc:CT
C1524334|CT Guidance for percutaneous vertebroplasty of Thoracic spine
C1524362|Elbow-R CT
C1524362|Elbow - right CT
C1524362|Multisection:Find:Pt:Elbow.right:Doc:CT
C1524362|Multisection:Finding:Point in time:Elbow.right:Document:Computerized Tomography
C1524366|Lower extremity X-ray tomograph
C1524366|LE XRTomo
C1524366|Multisection:Find:Pt:Lower extremity:Doc:XR.tomo
C1524366|Multisection:Finding:Point in time:Lower extremity:Document:XR.tomo
C1524767|Knee - right CT WO and W contrast IV
C1524767|Knee-R CT WO+W contr IV
C1524767|Multisection^WO & W contrast IV:Find:Pt:Knee.right:Doc:CT
C1524767|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee.right:Document:Computerized Tomography
C1524392|Forearm-R CT
C1524392|Forearm - right CT
C1524392|Multisection:Find:Pt:Forearm.right:Doc:CT
C1524392|Multisection:Finding:Point in time:Forearm.right:Document:Computerized Tomography
C1525079|Chest Flr PA+Lat
C1525079|Chest Fluoroscopy PA and lateral
C1525079|Views PA & lateral:Finding:Point in time:Chest:Document:XR.fluor
C1525079|Views PA & lateral:Find:Pt:Chest:Doc:XR.fluor
C1830202|Extr v-Bl DOP Ltd
C1830202|Extremity vein - bilateral US.doppler limited
C1830202|Multisection limited:Find:Pt:Extremity vein.bilateral:Doc:US.doppler
C1830202|Multisection limited:Finding:Point in time:Extremity vein.bilateral:Document:Ultrasound.doppler
C1830213|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.left>Vessels:Document:Computerized Tomography.angio
C1830213|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.left>Vessels:Doc:CT.angio
C1830213|Upper extremity - left Vessels CT angiogram WO and W contrast IV
C1830213|EU ves-L CT.Angio WO+W contr IV
C1830219|Abd CT WO+W red contr vol IV
C1830219|Multisection^WO & W reduced contrast volume IV:Find:Pt:Abdomen:Doc:CT
C1830219|Abdomen CT WO and W reduced contrast volume IV
C1830219|Multisection^WO & W reduced contrast volume Intravenous:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1830226|IAC CT W red contr vol IV
C1830226|Internal auditory canal CT W reduced contrast volume IV
C1830226|Multisection^W reduced contrast volume Intravenous:Finding:Point in time:Internal auditory canal:Document:Computerized Tomography
C1830226|Multisection^W reduced contrast volume IV:Find:Pt:Internal auditory canal:Doc:CT
C1830276|Teeth X-ray bitewing
C1830276|Teeth XR Bitewing
C1830276|Views bitewing:Find:Pt:Teeth:Doc:XR
C1830276|Views bitewing:Finding:Point in time:Teeth:Document:XR
C1830070|Chest Flr GE 4V
C1830070|Chest Fluoroscopy GE 4 views
C1830070|Views GE 4:Find:Pt:Chest:Doc:XR.fluor
C1830070|Views GE 4:Finding:Point in time:Chest:Document:XR.fluor
C1715384|Skull.base CT WO contr
C1715384|Skull.base CT WO contrast
C1715384|Multisection^WO contrast:Find:Pt:Skull.base:Doc:CT
C1715384|Multisection^WO contrast:Finding:Point in time:Skull.base:Document:Computerized Tomography
C1717314|Liver RI W 133Xe IH
C1717314|Views^W Xe-133 IH:Find:Pt:Liver:Doc:Radnuc
C1717314|Views^W Xe-133 Inhalation:Finding:Point in time:Liver:Document:Radnuc
C1717314|Liver Scan W Xe-133 IH
C1715438|Peripheral artery US limited
C1715438|Periph a US Ltd
C1715438|Multisection limited:Find:Pt:Peripheral artery:Doc:US
C1715438|Multisection limited:Finding:Point in time:Peripheral artery:Document:Ultrasound
C1715445|Views 2 limited:Finding:Point in time:Sinuses:Narrative:XR
C1715445|Deprecated Sinuses X-ray 2 views limited
C1715445|Deprecated Sinuses XR V2 Ltd
C1715445|Views 2 limited:Find:Pt:Sinuses:Nar:XR
C1715471|Ankle XR GE 3V
C1715471|Ankle X-ray GE 3 views
C1715471|Views GE 3:Finding:Point in time:Ankle:Document:XR
C1715471|Views GE 3:Find:Pt:Ankle:Doc:XR
C1715488|Kidney CT Ablation guid
C1715488|CT Guidance for ablation of tissue of Kidney
C1715488|Guidance for ablation of tissue:Find:Pt:Kidney:Doc:CT
C1715488|Guidance for ablation of tissue:Finding:Point in time:Kidney:Document:Computerized Tomography
C1645316|Guidance for removal of fluid:Find:Pt:Abdomen:Doc:CT
C1645316|Deprecated CT Guidance for removal of fluid from Abdomen
C1645316|Guidance for removal of fluid:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1645316|Deprecated Abd CT Fld rem guid
C1644148|LE a US Ltd
C1644148|Lower extremity artery US limited
C1644148|Multisection limited:Find:Pt:Lower extremity artery:Doc:US
C1644148|Multisection limited:Finding:Point in time:Lower extremity artery:Document:Ultrasound
C1648951|SPECT WB W Tc99mCEA IV
C1648951|SPECT whole body W Tc-99m Arcitumomab IV
C1648951|Multisection whole body^W Tc-99m Arcitumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1648951|Multisection whole body^W Tc-99m Arcitumomab IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1632340|Ribs-R XR 1V
C1632340|Ribs - right X-ray Single view
C1632340|View 1:Find:Pt:Ribs.right:Doc:XR
C1632340|View 1:Finding:Point in time:Ribs.right:Document:XR
C1645330|Ft.Sesamoids-L XR Axial
C1645330|Foot sesamoid bones - left X-ray axial
C1645330|View axial:Find:Pt:Foot.sesamoid bones.left:Doc:XR
C1645330|View axial:Finding:Point in time:Foot.sesamoid bones.left:Document:XR
C1638464|Views AP^WO & W L-bending:Finding:Point in time:Spine.lumbar:Document:XR
C1638464|Views AP^WO & W L-bending:Find:Pt:Spine.lumbar:Doc:XR
C1638464|L-spine XR AP WO+W L-bending
C1638464|Lumbar spine X-ray AP W and WO left bending
C1714902|Vessel Scan static
C1714902|Views static^W radionuclide IV:Find:Pt:Vessel:Doc:Radnuc
C1714902|Views static^W radionuclide Intravenous:Finding:Point in time:Vessel:Document:Radnuc
C1714902|Vesl RI Static W RNC IV
C1714944|Ankle-L MRI Dyn W contr IV
C1714944|Ankle - left MRI dynamic W contrast IV
C1714944|Multisection dynamic^W contrast IV:Find:Pt:Ankle.left:Doc:MRI
C1714944|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Ankle.left:Document:MRI
C1637281|T+L-spine XR Scoli AP+Lat sitting
C1637281|Views scoliosis AP & lateral^sitting:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1637281|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral sitting
C1637281|Views scoliosis AP & lateral^sitting:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1636069|T+L-spine XR Scoli Lat sitting
C1636069|View scoliosis lateral^sitting:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1636069|Spine Thoracic and Lumbar X-ray scoliosis lateral sitting
C1636069|View scoliosis lateral^sitting:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1623574|Humerus XR in Surg
C1623574|Humerus X-ray during surgery
C1623574|View^during surgery:Finding:Point in time:Humerus:Document:XR
C1623574|View^during surgery:Find:Pt:Humerus:Doc:XR
C1633399|L-spine CT Needle local guid
C1633399|Guidance for needle localization:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1633399|Guidance for needle localization:Find:Pt:Spine.lumbar:Doc:CT
C1633399|CT Guidance for needle localization of Lumbar spine
C1643244|Deprecated Views portable:Finding:Point in time:Tibia.right:Narrative:XR
C1643244|Deprecated Tib-R XR port
C1643244|Views portable:Find:Pt:Tibia.right:Nar:XR
C1643244|Views portable:Finding:Point in time:Tibia.right:Narrative:XR
C1643244|Deprecated Tibia Right X-ray Portable
C1978436|Views & (view AP^standing):Finding:Point in time:Knee.bilateral:Narrative:XR
C1978436|Knee-Bl XR +(AP 1V Stand)
C1978436|Knee - bilateral X-ray and (AP view standing)
C1978436|Views & (view AP^standing):Finding:Point in time:Knee.bilateral:Document:XR
C1978436|Views & (view AP^standing):Find:Pt:Knee.bilateral:Doc:XR
C1954152|Gastric emptying time^post 100 mg sodium octanoate PO:Time:Pt:Exhl gas:Qn:Radnuc
C1954152|Exhaled gas Scan Gastric emptying time post 100 mg sodium octanoate PO
C1954152|ExG RI GE time p 100mg Na octanoate PO
C1954152|Gastric emptying time^post 100 mg sodium octanoate Oral:Time:Point in time:Exhaled gas (breath):Quantitative:Radnuc
C1954304|UE v-Bl US
C1954304|Upper extremity vein - bilateral US
C1954304|Multisection:Finding:Point in time:Upper extremity vein.bilateral:Document:Ultrasound
C1954304|Multisection:Find:Pt:Upper extremity vein.bilateral:Doc:US
C1953041|Spine X-ray oblique
C1953041|Spine XR Obl
C1953041|Views oblique:Finding:Point in time:Spine:Document:XR
C1953041|Views oblique:Find:Pt:Spine:Doc:XR
C1953958|Multisection^WO & W contrast Intrathecal:Finding:Point in time:Spine.lumbar:Document:MRI
C1953958|L-spine MRI WO+W contr IT
C1953958|Multisection^WO & W contrast IT:Find:Pt:Spine.lumbar:Doc:MRI
C1953958|Lumbar spine MRI WO and W contrast IT
C1953962|Clavicle-R MRI W contr IV
C1953962|Clavicle - right MRI W contrast IV
C1953962|Multisection^W contrast IV:Find:Pt:Clavicle.right:Doc:MRI
C1953962|Multisection^W contrast Intravenous:Finding:Point in time:Clavicle.right:Document:MRI
C1954655|Deprecated Scan Guidance for injection of Joint space
C1954655|Deprecated Joint.space RI Inj guid
C1954655|Guidance for injection:Finding:Point in time:Joint.space.To be specified in another part of the message:Narrative:Radnuc
C1954655|Guidance for injection:Find:Pt:Joint.space.XXX:Nar:Radnuc
C2923070|Abdomen MRCP WO contrast
C2923070|Abd MRCP WO contr
C2923070|Guidance for endoscopy^WO contrast:Find:Pt:Liver+Biliary ducts+Pancreas:Doc:MRI
C2923070|Guidance for endoscopy^WO contrast:Finding:Point in time:Liver+Biliary ducts+Pancreas:Document:MRI
C2925712|Hrt MRI W stress+WO+W contr IV
C2925712|Multisection^W stress & WO & W contrast IV:Find:Pt:Heart:Doc:MRI
C2925712|Multisection^W stress & WO & W contrast Intravenous:Finding:Point in time:Heart:Document:MRI
C2925712|Heart MRI W stress and WO and W contrast IV
C2966670|Multisection^W air contrast PR:Find:Pt:Abdomen+Pelvis>Colon+Rectum:Doc:CT
C2966670|Multisection^W air contrast Rectal:Finding:Point in time:Abdomen+Pelvis>Colon+Rectum:Document:Computerized Tomography
C2966670|Colon+Rectum CT W Air contr PR
C2966670|Colon and Rectum CT W air contrast PR
C3533801|Pelvis MRI WO+W contr IV+endorectal coil
C3533801|Multisection^WO & W contrast Intravenous & W endorectal coil:Finding:Point in time:Pelvis:Document:MRI
C3533801|Pelvis MRI WO and W contrast IV and W endorectal coil
C3533801|Multisection^WO & W contrast IV & W endorectal coil:Find:Pt:Pelvis:Doc:MRI
C3262934|Extr-R CT WO contr
C3262934|Extremity - right CT WO contrast
C3262934|Multisection^WO contrast:Finding:Point in time:Extremity.right:Document:Computerized Tomography
C3262934|Multisection^WO contrast:Find:Pt:Extremity.right:Doc:CT
C3263011|Brst implant MRI WO contr
C3263011|Breast implant MRI WO contrast
C3263011|Multisection^WO contrast:Finding:Point in time:Breast implant:Document:MRI
C3263011|Multisection^WO contrast:Find:Pt:Breast implant:Doc:MRI
C3482437|T-spine CT Nerve Block guid
C3482437|Guidance for nerve block:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C3482437|Guidance for nerve block:Find:Pt:Spine.thoracic:Doc:CT
C3482437|CT Guidance for nerve block of Thoracic spine
C3263061|Renal a XRA PTA of ves W contr IA
C3263061|Renal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C3263061|Percutaneous transluminal angioplasty of vessel^W contrast Intra-arterial:Finding:Point in time:Renal artery:Document:XR.fluor.angio
C3263061|Percutaneous transluminal angioplasty of vessel^W contrast IA:Find:Pt:Renal artery:Doc:XR.fluor.angio
C1525318|Hip-Bl XR Lat Xtable
C1525318|Hip - bilateral X-ray lateral crosstable
C1525318|Hip - bilateral X-ray and lateral crosstable
C1525318|Hip-Bl XR +Lat Xtable
C1525318|Views & lateral crosstable:Find:Pt:Hip.bilateral:Doc:XR
C1525318|View lateral crosstable:Find:Pt:Hip.bilateral:Doc:XR
C1525318|Views & lateral crosstable:Finding:Point in time:Hip.bilateral:Document:XR
C1525318|View lateral crosstable:Finding:Point in time:Hip.bilateral:Document:XR
C3262922|Guidance for biopsy.needle:Find:Pt:Chest>Pleura:Doc:CT
C3262922|Guidance for biopsy.needle:Finding:Point in time:Chest>Pleura:Document:Computerized Tomography
C3262922|CT Guidance for needle biopsy of Chest Pleura
C3262922|Chest Pleura CT Bx needle guid
C0942153|Mastoid - right X-ray
C0942153|Mastoid-R XR
C0942153|Views:Finding:Point in time:Mastoid.right:Document:XR
C0942153|Views:Find:Pt:Mastoid.right:Doc:XR
C0942180|Wrist-L XR
C0942180|Wrist - left X-ray
C0942180|Views:Find:Pt:Wrist.left:Doc:XR
C0942180|Views:Finding:Point in time:Wrist.left:Document:XR
C0942202|Thigh-R MRI WO+W contr IV
C0942202|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thigh.right:Document:MRI
C0942202|Thigh - right MRI WO and W contrast IV
C0942202|Multisection^WO & W contrast IV:Find:Pt:Thigh.right:Doc:MRI
C0942208|Should-R MRI WO+W contr IV
C0942208|Multisection^WO & W contrast IV:Find:Pt:Shoulder.right:Doc:MRI
C0942208|Shoulder - right MRI WO and W contrast IV
C0942208|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder.right:Document:MRI
C0942223|Elbow-L MRI
C0942223|Elbow - left MRI
C0942223|Multisection:Find:Pt:Elbow.left:Doc:MRI
C0942223|Multisection:Finding:Point in time:Elbow.left:Document:MRI
C0942278|Knee - left X-ray Merchants
C0942278|Knee-L XR Merchants
C0942278|View Merchants:Find:Pt:Knee.left:Doc:XR
C0942278|View Merchants:Finding:Point in time:Knee.left:Document:XR
C0942295|Cent v-Bl LB Cath plac guid into ves
C0942295|Guidance for placement of large bore catheter into vessel in Central vein - bilateral
C0942295|Guidance for placement of large bore catheter into vessel:Finding:Point in time:Central vein.bilateral:Document
C0942295|Guidance for placement of large bore catheter into vessel:Find:Pt:Central vein.bilateral:Doc
C0942369|Humerus-Bl XR 2V
C0942369|Humerus - bilateral X-ray 2 views
C0942369|Views 2:Finding:Point in time:Humerus.bilateral:Document:XR
C0942369|Views 2:Find:Pt:Humerus.bilateral:Doc:XR
C0882022|Lymph RI W RNC Intra Lymph
C0882022|Lymphatics Scan W radionuclide intra lymphatic
C0882022|Views^W radionuclide intra lymphatic:Find:Pt:Lymphatics:Doc:Radnuc
C0882022|Views^W radionuclide intra lymphatic:Finding:Point in time:Lymphatics:Document:Radnuc
C0882025|Views:Finding:Point in time:Mastoid:Narrative:XR
C0882025|Mastoid XR
C0882025|Mastoid X-ray
C0882025|Views:Finding:Point in time:Mastoid:Document:XR
C0882025|Views:Find:Pt:Mastoid:Doc:XR
C0882030|Nasopharynx+Neck CT W contr IV
C0882030|Nasopharynx and Neck CT W contrast IV
C0882030|Multisection^W contrast Intravenous:Finding:Point in time:Nasopharynx+Neck:Document:Computerized Tomography
C0882030|Multisection^W contrast IV:Find:Pt:Nasopharynx+Neck:Doc:CT
C0882097|Sinuses MRI
C0882097|Multisection:Finding:Point in time:Sinuses:Document:MRI
C0882097|Multisection:Find:Pt:Sinuses:Doc:MRI
C0882117|C-spine MRI W contr IV
C0882117|Multisection^W contrast Intravenous:Finding:Point in time:Spine.cervical:Document:MRI
C0882117|Multisection^W contrast IV:Find:Pt:Spine.cervical:Doc:MRI
C0882117|Cervical spine MRI W contrast IV
C0882217|Unspecified body region Fluoroscopy 30 minutes
C0882217|XXX Flr 30M
C0882217|View:Find:30M:XXX:Doc:XR.fluor
C0882217|View:Finding:30 minutes:To be specified in another part of the message:Document:XR.fluor
C0882218|XXX Flr 45M
C0882218|Unspecified body region Fluoroscopy 45 minutes
C0882218|View:Finding:45 minutes:To be specified in another part of the message:Document:XR.fluor
C0882218|View:Find:45M:XXX:Doc:XR.fluor
C0942099|Should-L Flr W contr IS
C0942099|Views^W contrast IS:Find:Pt:Shoulder.left:Doc:XR.fluor
C0942099|Views^W contrast Intrasynovial:Finding:Point in time:Shoulder.left:Document:XR.fluor
C0942099|Shoulder - left Fluoroscopy W contrast IS
C0881842|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast:Narrative:Mam
C0881842|Mammogram Guidance for core needle percutaneous biopsy of Breast
C0881842|Brst Mam PC Bx CN guid
C0881842|Guidance for percutaneous biopsy.core needle:Find:Pt:Breast:Doc:Mam
C0881842|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast:Document:Mam
C0882193|Views:Finding:Point in time:Wrist:Narrative:XR
C0882193|Wrist XR
C0882193|Wrist X-ray
C0882193|Views:Find:Pt:Wrist:Doc:XR
C0882193|Views:Finding:Point in time:Wrist:Document:XR
C0881874|Chest XR PA+Lat Upr
C0881874|Chest X-ray PA and lateral upright
C0881874|Views PA & lateral upright:Finding:Point in time:Chest:Document:XR
C0881874|Views PA & lateral upright:Find:Pt:Chest:Doc:XR
C0881877|Chest XR R-Obl+L-Obl Upr
C0881877|Chest X-ray right oblique and left oblique upright
C0881877|Views R-oblique & L-oblique upright:Find:Pt:Chest:Doc:XR
C0881877|Views R-oblique & L-oblique upright:Finding:Point in time:Chest:Document:XR
C0881891|Colon Flr W Air+Ba PR
C0881891|Colon Fluoroscopy W air and barium contrast PR
C0881891|Views^W air & barium contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C0881891|Views^W air & barium contrast PR:Find:Pt:Colon:Doc:XR.fluor
C0881892|Colon Fluoroscopy W contrast PR
C0881892|Colon Flr W contr PR
C0881892|Views^W contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C0881892|Views^W contrast PR:Find:Pt:Colon:Doc:XR.fluor
C0881897|Diaphragm US Motion
C0881897|Motion:Find:Pt:Diaphragm:Doc:US
C0881897|Motion:Finding:Point in time:Diaphragm:Document:Ultrasound
C0881915|US Guidance for drainage of Extremity
C0881915|Extr US Drain guid
C0881915|Guidance for drainage:Finding:Point in time:Extremity:Document:Ultrasound
C0881915|Guidance for drainage:Find:Pt:Extremity:Doc:US
C0882530|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thigh:Document:MRI
C0882530|Thigh MRI WO+W contr IV
C0882530|Multisection^WO & W contrast IV:Find:Pt:Thigh:Doc:MRI
C0882530|Thigh MRI WO and W contrast IV
C0882008|Knee X-ray standing
C0882008|Knee XR stand
C0882008|Views^standing:Finding:Point in time:Knee:Document:XR
C0882008|Views^standing:Find:Pt:Knee:Doc:XR
C1114497|Deprecated Kidney - bilateral and Collecting system MRI WO contrast
C1114497|Multisection^WO contrast:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:MRI
C1114497|Multisection^WO contrast:Find:Pt:Kidney.bilateral+Collecting system:Nar:MRI
C1114497|Deprecated KD-Bl+CS MRI WO contr
C1114587|Finger fourth X-ray
C1114587|Finger.4th XR
C1114587|Views:Finding:Point in time:Finger.fourth:Document:XR
C1114587|Views:Find:Pt:Finger.fourth:Doc:XR
C1114614|Fluoroscopy Guidance for injection of Spine Cervical Facet Joint
C1114614|C-Spine facet joint Flr Inj guid
C1114614|Guidance for injection:Find:Pt:Spine.cervical facet joint:Doc:XR.fluor
C1114614|Guidance for injection:Finding:Point in time:Spine.cervical facet joint:Document:XR.fluor
C1114951|Epidural vv XRA W contr IV
C1114951|Epidural veins Fluoroscopic angiogram W contrast IV
C1114951|Views^W contrast Intravenous:Finding:Point in time:Epidural veins:Document:XR.fluor.angio
C1114951|Views^W contrast IV:Find:Pt:Epidural veins:Doc:XR.fluor.angio
C1114623|Head+Neck a XRA W contr IA
C1114623|Head artery and Neck artery Fluoroscopic angiogram W contrast IA
C1114623|Views^W contrast IA:Find:Pt:Head artery+Neck artery:Doc:XR.fluor.angio
C1114623|Views^W contrast Intra-arterial:Finding:Point in time:Head artery+Neck artery:Document:XR.fluor.angio
C1114636|Ab Ao XRA W contr IA
C1114636|Aorta abdominal Fluoroscopic angiogram W contrast IA
C1114636|Views^W contrast IA:Find:Pt:Aorta.abdominal:Doc:XR.fluor.angio
C1114636|Views^W contrast Intra-arterial:Finding:Point in time:Aorta.abdominal:Document:XR.fluor.angio
C1114639|Lymphatics abdominal - bilateral Fluoroscopy W contrast intra lymphatic
C1114639|Lymph Abd-Bl Flr W contr IL
C1114639|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.abdominal.bilateral:Document:XR.fluor
C1114639|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.abdominal.bilateral:Doc:XR.fluor
C1114665|Lower leg MRI WO contrast
C1114665|Lower leg MRI WO contr
C1114665|Multisection^WO contrast:Finding:Point in time:Lower leg:Document:MRI
C1114665|Multisection^WO contrast:Find:Pt:Lower leg:Doc:MRI
C1543452|Ankle-R XR AP+Lat stand
C1543452|Ankle - right X-ray AP and lateral standing
C1543452|Views AP & lateral^standing:Finding:Point in time:Ankle.right:Document:XR
C1543452|Views AP & lateral^standing:Find:Pt:Ankle.right:Doc:XR
C1543460|Knee - right X-ray 2 views and Sunrise and tunnel
C1543460|Knee-R XR 2V+Sunrise+Tunnel
C1543460|Views 2 & Sunrise & tunnel:Finding:Point in time:Knee.right:Document:XR
C1543460|Views 2 & Sunrise & tunnel:Find:Pt:Knee.right:Doc:XR
C1543470|Should-R XR V(w IR+ER)+Ax
C1543470|Shoulder - right X-ray (W internal rotation and W external rotation) and axillary
C1543470|Views (W internal rotation & W external rotation) & axillary:Find:Pt:Shoulder.right:Doc:XR
C1543470|Views (W internal rotation & W external rotation) & axillary:Finding:Point in time:Shoulder.right:Document:XR
C1543872|RI for Inf WB W Ga-67 IV
C1543872|Views for infection whole body^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543872|Views for infection whole body^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543872|Scan for infection whole body W Ga-67 IV
C1543894|Heart Scan first pass
C1543894|Hrt RI FP W RNC IV
C1543894|Views first pass^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543894|Views first pass^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543915|Hrt RI Flow for Shunt Det W RNC IV
C1543915|Heart Scan flow for shunt detection
C1543915|Views flow for shunt detection^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543915|Views flow for shunt detection^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543934|Hrt RI FP+WM+VV+EF W RNC IV
C1543934|Heart Scan first pass and wall motion and ventricular volume and ejection fraction
C1543934|Views first pass & wall motion & ventricular volume & ejection fraction^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543934|Views first pass & wall motion & ventricular volume & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543514|Multisection:Find:Pt:Carotid artery.right:Nar:US.doppler
C1543514|Deprecated Carotid artery Right US.doppler Multisection
C1543514|Deprecated Carot a-R US.doppler
C1543514|Multisection:Finding:Point in time:Carotid artery.right:Narrative:Ultrasound.doppler
C1543181|Ribs XR 2V
C1543181|Ribs X-ray 2 views
C1543181|Views 2:Finding:Point in time:Ribs:Document:XR
C1543181|Views 2:Find:Pt:Ribs:Doc:XR
C1543182|Sacrum+Coccyx XR 3V
C1543182|Sacrum and Coccyx X-ray 3 views
C1543182|Views 3:Finding:Point in time:Sacrum+Coccyx:Document:XR
C1543182|Views 3:Find:Pt:Sacrum+Coccyx:Doc:XR
C1543265|Gastrointestine upper Fluoroscopy W air contrast PO
C1543265|UGI Flr W Air contr PO
C1543265|View^W air contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1543265|View^W air contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1525166|Scapula-R MRI WO contr
C1525166|Scapula - right MRI WO contrast
C1525166|Multisection^WO contrast:Find:Pt:Scapula.right:Doc:MRI
C1525166|Multisection^WO contrast:Finding:Point in time:Scapula.right:Document:MRI
C1543697|Brain RI W Tl-201 IV
C1543697|Brain Scan W Tl-201 IV
C1543697|Views^W Tl-201 IV:Find:Pt:Brain:Doc:Radnuc
C1543697|Views^W Tl-201 Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1543705|Brain vv RI W RNC IV
C1543705|Brain veins Scan
C1543705|Views^W radionuclide IV:Find:Pt:Brain veins:Doc:Radnuc
C1543705|Views^W radionuclide Intravenous:Finding:Point in time:Brain veins:Document:Radnuc
C1543418|L-spine XR AP+Lat stand
C1543418|Views AP & lateral^standing:Find:Pt:Spine.lumbar:Doc:XR
C1543418|Views AP & lateral^standing:Finding:Point in time:Spine.lumbar:Document:XR
C1543418|Lumbar spine X-ray AP and lateral standing
C1525107|Abd vv MRI.Angio
C1525107|Abdominal veins MRI angiogram
C1525107|Multisection:Find:Pt:Abdominal veins:Doc:MRI.angio
C1525107|Multisection:Finding:Point in time:Abdominal veins:Document:MRI.angio
C1525172|LE ves-R MRI.Angio
C1525172|Lower extremity vessels - right MRI angiogram
C1525172|Multisection:Find:Pt:Lower extremity vessels.right:Doc:MRI.angio
C1525172|Multisection:Finding:Point in time:Lower extremity vessels.right:Document:MRI.angio
C1525289|Deprecated Maxillofacial region CT and 3D reconstruction
C1525289|Deprecated Maxillofacial CT +3DR
C1525289|Multisection & 3D reconstruction:Finding:Point in time:Maxillofacial region:Document:Computerized Tomography
C1525289|Multisection & 3D reconstruction:Find:Pt:Maxillofacial region:Doc:CT
C1525192|Temporal bone-R CT W contr IV
C1525192|Temporal bone - right CT W contrast IV
C1525192|Multisection^W contrast IV:Find:Pt:Temporal bone.right:Doc:CT
C1525192|Multisection^W contrast Intravenous:Finding:Point in time:Temporal bone.right:Document:Computerized Tomography
C1525203|Abd ves CT.Angio W contr IV
C1525203|Abdominal vessels CT angiogram W contrast IV
C1525203|Multisection^W contrast IV:Find:Pt:Abdomen>Vessels:Doc:CT.angio
C1525203|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen>Vessels:Document:Computerized Tomography.angio
C1525217|Multisection^WO & W contrast IV:Find:Pt:Orbit.left:Doc:MRI
C1525217|Multisection^WO & W contrast Intravenous:Finding:Point in time:Orbit.left:Document:MRI
C1525217|Orbit - left MRI WO and W contrast IV
C1525217|Orbit-L MRI WO+W contr IV
C1525234|Multisection^WO & W contrast IV:Find:Pt:Upper extremity vessels.left:Doc:MRI.angio
C1525234|Upper extremity vessels - left MRI angiogram WO and W contrast IV
C1525234|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity vessels.left:Document:MRI.angio
C1525234|UE ves-L MRI.Angio WO+W contr IV
C1527092|Orbit MRI WO contrast
C1527092|Orbit MRI WO contr
C1527092|Multisection^WO contrast:Find:Pt:Orbit:Doc:MRI
C1527092|Multisection^WO contrast:Finding:Point in time:Orbit:Document:MRI
C1525265|Pituitary and Sella turcica CT
C1525265|Multisection:Find:Pt:Head>Pituitary+Sella turcica:Doc:CT
C1525265|Multisection:Finding:Point in time:Head>Pituitary+Sella turcica:Document:Computerized Tomography
C1525265|Head Pit+Slla turc CT
C1525502|Hip XR AP+Lat Frog
C1525502|Hip X-ray AP and lateral frog
C1525502|Views AP & lateral frog:Find:Pt:Hip:Doc:XR
C1525502|Views AP & lateral frog:Finding:Point in time:Hip:Document:XR
C1524244|Ankle-Bl XR AP+Lat+Mortise
C1524244|Ankle - bilateral X-ray AP and lateral and Mortise
C1524244|Views AP & lateral & Mortise:Finding:Point in time:Ankle.bilateral:Document:XR
C1524244|Views AP & lateral & Mortise:Find:Pt:Ankle.bilateral:Doc:XR
C1525545|Chest XR PA+Lat+L-Obl
C1525545|Chest X-ray PA and lateral and left oblique
C1525545|Views PA & lateral & L-oblique:Find:Pt:Chest:Doc:XR
C1525545|Views PA & lateral & L-oblique:Finding:Point in time:Chest:Document:XR
C1525555|Knee-L XR Sunrise+Tunnel
C1525555|Knee - left X-ray Sunrise and tunnel
C1525555|Views Sunrise & tunnel:Find:Pt:Knee.left:Doc:XR
C1525555|Views Sunrise & tunnel:Finding:Point in time:Knee.left:Document:XR
C1525567|Hip X-ray portable
C1525567|Hip XR port
C1525567|Views portable:Find:Pt:Hip:Doc:XR
C1525567|Views portable:Finding:Point in time:Hip:Document:XR
C1525600|Lower extremity X-ray standing
C1525600|LE XR stand
C1525600|Views^standing:Finding:Point in time:Lower extremity:Document:XR
C1525600|Views^standing:Find:Pt:Lower extremity:Doc:XR
C1525603|Hip - left X-ray standing
C1525603|Hip-L XR stand
C1525603|View^standing:Find:Pt:Hip.left:Doc:XR
C1525603|View^standing:Finding:Point in time:Hip.left:Document:XR
C1525632|Lower Extremity Joint CT W contrast IS
C1525632|Multisection^W contrast Intrasynovial:Finding:Point in time:Lower extremity.joint:Document:Computerized Tomography
C1525632|Multisection^W contrast IS:Find:Pt:Lower extremity.joint:Doc:CT
C1525632|LE.joint CT W contr IS
C1525654|Temporomandibular joint MRI WO and W contrast IV
C1525654|Multisection^WO & W contrast Intravenous:Finding:Point in time:Temporomandibular joint:Document:MRI
C1525654|TMJ MRI WO+W contr IV
C1525654|Multisection^WO & W contrast IV:Find:Pt:Temporomandibular joint:Doc:MRI
C1525673|Multisection anteversion measurement:Finding:Point in time:Femur+Hip:Document:Computerized Tomography
C1525673|Deprecated Femur and Hip CT anteversion measurement
C1525673|Multisection anteversion measurement:Find:Pt:Femur+Hip:Doc:CT
C1525673|Deprecated Femur+Hip CT Anteversion Meas
C1525719|Carotid artery+Vertebral artery - left Fluoroscopic angiogram W contrast IA
C1525719|Carot a+VA-L XRA W contr IA
C1525719|Views^W contrast IA:Find:Pt:Carotid artery+Vertebral artery.left:Doc:XR.fluor.angio
C1525719|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Vertebral artery.left:Document:XR.fluor.angio
C1525765|Wrist-L CT WO+W contr IV
C1525765|Multisection^WO & W contrast IV:Find:Pt:Wrist.left:Doc:CT
C1525765|Multisection^WO & W contrast Intravenous:Finding:Point in time:Wrist.left:Document:Computerized Tomography
C1525765|Wrist - left CT WO and W contrast IV
C1525810|Lumbar Spine vessels MRI angiogram WO and W contrast IV
C1525810|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.lumbar vessels:Document:MRI.angio
C1525810|L-spine ves MRI.Angio WO+W contr IV
C1525810|Multisection^WO & W contrast IV:Find:Pt:Spine.lumbar vessels:Doc:MRI.angio
C1526127|Toes-R XR AP+Lat
C1526127|Toes - right X-ray AP and lateral
C1526127|Views AP & lateral:Finding:Point in time:Toes.right:Document:XR
C1526127|Views AP & lateral:Find:Pt:Toes.right:Doc:XR
C1526059|Knee - right X-ray 4 views
C1526059|Knee-R XR 4V
C1526059|Views 4:Find:Pt:Knee.right:Doc:XR
C1526059|Views 4:Finding:Point in time:Knee.right:Document:XR
C1526067|Knee - right X-ray lateral
C1526067|Knee-R XR Lat
C1526067|View lateral:Finding:Point in time:Knee.right:Document:XR
C1526067|View lateral:Find:Pt:Knee.right:Doc:XR
C1526099|Shoulder - right X-ray 4 views
C1526099|Should-R XR 4V
C1526099|Views 4:Find:Pt:Shoulder.right:Doc:XR
C1526099|Views 4:Finding:Point in time:Shoulder.right:Document:XR
C1526163|Skull XR Lat+Caldwell+Waters+Towne
C1526163|Skull X-ray lateral and Caldwell and Waters and Towne
C1526163|Views lateral & Caldwell & Waters & Towne:Find:Pt:Skull:Doc:XR
C1526163|Views lateral & Caldwell & Waters & Towne:Finding:Point in time:Skull:Document:XR
C1526166|Skull X-ray tomograph
C1526166|Skull XRTomo
C1526166|Multisection:Find:Pt:Skull:Doc:XR.tomo
C1526166|Multisection:Finding:Point in time:Skull:Document:XR.tomo
C1526230|Sternoclavicular joint - right X-ray
C1526230|SC joint-R XR
C1526230|Views:Find:Pt:Sternoclavicular joint.right:Doc:XR
C1526230|Views:Finding:Point in time:Sternoclavicular joint.right:Document:XR
C1525140|Upper extremity artery - bilateral US
C1525140|UE a-Bl US
C1525140|Multisection:Find:Pt:Upper extremity artery.bilateral:Doc:US
C1525140|Multisection:Finding:Point in time:Upper extremity artery.bilateral:Document:Ultrasound
C1525920|US Guidance for deep aspiration.fine needle of Tissue
C1525920|tiss US Guide for deep FNA
C1525920|Guidance for deep aspiration.fine needle:Finding:Point in time:Tissue:Document:Ultrasound
C1525920|Guidance for deep aspiration.fine needle:Find:Pt:Tissue:Doc:US
C1526329|Wrist - right X-ray scaphoid
C1526329|Wrist-R XR Scaphoid
C1526329|Views scaphoid:Finding:Point in time:Wrist.right:Document:XR
C1526329|Views scaphoid:Find:Pt:Wrist.right:Doc:XR
C1524505|Elbow-R CT W contr IV
C1524505|Elbow - right CT W contrast IV
C1524505|Multisection^W contrast IV:Find:Pt:Elbow.right:Doc:CT
C1524505|Multisection^W contrast Intravenous:Finding:Point in time:Elbow.right:Document:Computerized Tomography
C1524544|Upper arm-L MRI W contr IV
C1524544|Upper arm - left MRI W contrast IV
C1524544|Multisection^W contrast IV:Find:Pt:Upper arm.left:Doc:MRI
C1524544|Multisection^W contrast Intravenous:Finding:Point in time:Upper arm.left:Document:MRI
C1524579|Sacrum CT W contr IV
C1524579|Sacrum CT W contrast IV
C1524579|Multisection^W contrast IV:Find:Pt:Sacrum:Doc:CT
C1524579|Multisection^W contrast Intravenous:Finding:Point in time:Sacrum:Document:Computerized Tomography
C1524935|Ft XR 1V
C1524935|Foot X-ray Single view
C1524935|View 1:Find:Pt:Foot:Doc:XR
C1524935|View 1:Finding:Point in time:Foot:Document:XR
C1524614|Multisection^WO & W contrast IV:Find:Pt:Lower extremity:Doc:CT
C1524614|Lower extremity CT WO and W contrast IV
C1524614|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity:Document:Computerized Tomography
C1524614|LE CT WO+W contr IV
C1524966|Hip-Bl XR Obl 1V
C1524966|Hip - bilateral X-ray oblique single view
C1524966|View oblique:Finding:Point in time:Hip.bilateral:Document:XR
C1524966|View oblique:Find:Pt:Hip.bilateral:Doc:XR
C1524974|Brst-Bl Mam
C1524974|Breast - bilateral Mammogram
C1524974|Views:Finding:Point in time:Breast.bilateral:Document:Mam
C1524974|Views:Find:Pt:Breast.bilateral:Doc:Mam
C1526998|Aorta thoracic MRI
C1526998|TA MRI
C1526998|Multisection:Find:Pt:Aorta.thoracic:Doc:MRI
C1526998|Multisection:Finding:Point in time:Aorta.thoracic:Document:MRI
C1524631|Foot X-ray 3 views
C1524631|Ft XR 3V
C1524631|Views 3:Finding:Point in time:Foot:Document:XR
C1524631|Views 3:Find:Pt:Foot:Doc:XR
C1524649|Elbow - left X-ray 4 views
C1524649|Elbow-L XR 4V
C1524649|Views 4:Find:Pt:Elbow.left:Doc:XR
C1524649|Views 4:Finding:Point in time:Elbow.left:Document:XR
C1524658|L-spine XR 4V
C1524658|Views 4:Finding:Point in time:Spine.lumbar:Document:XR
C1524658|Views 4:Find:Pt:Spine.lumbar:Doc:XR
C1524658|Lumbar spine X-ray 4 views
C1525016|Shoulder - left X-ray 5 views
C1525016|Should-L XR 5V
C1525016|Views 5:Find:Pt:Shoulder.left:Doc:XR
C1525016|Views 5:Finding:Point in time:Shoulder.left:Document:XR
C1524371|Lower extremity - left X-ray tomograph
C1524371|LE-L XRTomo
C1524371|Multisection:Find:Pt:Lower extremity.left:Doc:XR.tomo
C1524371|Multisection:Finding:Point in time:Lower extremity.left:Document:XR.tomo
C1527032|Forearm CT
C1527032|Multisection:Find:Pt:Forearm:Doc:CT
C1527032|Multisection:Finding:Point in time:Forearm:Document:Computerized Tomography
C1524667|Ft CT WO+W contr IV
C1524667|Foot CT WO and W contrast IV
C1524667|Multisection^WO & W contrast Intravenous:Finding:Point in time:Foot:Document:Computerized Tomography
C1524667|Multisection^WO & W contrast IV:Find:Pt:Foot:Doc:CT
C1524735|Forearm - left MRI WO and W contrast IV
C1524735|Forearm-L MRI WO+W contr IV
C1524735|Multisection^WO & W contrast IV:Find:Pt:Forearm.left:Doc:MRI
C1524735|Multisection^WO & W contrast Intravenous:Finding:Point in time:Forearm.left:Document:MRI
C1524740|Hand - left MRI WO and W contrast IV
C1524740|Hand-L MRI WO+W contr IV
C1524740|Multisection^WO & W contrast IV:Find:Pt:Hand.left:Doc:MRI
C1524740|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hand.left:Document:MRI
C1524396|Hand-L CT
C1524396|Hand - left CT
C1524396|Multisection:Find:Pt:Hand.left:Doc:CT
C1524396|Multisection:Finding:Point in time:Hand.left:Document:Computerized Tomography
C1524671|Knee-L XR AP+Lat+Obl
C1524671|Knee - left X-ray AP and lateral and oblique
C1524671|Views AP & lateral & oblique:Finding:Point in time:Knee.left:Document:XR
C1524671|Views AP & lateral & oblique:Find:Pt:Knee.left:Doc:XR
C1830211|Multisection^WO & W contrast Intravenous:Finding:Point in time:Orbit+Face+Neck:Document:MRI
C1830211|Orbit and Face and Neck MRI WO and W contrast IV
C1830211|Orbit+Face+Neck MRI WO+W contr IV
C1830211|Multisection^WO & W contrast IV:Find:Pt:Orbit+Face+Neck:Doc:MRI
C1830258|Colon Flr W Air contr PR
C1830258|Colon Fluoroscopy W air contrast PR
C1830258|Views^W air contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C1830258|Views^W air contrast PR:Find:Pt:Colon:Doc:XR.fluor
C1830259|Multisection whole body:Finding:Point in time:^Patient:Narrative:MRI
C1830259|MRI whole body
C1830259|MRI WB
C1830259|Multisection whole body:Finding:Point in time:^Patient:Document:MRI
C1830259|Multisection whole body:Find:Pt:^Patient:Doc:MRI
C1830087|Chest SPECT Tube plac guid W RNC IV
C1830087|SPECT Guidance for placement of tube in Chest
C1830087|Guidance for placement of tube^W radionuclide Intravenous:Finding:Point in time:Chest:Document:Radnuc.SPECT
C1830087|Guidance for placement of tube^W radionuclide IV:Find:Pt:Chest:Doc:Radnuc.SPECT
C1830088|Cerebral artery US
C1830088|Cerebral a US
C1830088|Multisection:Find:Pt:Cerebral artery:Doc:US
C1830088|Multisection:Finding:Point in time:Cerebral artery:Document:Ultrasound
C1830283|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Head:Document:Computerized Tomography
C1830283|Deprecated Head CT dynamic W contrast IV
C1830283|Deprecated Head CT Dyn W contr IV
C1830283|Multisection dynamic^W contrast IV:Find:Pt:Head:Doc:CT
C1715376|Guidance for aspiration.fine needle:Find:Pt:Chest>Mediastinum:Doc:CT
C1715376|Guidance for aspiration.fine needle:Finding:Point in time:Chest>Mediastinum:Document:Computerized Tomography
C1715376|Chest medias CT FNA Asp
C1715376|CT Guidance for fine needle aspiration of Chest Mediastinum
C1715406|Multisection:Finding:Point in time:To be specified in another part of the message:Narrative:Radnuc.PET
C1715406|Unspecified body region PET
C1715406|XXX PET
C1715406|Multisection:Find:Pt:XXX:Doc:Radnuc.PET
C1715406|Multisection:Finding:Point in time:To be specified in another part of the message:Document:Radnuc.PET
C1715429|Lung US Bx guid
C1715429|US Guidance for biopsy of Lung
C1715429|Guidance for biopsy:Finding:Point in time:Lung:Document:Ultrasound
C1715429|Guidance for biopsy:Find:Pt:Lung:Doc:US
C1715470|Sinuses XR Ltd
C1715470|Sinuses X-ray limited
C1715470|Views limited:Finding:Point in time:Sinuses:Document:XR
C1715470|Views limited:Find:Pt:Sinuses:Doc:XR
C1715479|Fluoroscopy Guidance for fine needle aspiration of Lymph node
C1715479|LN Flr FNA Asp
C1715479|Guidance for aspiration.fine needle:Finding:Point in time:Lymph node:Document:XR.fluor
C1715479|Guidance for aspiration.fine needle:Find:Pt:Lymph node:Doc:XR.fluor
C1715492|Kdny-Bl RI WO+W Tc99mDTPA IV
C1715492|Views^WO & W Tc-99m DTPA IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1715492|Kidney - bilateral Scan WO and W Tc-99m DTPA IV
C1715492|Views^WO & W Tc-99m DTPA Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1714909|Axilla - left MRI
C1714909|Axilla-L MRI
C1714909|Multisection:Finding:Point in time:Axilla.left:Document:MRI
C1714909|Multisection:Find:Pt:Axilla.left:Doc:MRI
C1715027|Liver SPECT Flow W RNC IV
C1715027|Liver SPECT flow
C1715027|Multisection flow^W radionuclide IV:Find:Pt:Liver:Doc:Radnuc.SPECT
C1715027|Multisection flow^W radionuclide Intravenous:Finding:Point in time:Liver:Document:Radnuc.SPECT
C1715032|Deprecated Views^W Tc-99m Mertiatide Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system+Renal vessels:Narrative:Radnuc
C1715032|Views^W Tc-99m Mertiatide IV:Find:Pt:Kidney.bilateral+Collecting system+Renal vessels:Nar:Radnuc
C1715032|Deprecated KD-Bl+CS+Renal ves RI W Tc99m
C1715032|Views^W Tc-99m Mertiatide Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system+Renal vessels:Narrative:Radnuc
C1715032|Deprecated Kidney Bilateral & Collecting System & Renal Vessels Radnuc Views W Tc-99m Mertiatide IV
C1636068|Wrist - bilateral X-ray Single view
C1636068|Wrist-Bl XR 1V
C1636068|View 1:Finding:Point in time:Wrist.bilateral:Document:XR
C1636068|View 1:Find:Pt:Wrist.bilateral:Doc:XR
C1633467|Knee-R XR 30 Deg stand
C1633467|Knee - right X-ray 30 degree standing
C1633467|View 30 degree^standing:Finding:Point in time:Knee.right:Document:XR
C1633467|View 30 degree^standing:Find:Pt:Knee.right:Doc:XR
C1639385|Iliac graft US.doppler
C1639385|Iliac Graft DOP
C1639385|Multisection:Find:Pt:Iliac graft:Doc:US.doppler
C1639385|Multisection:Finding:Point in time:Iliac graft:Document:Ultrasound.doppler
C1639908|Extr ves XRA W contr IV
C1639908|Extremity vessels Fluoroscopic angiogram W contrast IV
C1639908|Views^W contrast IV:Find:Pt:Extremity vessels:Doc:XR.fluor.angio
C1639908|Views^W contrast Intravenous:Finding:Point in time:Extremity vessels:Document:XR.fluor.angio
C1631253|XXX CT Bx guid W contr IV
C1631253|CT Guidance for biopsy of Unspecified body region-- W contrast IV
C1631253|Guidance for biopsy^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1631253|Guidance for biopsy^W contrast IV:Find:Pt:XXX:Doc:CT
C1642594|Elbow - right X-ray limited
C1642594|Elbow-R XR Ltd
C1642594|Views limited:Find:Pt:Elbow.right:Doc:XR
C1642594|Views limited:Finding:Point in time:Elbow.right:Document:XR
C1624131|Bone RI W Tc99mWBC IV
C1624131|Bone Scan W Tc-99m tagged WBC IV
C1624131|Views^W Tc-99m tagged WBC IV:Find:Pt:Bone:Doc:Radnuc
C1624131|Views^W Tc-99m tagged WBC Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1652987|Liver Scan blood pool
C1652987|Liver RI BP W RNC IV
C1652987|Views blood pool^W radionuclide Intravenous:Finding:Point in time:Liver:Document:Radnuc
C1652987|Views blood pool^W radionuclide IV:Find:Pt:Liver:Doc:Radnuc
C1954307|Lower extremity artery US
C1954307|LE a US
C1954307|Multisection:Finding:Point in time:Lower extremity artery:Document:Ultrasound
C1954307|Multisection:Find:Pt:Lower extremity artery:Doc:US
C1954366|Wrist+Hand XR 3V
C1954366|Wrist and Hand X-ray 3 views
C1954366|Views 3:Find:Pt:Wrist+Hand:Doc:XR
C1954366|Views 3:Finding:Point in time:Wrist+Hand:Document:XR
C1954367|Wrist+Hand-Bl XR 3V
C1954367|Wrist - bilateral and Hand - bilateral X-ray 3 views
C1954367|Views 3:Finding:Point in time:Wrist.bilateral+Hand.bilateral:Document:XR
C1954367|Views 3:Find:Pt:Wrist.bilateral+Hand.bilateral:Doc:XR
C2925707|XXX US Ablation guid
C2925707|US Guidance for ablation of tissue of Unspecified body region
C2925707|Guidance for ablation of tissue:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C2925707|Guidance for ablation of tissue:Find:Pt:XXX:Doc:US
C3533807|Multisection^WO & W contrast Intravenous:Finding:Point in time:Toes.right:Document:MRI
C3533807|Toes - right MRI WO and W contrast IV
C3533807|Multisection^WO & W contrast IV:Find:Pt:Toes.right:Doc:MRI
C3533807|Toes-R MRI WO+W contr IV
C3533798|Abdomen MRCP with and without contrast IV
C3533798|Abd MRCP W+WO contr IV
C3533798|Guidance for endoscopy^WO & W contrast IV:Find:Pt:Liver+Biliary ducts+Pancreas:Doc:MRI
C3533798|Guidance for endoscopy^WO & W contrast Intravenous:Finding:Point in time:Liver+Biliary ducts+Pancreas:Document:MRI
C3533796|Small bowel CT W contrast PO and W contrast IV
C3533796|Small bowel CT W contrast PO+IV
C3533796|Multisection^W contrast PO+W contrast IV:Find:Pt:Abdomen+Pelvis>Small bowel:Doc:CT
C3533796|Multisection^W contrast Oral+W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis>Small bowel:Document:Computerized Tomography
C3262943|Guidance for drainage of abscess:Finding:Point in time:Neck:Document:XR.fluor
C3262943|Guidance for drainage of abscess:Find:Pt:Neck:Doc:XR.fluor
C3262943|Fluoroscopy Guidance for drainage of abscess of Neck
C3262943|Neck Flr Abscess drain guid
C3482445|Deprecated T-spine CT Stereo
C3482445|Multisection stereotactic:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C3482445|Multisection stereotactic:Find:Pt:Spine.thoracic:Doc:CT
C3482445|Deprecated Spine Thoracic CT stereotactic
C3261719|Umbilical artery US.doppler
C3261719|Umb a DOP
C3261719|Multisection:Find:Pt:Umbilical artery:Doc:US.doppler
C3261719|Multisection:Finding:Point in time:Umbilical artery:Document:Ultrasound.doppler
C3263087|US Guidance for aspiration of Lymph node
C3263087|LN US Asp guid
C3263087|Guidance for aspiration:Find:Pt:Lymph node:Doc:US
C3263087|Guidance for aspiration:Finding:Point in time:Lymph node:Document:Ultrasound
C3263100|Kidney Transplant US Ltd
C3263100|Kidney transplant US limited
C3263100|Multisection limited:Find:Pt:Kidney transplant:Doc:US
C3263100|Multisection limited:Finding:Point in time:Kidney transplant:Document:Ultrasound
C3263109|Humerus-R XR 1V
C3263109|Humerus - right X-ray Single view
C3263109|View 1:Finding:Point in time:Humerus.right:Document:XR
C3263109|View 1:Find:Pt:Humerus.right:Doc:XR
C3263211|Mesenteric a US
C3263211|Mesenteric artery US
C3263211|Multisection:Find:Pt:Mesenteric artery:Doc:US
C3263211|Multisection:Finding:Point in time:Mesenteric artery:Document:Ultrasound
C3262889|Abd ves XRA W contr IV
C3262889|Abdominal vessels Fluoroscopic angiogram W contrast IV
C3262889|Views^W contrast Intravenous:Finding:Point in time:Abdominal vessels:Document:XR.fluor.angio
C3262889|Views^W contrast IV:Find:Pt:Abdominal vessels:Doc:XR.fluor.angio
C0942156|Optic foramen-R XR
C0942156|Optic foramen - right X-ray
C0942156|Views:Find:Pt:Optic foramen.right:Doc:XR
C0942156|Views:Finding:Point in time:Optic foramen.right:Document:XR
C0945324|LE.joint-Bl MRI
C0945324|Lower extremity joint - bilateral MRI
C0945324|Multisection:Finding:Point in time:Lower extremity.joint.bilateral:Document:MRI
C0945324|Multisection:Find:Pt:Lower extremity.joint.bilateral:Doc:MRI
C0942242|Forearm - bilateral MRI
C0942242|Forearm-Bl MRI
C0942242|Multisection:Find:Pt:Forearm.bilateral:Doc:MRI
C0942242|Multisection:Finding:Point in time:Forearm.bilateral:Document:MRI
C0942302|Mammogram Guidance for needle localization of mass of Breast - bilateral
C0942302|Brst-Bl Mam Needle local mass guid
C0942302|Guidance for needle localization of mass:Finding:Point in time:Breast.bilateral:Document:Mam
C0942302|Guidance for needle localization of mass:Find:Pt:Breast.bilateral:Doc:Mam
C0942319|Cent v-L XRA CC change guid W contr IV
C0942319|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - left-- W contrast IV
C0942319|Guidance for change of central catheter^W contrast Intravenous:Finding:Point in time:Central vein.left:Document:XR.fluor.angio
C0942319|Guidance for change of central catheter^W contrast IV:Find:Pt:Central vein.left:Doc:XR.fluor.angio
C0942325|US Guidance for biopsy of Kidney - bilateral
C0942325|Guidance for biopsy:Finding:Point in time:Kidney.bilateral:Document:Ultrasound
C0942325|Guidance for biopsy:Find:Pt:Kidney.bilateral:Doc:US
C0942325|Kdny-Bl US Bx guid
C0942336|Wrist+Hand-R XR Bone Age
C0942336|Wrist - right and Hand - right X-ray bone age
C0942336|Views bone age:Finding:Point in time:Wrist.right+Hand.right:Document:XR
C0942336|Views bone age:Find:Pt:Wrist.right+Hand.right:Doc:XR
C0882029|Nasopharynx+Neck CT
C0882029|Nasopharynx and Neck CT
C0882029|Multisection:Find:Pt:Nasopharynx+Neck:Doc:CT
C0882029|Multisection:Finding:Point in time:Nasopharynx+Neck:Document:Computerized Tomography
C0882083|Views:Finding:Point in time:Sacroiliac joint:Narrative:XR
C0882083|SIJ XR
C0882083|Sacroiliac Joint X-ray
C0882083|Views:Finding:Point in time:Sacroiliac joint:Document:XR
C0882083|Views:Find:Pt:Sacroiliac joint:Doc:XR
C0882084|SIJ CT Inj guid
C0882084|CT Guidance for injection of Sacroiliac Joint
C0882084|Guidance for injection:Find:Pt:Sacroiliac joint:Doc:CT
C0882084|Guidance for injection:Finding:Point in time:Sacroiliac joint:Document:Computerized Tomography
C0882091|Should XR 3V
C0882091|Shoulder X-ray 3 views
C0882091|Views 3:Find:Pt:Shoulder:Doc:XR
C0882091|Views 3:Finding:Point in time:Shoulder:Document:XR
C0882096|Sinuses CT Ltd
C0882096|Sinuses CT limited
C0882096|Multisection limited:Finding:Point in time:Head>Sinuses:Document:Computerized Tomography
C0882096|Multisection limited:Find:Pt:Head>Sinuses:Doc:CT
C0882166|Thyroid RI W I-131 IV
C0882166|Thyroid Scan W I-131 IV
C0882166|Views^W I-131 Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C0882166|Views^W I-131 IV:Find:Pt:Thyroid:Doc:Radnuc
C0882209|XXX MRI Add'l seq
C0882209|Unspecified body region MRI additional sequence
C0882209|Multisection additional sequence:Find:Pt:XXX:Doc:MRI
C0882209|Multisection additional sequence:Finding:Point in time:To be specified in another part of the message:Document:MRI
C0947253|Knee-L RI W RNC IV
C0947253|Knee - left Scan
C0947253|Views^W radionuclide Intravenous:Finding:Point in time:Knee.left:Document:Radnuc
C0947253|Views^W radionuclide IV:Find:Pt:Knee.left:Doc:Radnuc
C0882515|Views:Finding:Point in time:Acromioclavicular joint:Narrative:XR
C0882515|Acromioclavicular Joint X-ray
C0882515|AC joint XR
C0882515|Views:Finding:Point in time:Acromioclavicular joint:Document:XR
C0882515|Views:Find:Pt:Acromioclavicular joint:Doc:XR
C0881884|Chest ves MRI.Angio W contr IV
C0881884|Chest vessels MRI angiogram W contrast IV
C0881884|Multisection^W contrast IV:Find:Pt:Chest vessels:Doc:MRI.angio
C0881884|Multisection^W contrast Intravenous:Finding:Point in time:Chest vessels:Document:MRI.angio
C0881978|Views 3 serial^WO & W contrast IV:Find:Pt:Kidney.bilateral:Doc:XR
C0881978|Kdny-Bl XR 3V Serial WO+W contr IV
C0881978|Views 3 serial^WO & W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:XR
C0881978|Kidney - bilateral X-ray 3 views serial WO and W contrast IV
C0882000|Views^W contrast Intrasynovial:Finding:Point in time:Knee:Document:XR.fluor
C0882000|Knee Flr W contr IS
C0882000|Knee Fluoroscopy W contrast IS
C0882000|Views^W contrast IS:Find:Pt:Knee:Doc:XR.fluor
C0882016|Liver+Spleen RI W Tc99mCa colloid IV
C0882016|Liver and Spleen Scan W Tc-99m calcium colloid IV
C0882016|Views^W Tc-99m calcium colloid IV:Find:Pt:Liver+Spleen:Doc:Radnuc
C0882016|Views^W Tc-99m calcium colloid Intravenous:Finding:Point in time:Liver+Spleen:Document:Radnuc
C1114492|Multisection^WO & W contrast Intravenous:Finding:Point in time:Liver:Document:MRI
C1114492|Liver MRI WO+W contr IV
C1114492|Multisection^WO & W contrast IV:Find:Pt:Liver:Doc:MRI
C1114492|Liver MRI WO and W contrast IV
C1114551|Chest XR L-Lat port
C1114551|Chest X-ray left lateral portable
C1114551|View L-lateral portable:Finding:Point in time:Chest:Document:XR
C1114551|View L-lateral portable:Find:Pt:Chest:Doc:XR
C1114638|Lymphatics abdominal Fluoroscopy W contrast intra lymphatic
C1114638|Lymph Abd Flr W contr IL
C1114638|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.abdominal:Document:XR.fluor
C1114638|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.abdominal:Doc:XR.fluor
C1114683|Tibioperoneal ves MRI.Angio
C1114683|Tibioperoneal vessels MRI angiogram
C1114683|Multisection:Find:Pt:Tibioperoneal vessels:Doc:MRI.angio
C1114683|Multisection:Finding:Point in time:Tibioperoneal vessels:Document:MRI.angio
C1114443|Pelvis CT WO contr
C1114443|Pelvis CT WO contrast
C1114443|Multisection^WO contrast:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1114443|Multisection^WO contrast:Find:Pt:Pelvis:Doc:CT
C1114461|UGI Flr +AP W contr PO
C1114461|Gastrointestine upper Fluoroscopy and AP W contrast PO
C1114461|Views & AP^W contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1114461|Views & AP^W contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1543421|Should-Bl XR AP(w IR+ER)+Ax
C1543421|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation) and axillary
C1543421|Views AP (W internal rotation & W external rotation) & axillary:Finding:Point in time:Shoulder.bilateral:Document:XR
C1543421|Views AP (W internal rotation & W external rotation) & axillary:Find:Pt:Shoulder.bilateral:Doc:XR
C1543427|Deprecated Chest X-ray PA & oblique W nipple markers
C1543427|Deprecated Chest XR PA+Obl W nipple mark
C1543427|Views PA & oblique^W nipple markers:Find:Pt:Chest:Nar:XR
C1543427|Views PA & oblique^W nipple markers:Finding:Point in time:Chest:Narrative:XR
C1543737|SPECT for Abscess W Ga-67 IV
C1543737|Multisection for abscess^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543737|Multisection for abscess^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1765325|Liver RI W Tc99mRBC IV
C1765325|Liver Scan W Tc-99m tagged RBC IV
C1765325|Views^W Tc-99m tagged RBC IV:Find:Pt:Liver:Doc:Radnuc
C1765325|Views^W Tc-99m tagged RBC Intravenous:Finding:Point in time:Liver:Document:Radnuc
C1543744|Liver SPECT
C1543744|Liver SPECT W RNC IV
C1543744|Multisection^W radionuclide IV:Find:Pt:Liver:Doc:Radnuc.SPECT
C1543744|Multisection^W radionuclide Intravenous:Finding:Point in time:Liver:Document:Radnuc.SPECT
C1543754|Hrt RI PF W DBM+Tc99mMIBI IV
C1543754|Heart Scan perfusion W dobutamine and W Tc-99m Sestamibi IV
C1543754|Views perfusion^W dobutamine & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543754|Views perfusion^W dobutamine & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543778|Hrt RI PF Rest+stress+W RNC IV
C1543778|Heart Scan perfusion at rest and W stress and W radionuclide IV
C1543778|Views perfusion^at rest & W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543778|Views perfusion^at rest & W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543790|Abd RI W In-111 Satmb IV
C1543790|Abdomen Scan W In-111 Satumomab IV
C1543790|Views^W In-111 Satumomab Intravenous:Finding:Point in time:Abdomen:Document:Radnuc
C1543790|Views^W In-111 Satumomab IV:Find:Pt:Abdomen:Doc:Radnuc
C1543876|RI W In-111 Satmb IV
C1543876|Scan W In-111 Satumomab IV
C1543876|Views^W In-111 Satumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543876|Views^W In-111 Satumomab IV:Find:Pt:^Patient:Doc:Radnuc
C1543902|Bone RI 2 Phase W RNC IV
C1543902|Bone Scan 2 views phase
C1543902|Views 2 phase^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543902|Views 2 phase^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543921|Salivary gland RI Flow W RNC IV
C1543921|Salivary gland Scan flow
C1543921|Views flow^W radionuclide Intravenous:Finding:Point in time:Salivary gland:Document:Radnuc
C1543921|Views flow^W radionuclide IV:Find:Pt:Salivary gland:Doc:Radnuc
C1543960|Lung RI V+EQ W RNC IH SB
C1543960|Views ventilation & equilibrium^W radionuclide IH single breath:Find:Pt:Lung:Doc:Radnuc
C1543960|Lung Scan ventilation and equilibrium W radionuclide IH single breath
C1543960|Views ventilation & equilibrium^W radionuclide Inhalation single breath:Finding:Point in time:Lung:Document:Radnuc
C1543967|Vein RI for Thrombosis W RNC IV
C1543967|Vein Scan for thrombosis
C1543967|Views for thrombosis^W radionuclide Intravenous:Finding:Point in time:Vein:Document:Radnuc
C1543967|Views for thrombosis^W radionuclide IV:Find:Pt:Vein:Doc:Radnuc
C1543502|Renal vessels US.doppler
C1543502|Renal ves DOP
C1543502|Multisection:Finding:Point in time:Renal vessels:Document:Ultrasound.doppler
C1543502|Multisection:Find:Pt:Renal vessels:Doc:US.doppler
C1543170|T+L-spine XR AP 1V
C1543170|Spine Thoracic and Lumbar X-ray AP single view
C1543170|View AP:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1543170|View AP:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1543189|Ft XR AP+Lat stand
C1543189|Foot X-ray AP and lateral standing
C1543189|Views AP & lateral^standing:Find:Pt:Foot:Doc:XR
C1543189|Views AP & lateral^standing:Finding:Point in time:Foot:Document:XR
C1543591|Shoulder X-ray Stryker Notch
C1543591|Should XR Stryker Notch
C1543591|View Stryker Notch:Find:Pt:Shoulder:Doc:XR
C1543591|View Stryker Notch:Finding:Point in time:Shoulder:Document:XR
C1543595|Skull XR PA+R-Lat+L-Lat+Towne
C1543595|Skull X-ray PA and right lateral and left lateral and Towne
C1543595|Views PA & R-lateral & L-lateral & Towne:Find:Pt:Skull:Doc:XR
C1543595|Views PA & R-lateral & L-lateral & Towne:Finding:Point in time:Skull:Document:XR
C1543718|Heart SPECT for infarct
C1543718|Hrt SPECT for Infarct W RNC IV
C1543718|Multisection for infarct^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543718|Multisection for infarct^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543728|Hrt RI W Stress+W 201 TH IV
C1543728|Heart Scan W stress and W 201 Th IV
C1543728|Views^W stress & W 201 TH IV:Find:Pt:Heart:Doc:Radnuc
C1543728|Views^W stress & W 201 TH Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1526782|Parotid gland - right Fluoroscopy W contrast intra salivary duct
C1526782|Parotid gland-R Flr W contr intra SD
C1526782|Views^W contrast intra salivary duct:Finding:Point in time:Parotid gland.right:Document:XR.fluor
C1526782|Views^W contrast intra salivary duct:Find:Pt:Parotid gland.right:Doc:XR.fluor
C1524845|Femur CT WO contr
C1524845|Femur CT WO contrast
C1524845|Multisection^WO contrast:Finding:Point in time:Femur:Document:Computerized Tomography
C1524845|Multisection^WO contrast:Find:Pt:Femur:Doc:CT
C1525178|Orbit vessels MRI angiogram
C1525178|Orbit ves MRI.Angio
C1525178|Multisection:Finding:Point in time:Orbit vessels:Document:MRI.angio
C1525178|Multisection:Find:Pt:Orbit vessels:Doc:MRI.angio
C1524240|L-spine MRI Ltd WO contr
C1524240|Multisection limited^WO contrast:Find:Pt:Spine.lumbar:Doc:MRI
C1524240|Multisection limited^WO contrast:Finding:Point in time:Spine.lumbar:Document:MRI
C1524240|Lumbar spine MRI limited WO contrast
C1524242|Kidney MRI W contr IV
C1524242|Kidney MRI W contrast IV
C1524242|Multisection^W contrast IV:Find:Pt:Kidney:Doc:MRI
C1524242|Multisection^W contrast Intravenous:Finding:Point in time:Kidney:Document:MRI
C1525189|Abd+Pelvis CT W contr IV
C1525189|Abdomen and Pelvis CT W contrast IV
C1525189|Multisection^W contrast IV:Find:Pt:Abdomen+Pelvis:Doc:CT
C1525189|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis:Document:Computerized Tomography
C1525228|Multisection^WO & W contrast IV:Find:Pt:Pelvis veins:Doc:MRI.angio
C1525228|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pelvis veins:Document:MRI.angio
C1525228|Pelvis veins MRI angiogram WO and W contrast IV
C1525228|Pelvis vv MRI.Angio WO+W contr IV
C1525334|Knee - left X-ray lateral standing
C1525334|Knee-L XR Lat stand
C1525334|View lateral^standing:Find:Pt:Knee.left:Doc:XR
C1525334|View lateral^standing:Finding:Point in time:Knee.left:Document:XR
C1525335|L-spine XR Lat stand
C1525335|View lateral^standing:Find:Pt:Spine.lumbar:Doc:XR
C1525335|View lateral^standing:Finding:Point in time:Spine.lumbar:Document:XR
C1525335|Lumbar spine X-ray lateral standing
C1525345|Views ski jump:Finding:Point in time:Calcaneus.left:Document:XR
C1525345|Views ski jump:Find:Pt:Calcaneus.left:Doc:XR
C1525345|Deprecated Calcaneus - left X-ray ski jump
C1525345|Deprecated Heel-L XR Ski Jump
C1524223|Shoulder - left X-ray Velpeau axillary
C1524223|Should-L XR Velpeau Ax
C1524223|View Velpeau axillary:Find:Pt:Shoulder.left:Doc:XR
C1524223|View Velpeau axillary:Finding:Point in time:Shoulder.left:Document:XR
C1525479|Foot - bilateral X-ray 2 views standing
C1525479|Ft-Bl XR 2V stand
C1525479|Views 2^standing:Find:Pt:Foot.bilateral:Doc:XR
C1525479|Views 2^standing:Finding:Point in time:Foot.bilateral:Document:XR
C1525484|L-spine XR 5V stand
C1525484|Views 5^standing:Finding:Point in time:Spine.lumbar:Document:XR
C1525484|Views 5^standing:Find:Pt:Spine.lumbar:Doc:XR
C1525484|Lumbar spine X-ray 5 views standing
C1525490|C-spine XR AP+Lat+Odont port
C1525490|Views AP & lateral & odontoid portable:Find:Pt:Spine.cervical:Doc:XR
C1525490|Views AP & lateral & odontoid portable:Finding:Point in time:Spine.cervical:Document:XR
C1525490|Cervical spine X-ray AP and lateral and odontoid portable
C1525500|Pelvis+Hip XR AP+Lat Xtable
C1525500|Pelvis and Hip X-ray AP and lateral crosstable
C1525500|Views AP & lateral crosstable:Finding:Point in time:Pelvis+Hip:Document:XR
C1525500|Views AP & lateral crosstable:Find:Pt:Pelvis+Hip:Doc:XR
C1114579|Views portable:Finding:Point in time:Spine.lumbar:Narrative:XR
C1114579|L-spine XR port
C1114579|Views portable:Finding:Point in time:Spine.lumbar:Document:XR
C1114579|Views portable:Find:Pt:Spine.lumbar:Doc:XR
C1114579|Lumbar spine X-ray portable
C1525592|LE vv-L XRA W contr IV
C1525592|Lower extremity veins - left Fluoroscopic angiogram W contrast IV
C1525592|Views^W contrast IV:Find:Pt:Lower extremity veins.left:Doc:XR.fluor.angio
C1525592|Views^W contrast Intravenous:Finding:Point in time:Lower extremity veins.left:Document:XR.fluor.angio
C1525614|Brain.temporal MRI
C1525614|Multisection:Finding:Point in time:Brain.temporal:Document:MRI
C1525614|Multisection:Find:Pt:Brain.temporal:Doc:MRI
C1525625|TMJ-L MRI
C1525625|Temporomandibular joint - left MRI
C1525625|Multisection:Find:Pt:Temporomandibular joint.left:Doc:MRI
C1525625|Multisection:Finding:Point in time:Temporomandibular joint.left:Document:MRI
C1525669|TMJ-R MRI WO contr
C1525669|Temporomandibular joint - right MRI WO contrast
C1525669|Multisection^WO contrast:Find:Pt:Temporomandibular joint.right:Doc:MRI
C1525669|Multisection^WO contrast:Finding:Point in time:Temporomandibular joint.right:Document:MRI
C1525699|C+T-spine XR AP+Lat
C1525699|Spine Cervical and Spine Thoracic X-ray AP and lateral
C1525699|Views AP & lateral:Finding:Point in time:Spine.cervical+Spine.thoracic:Document:XR
C1525699|Views AP & lateral:Find:Pt:Spine.cervical+Spine.thoracic:Doc:XR
C1525706|Ac arch+Brach a XRA W contr IA
C1525706|Aortic arch and Brachial artery Fluoroscopic angiogram W contrast IA
C1525706|Views^W contrast IA:Find:Pt:Aortic arch+Brachial artery:Doc:XR.fluor.angio
C1525706|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Brachial artery:Document:XR.fluor.angio
C1525723|Gastric artery Fluoroscopic angiogram W contrast IA
C1525723|Gastric a XRA W contr IA
C1525723|Views^W contrast Intra-arterial:Finding:Point in time:Gastric artery:Document:XR.fluor.angio
C1525723|Views^W contrast IA:Find:Pt:Gastric artery:Doc:XR.fluor.angio
C1525737|Extr vv-L XRA W contr IV
C1525737|Extremity veins - left Fluoroscopic angiogram W contrast IV
C1525737|Views^W contrast Intravenous:Finding:Point in time:Extremity veins.left:Document:XR.fluor.angio
C1525737|Views^W contrast IV:Find:Pt:Extremity veins.left:Doc:XR.fluor.angio
C1525790|Ankle XR Broden W Stress
C1525790|Ankle X-ray Broden W manual stress
C1525790|Views Broden^W manual stress:Find:Pt:Ankle:Doc:XR
C1525790|Views Broden^W manual stress:Finding:Point in time:Ankle:Document:XR
C1524140|Lymph Abd+Pelvic Flr W contr IL
C1524140|Lymphatics abdominal and Lymphatics pelvic Fluoroscopy W contrast intra lymphatic
C1524140|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.abdominal+Lymphatics.pelvic:Doc:XR.fluor
C1524140|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.abdominal+Lymphatics.pelvic:Document:XR.fluor
C1525887|Ribs-L+Chest XR Lat+PA Chst
C1525887|Ribs - left and Chest X-ray lateral and PA chest
C1525887|Views lateral & PA chest:Finding:Point in time:Ribs.left+Chest:Document:XR
C1525887|Views lateral & PA chest:Find:Pt:Ribs.left+Chest:Doc:XR
C1525826|Finger.3rd-Bl XR
C1525826|Finger third - bilateral X-ray
C1525826|Views:Find:Pt:Finger.third.bilateral:Doc:XR
C1525826|Views:Finding:Point in time:Finger.third.bilateral:Document:XR
C1525980|Acetabulum - right X-ray 2 views
C1525980|Acetabulum-R XR 2V
C1525980|Views 2:Finding:Point in time:Acetabulum.right:Document:XR
C1525980|Views 2:Find:Pt:Acetabulum.right:Doc:XR
C1526008|Femur-R XR AP+Lat
C1526008|Femur - right X-ray AP and lateral
C1526008|Views AP & lateral:Find:Pt:Femur.right:Doc:XR
C1526008|Views AP & lateral:Finding:Point in time:Femur.right:Document:XR
C1526112|Should-R XR Ax+Y
C1526112|Shoulder - right X-ray axillary and Y
C1526112|Views axillary & Y:Finding:Point in time:Shoulder.right:Document:XR
C1526112|Views axillary & Y:Find:Pt:Shoulder.right:Doc:XR
C1525898|Wrist-R XR 4V
C1525898|Wrist - right X-ray 4 views
C1525898|Views 4:Find:Pt:Wrist.right:Doc:XR
C1525898|Views 4:Finding:Point in time:Wrist.right:Document:XR
C1525898|VIEWS 4:FINDING:POINT IN TIME:WRIST.RIGHT:NARRATIVE:XR
C1526061|Knee-R XR AP+Lat
C1526061|Knee - right X-ray AP and lateral
C1526061|Views AP & lateral:Finding:Point in time:Knee.right:Document:XR
C1526061|Views AP & lateral:Find:Pt:Knee.right:Doc:XR
C1525125|Breast - right Mammogram roll
C1525125|Brst-R Mam Roll
C1525125|Views roll:Find:Pt:Breast.right:Doc:Mam
C1525125|Views roll:Finding:Point in time:Breast.right:Document:Mam
C1526150|Sinuses XR Lat
C1526150|Sinuses X-ray lateral
C1526150|View lateral:Find:Pt:Sinuses:Doc:XR
C1526150|View lateral:Finding:Point in time:Sinuses:Document:XR
C1524275|Subclavian artery Fluoroscopic angiogram W contrast IA
C1524275|Subclavian a XRA W contr IA
C1524275|Views^W contrast IA:Find:Pt:Subclavian artery:Doc:XR.fluor.angio
C1524275|Views^W contrast Intra-arterial:Finding:Point in time:Subclavian artery:Document:XR.fluor.angio
C1524278|Thumb XR AP+Lat
C1524278|Thumb X-ray AP and lateral
C1524278|Views AP & lateral:Find:Pt:Thumb:Doc:XR
C1524278|Views AP & lateral:Finding:Point in time:Thumb:Document:XR
C1526177|Tib+Fib XR AP 1V
C1526177|Tibia and Fibula X-ray AP single view
C1526177|View AP:Finding:Point in time:Tibia+Fibula:Document:XR
C1526177|View AP:Find:Pt:Tibia+Fibula:Doc:XR
C1526190|T-spine XR Lat stand
C1526190|View lateral^standing:Find:Pt:Spine.thoracic:Doc:XR
C1526190|View lateral^standing:Finding:Point in time:Spine.thoracic:Document:XR
C1526190|Thoracic spine X-ray lateral standing
C1526231|Subclavian a-R XRA W contr IA
C1526231|Subclavian artery - right Fluoroscopic angiogram W contrast IA
C1526231|Views^W contrast IA:Find:Pt:Subclavian artery.right:Doc:XR.fluor.angio
C1526231|Views^W contrast Intra-arterial:Finding:Point in time:Subclavian artery.right:Document:XR.fluor.angio
C1526292|C+T+L+Sacrum MRI W contr IV
C1526292|Spine Cervical and Spine Thoracic and Spine Lumbar and Sacrum MRI W contrast IV
C1526292|Multisection^W contrast Intravenous:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar+Sacrum:Document:MRI
C1526292|Multisection^W contrast IV:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar+Sacrum:Doc:MRI
C1525914|Iliac ves-Bl US
C1525914|Iliac vessels - bilateral US
C1525914|Multisection:Finding:Point in time:Iliac vessels.bilateral:Document:Ultrasound
C1525914|Multisection:Find:Pt:Iliac vessels.bilateral:Doc:US
C1526341|Toe 2nd-R XR
C1526341|Toe second - right X-ray
C1526341|Views:Finding:Point in time:Toe.second.right:Document:XR
C1526341|Views:Find:Pt:Toe.second.right:Doc:XR
C1526348|Wrist XR 4V
C1526348|Wrist X-ray 4 views
C1526348|Views 4:Find:Pt:Wrist:Doc:XR
C1526348|Views 4:Finding:Point in time:Wrist:Document:XR
C1524892|Knee - left CT WO contrast
C1524892|Knee-L CT WO contr
C1524892|Multisection^WO contrast:Finding:Point in time:Knee.left:Document:Computerized Tomography
C1524892|Multisection^WO contrast:Find:Pt:Knee.left:Doc:CT
C1524513|UE-L CT W contr IV
C1524513|Upper extremity - left CT W contrast IV
C1524513|Multisection^W contrast IV:Find:Pt:Upper extremity.left:Doc:CT
C1524513|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.left:Document:Computerized Tomography
C1524520|Femur-R CT W contr IV
C1524520|Femur - right CT W contrast IV
C1524520|Multisection^W contrast Intravenous:Finding:Point in time:Femur.right:Document:Computerized Tomography
C1524520|Multisection^W contrast IV:Find:Pt:Femur.right:Doc:CT
C1524530|Forearm MRI W contr IV
C1524530|Forearm MRI W contrast IV
C1524530|Multisection^W contrast Intravenous:Finding:Point in time:Forearm:Document:MRI
C1524530|Multisection^W contrast IV:Find:Pt:Forearm:Doc:MRI
C1524537|Hand-L CT W contr IV
C1524537|Hand - left CT W contrast IV
C1524537|Multisection^W contrast IV:Find:Pt:Hand.left:Doc:CT
C1524537|Multisection^W contrast Intravenous:Finding:Point in time:Hand.left:Document:Computerized Tomography
C1524164|Deprecated Heel CT W contr IV
C1524164|Multisection^W contrast IV:Find:Pt:Calcaneus:Doc:CT
C1524164|Deprecated Calcaneus CT W contrast IV
C1524164|Multisection^W contrast Intravenous:Finding:Point in time:Calcaneus:Document:Computerized Tomography
C1524920|Renal v MRI.Angio WO contr
C1524920|Renal vein MRI angiogram WO contrast
C1524920|Multisection^WO contrast:Find:Pt:Renal vein:Doc:MRI.angio
C1524920|Multisection^WO contrast:Finding:Point in time:Renal vein:Document:MRI.angio
C1524578|Prostate MRI W contr IV
C1524578|Prostate MRI W contrast IV
C1524578|Multisection^W contrast Intravenous:Finding:Point in time:Prostate:Document:MRI
C1524578|Multisection^W contrast IV:Find:Pt:Prostate:Doc:MRI
C1524215|Knee-Bl XR AP 1V
C1524215|Knee - bilateral X-ray AP single view
C1524215|View AP:Finding:Point in time:Knee.bilateral:Document:XR
C1524215|View AP:Find:Pt:Knee.bilateral:Doc:XR
C1524949|Hand - left X-ray lateral
C1524949|Hand-L XR Lat
C1524949|View lateral:Find:Pt:Hand.left:Doc:XR
C1524949|View lateral:Finding:Point in time:Hand.left:Document:XR
C1524322|Chest CT Drain guid W contr IV
C1524322|CT Guidance for drainage of Chest-- W contrast IV
C1524322|Guidance for drainage^W contrast IV:Find:Pt:Chest:Doc:CT
C1524322|Guidance for drainage^W contrast Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C1524356|Multisection:Finding:Point in time:Clavicle:Narrative:MRI
C1524356|Clavicle MRI
C1524356|Multisection:Find:Pt:Clavicle:Doc:MRI
C1524356|Multisection:Finding:Point in time:Clavicle:Document:MRI
C1524359|Elbow - bilateral CT
C1524359|Elbow-Bl CT
C1524359|Multisection:Find:Pt:Elbow.bilateral:Doc:CT
C1524359|Multisection:Finding:Point in time:Elbow.bilateral:Document:Computerized Tomography
C1524360|Elbow - left CT
C1524360|Elbow-L CT
C1524360|Multisection:Find:Pt:Elbow.left:Doc:CT
C1524360|Multisection:Finding:Point in time:Elbow.left:Document:Computerized Tomography
C1524373|Lower extremity - right CT
C1524373|LE-R CT
C1524373|Multisection:Finding:Point in time:Lower extremity.right:Document:Computerized Tomography
C1524373|Multisection:Find:Pt:Lower extremity.right:Doc:CT
C1524375|Upper extremity CT
C1524375|UE CT
C1524375|Multisection:Find:Pt:Upper extremity:Doc:CT
C1524375|Multisection:Finding:Point in time:Upper extremity:Document:Computerized Tomography
C1524384|Fetal MRI
C1524384|Fet MRI
C1524384|Multisection:Find:Pt:^Fetus:Doc:MRI
C1524384|Multisection:Finding:Point in time:^Fetus:Document:MRI
C1524387|Foot - left CT
C1524387|Ft-L CT
C1524387|Multisection:Find:Pt:Foot.left:Doc:CT
C1524387|Multisection:Finding:Point in time:Foot.left:Document:Computerized Tomography
C1524666|Multisection^WO & W contrast IV:Find:Pt:Femur.right:Doc:CT
C1524666|Femur - right CT WO and W contrast IV
C1524666|Femur-R CT WO+W contr IV
C1524666|Multisection^WO & W contrast Intravenous:Finding:Point in time:Femur.right:Document:Computerized Tomography
C1524757|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.joint:Doc:MRI
C1524757|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.joint:Document:MRI
C1524757|Lower Extremity Joint MRI WO and W contrast IV
C1524757|LE.joint MRI WO+W contr IV
C1525043|Hip-L XR AP+Lat
C1525043|Hip - left X-ray AP and lateral
C1525043|Views AP & lateral:Finding:Point in time:Hip.left:Document:XR
C1525043|Views AP & lateral:Find:Pt:Hip.left:Doc:XR
C1525091|Fem a+Popliteal a XRA Angpsty W contr IA
C1525091|Femoral artery and Popliteal artery Fluoroscopic angiogram Angioplasty W contrast IA
C1525091|Angioplasty^W contrast IA:Find:Pt:Femoral artery+Popliteal artery:Doc:XR.fluor.angio
C1525091|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Femoral artery+Popliteal artery:Document:XR.fluor.angio
C1830188|Guidance for biopsy.needle:Finding:Point in time:To be specified in another part of the message:Narrative:COMPUTERIZED TOMOGRAPHY
C1830188|CT Guidance for needle biopsy of Unspecified body region
C1830188|XXX CT Bx needle guid
C1830188|Guidance for biopsy.needle:Find:Pt:XXX:Doc:CT
C1830188|Guidance for biopsy.needle:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1830199|Mastoid-Bl CT
C1830199|Mastoid - bilateral CT
C1830199|Multisection:Finding:Point in time:Mastoid.bilateral:Document:Computerized Tomography
C1830199|Multisection:Find:Pt:Mastoid.bilateral:Doc:CT
C1830253|Breast duct Mammogram during surgery W contrast intra duct
C1830253|Brst.duct Mam in Surg W contr intra Dct
C1830253|Views^during surgery W contrast intra duct:Find:Pt:Breast.duct:Doc:Mam
C1830253|Views^during surgery W contrast intra duct:Finding:Point in time:Breast.duct:Document:Mam
C1830089|Artery US
C1830089|Multisection:Finding:Point in time:To be specified in another part of the message artery:Document:Ultrasound
C1830089|Multisection:Find:Pt:XXX artery:Doc:US
C1831072|Knee-L XR GE 4V
C1831072|Knee - left X-ray GE 4 views
C1831072|Views GE 4:Find:Pt:Knee.left:Doc:XR
C1831072|Views GE 4:Finding:Point in time:Knee.left:Document:XR
C1715432|US Guidance for drainage of abscess of Subphrenic space
C1715432|Guidance for drainage of abscess:Finding:Point in time:Subphrenic space:Document:Ultrasound
C1715432|Subphrenic Space US Abscess drain guid
C1715432|Guidance for drainage of abscess:Find:Pt:Subphrenic space:Doc:US
C1715494|SM ves DOP
C1715494|Superior mesenteric vessels US.doppler
C1715494|Multisection:Find:Pt:Superior mesenteric vessels:Doc:US.doppler
C1715494|Multisection:Finding:Point in time:Superior mesenteric vessels:Document:Ultrasound.doppler
C1644646|Upper extremity artery - right US
C1644646|UE a-R US
C1644646|Multisection:Find:Pt:Upper extremity artery.right:Doc:US
C1644646|Multisection:Finding:Point in time:Upper extremity artery.right:Document:Ultrasound
C1648287|LE a-R US
C1648287|Lower extremity artery - right US
C1648287|Multisection:Find:Pt:Lower extremity artery.right:Doc:US
C1648287|Multisection:Finding:Point in time:Lower extremity artery.right:Document:Ultrasound
C1644151|Hand - left X-ray limited
C1644151|Hand-L XR Ltd
C1644151|Views limited:Find:Pt:Hand.left:Doc:XR
C1644151|Views limited:Finding:Point in time:Hand.left:Document:XR
C1644154|Prostate SPECT W In-111 Satmb IV
C1644154|Prostate SPECT W In-111 Satumomab IV
C1644154|Multisection^W In-111 Satumomab Intravenous:Finding:Point in time:Prostate:Document:Radnuc.SPECT
C1644154|Multisection^W In-111 Satumomab IV:Find:Pt:Prostate:Doc:Radnuc.SPECT
C1634507|Ankle-L XR Lat+Mortise+Broden W Stress
C1634507|Ankle - left X-ray lateral and Mortise and Broden W manual stress
C1634507|Views lateral & Mortise & Broden^W manual stress:Finding:Point in time:Ankle.left:Document:XR
C1634507|Views lateral & Mortise & Broden^W manual stress:Find:Pt:Ankle.left:Doc:XR
C1635006|Foot sesamoid bones - bilateral X-ray
C1635006|Views:Find:Pt:Foot.sesamoid bones.bilateral:Doc:XR
C1635006|Views:Finding:Point in time:Foot.sesamoid bones.bilateral:Document:XR
C1635006|Ft.Sesamoids-Bl XR
C1644666|Unspecified body region X-ray post mortem
C1644666|XXX XR PM
C1644666|Views post mortem:Finding:Point in time:To be specified in another part of the message:Document:XR
C1644666|Views post mortem:Find:Pt:XXX:Doc:XR
C1714798|Views^W furosemide & W radionuclide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1714798|Kidney - bilateral Scan W furosemide and W radionuclide IV
C1714798|Views^W furosemide & W radionuclide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1714798|Kdny-Bl RI W Furosemide+RNC IV
C1714818|Knee - right X-ray GE 3 views
C1714818|Knee-R XR GE 3V
C1714818|Views GE 3:Find:Pt:Knee.right:Doc:XR
C1714818|Views GE 3:Finding:Point in time:Knee.right:Document:XR
C1714784|Multisection for tumor whole body:Find:Pt:^Patient:Doc:CT
C1714784|Deprecated CT for tumor whole body
C1714784|Multisection for tumor whole body:Finding:Point in time:^Patient:Document:Computerized Tomography
C1714784|Deprecated CT for Tumor WB
C1635611|L-spine XR AP+Lat+Obl+Spot stand
C1635611|Views AP & lateral & oblique & spot^standing:Find:Pt:Spine.lumbar:Doc:XR
C1635611|Views AP & lateral & oblique & spot^standing:Finding:Point in time:Spine.lumbar:Document:XR
C1635611|Lumbar spine X-ray AP and lateral and oblique and spot standing
C1638455|Should-L XR 90 Deg Abduction
C1638455|Shoulder - left X-ray 90 degree abduction
C1638455|Views 90 degree abduction:Find:Pt:Shoulder.left:Doc:XR
C1638455|Views 90 degree abduction:Finding:Point in time:Shoulder.left:Document:XR
C1639906|Extr v-L US
C1639906|Extremity vein - left US
C1639906|Multisection:Finding:Point in time:Extremity vein.left:Document:Ultrasound
C1639906|Multisection:Find:Pt:Extremity vein.left:Doc:US
C1633388|Gastrointestine upper Fluoroscopy W gastrografin PO
C1633388|UGI Flr W Gastrografin PO
C1633388|Views^W gastrografin Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1633388|Views^W gastrografin PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1633403|Liver Flr Tube plac guid
C1633403|Fluoroscopy Guidance for placement of tube in Liver
C1633403|Guidance for placement of tube:Finding:Point in time:Liver:Document:XR.fluor
C1633403|Guidance for placement of tube:Find:Pt:Liver:Doc:XR.fluor
C1644664|Orbit+Face MRI
C1644664|Orbit and Face MRI
C1644664|Multisection:Find:Pt:Orbit+Face:Doc:MRI
C1644664|Multisection:Finding:Point in time:Orbit+Face:Document:MRI
C1954874|Views^W radionuclide Intravenous:Finding:Point in time:To be specified in another part of the message:Narrative:Radnuc
C1954874|Unspecified body region Scan
C1954874|XXX RI W RNC IV
C1954874|Views^W radionuclide IV:Find:Pt:XXX:Doc:Radnuc
C1954874|Views^W radionuclide Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Radnuc
C1977325|Heart SPECT perfusion and wall motion at rest and W stress and W Tl-201 IV and W Tc-99m Sestamibi IV
C1977325|Hrt SPECT PF+WM R+S+W Tl201+Tc99mMIBI IV
C1977325|Multisection perfusion & wall motion^at rest & W stress & W Tl-201 IV & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1977325|Multisection perfusion & wall motion^at rest & W stress & W Tl-201 Intravenous & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1977329|RI Ltd W I-131 mIBG IV
C1977329|Scan limited W I-131 MIBG IV
C1977329|Views limited^W I-131 MIBG Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1977329|Views limited^W I-131 MIBG IV:Find:Pt:^Patient:Doc:Radnuc
C2925708|Multisection & 3D reconstruction^W contrast Intravenous:Finding:Point in time:Chest>Coronary arteries:Document:Computerized Tomography.angio
C2925708|Multisection & 3D reconstruction^W contrast IV:Find:Pt:Chest>Coronary arteries:Doc:CT.angio
C2925708|Deprecated Chest>CA CT.Angio +3DR W cont
C2925708|Deprecated Chest>Coronary arteries CT angiogram and 3D reconstruction W contrast IV
C3533558|Guidance for removal of percutaneous nephrostomy tube^W contrast:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C3533558|Fluoroscopy Guidance for removal of percutaneous nephrostomy tube from Kidney - bilateral-- W contrast
C3533558|Guidance for removal of percutaneous nephrostomy tube^W contrast:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C3533558|Kdny-Bl Flr PNT removal guid W contr
C3533548|Guidance for trigger point injection:Find:Pt:Muscle:Doc:XR.fluor
C3533548|Fluoroscopy Guidance for trigger point injection of Muscle
C3533548|Muscle Flr TPI guid
C3533548|Guidance for trigger point injection:Finding:Point in time:Muscle:Document:XR.fluor
C3262930|Multisection^W contrast IS:Find:Pt:Wrist.left:Doc:CT
C3262930|Wrist - left CT W contrast IS
C3262930|Multisection^W contrast Intrasynovial:Finding:Point in time:Wrist.left:Document:Computerized Tomography
C3262930|Wrist-L CT W contr IS
C3262940|Scapula CT
C3262940|Multisection:Finding:Point in time:Scapula:Document:Computerized Tomography
C3262940|Multisection:Find:Pt:Scapula:Doc:CT
C3262950|Guidance for biopsy.needle:Find:Pt:Chest>Pleura:Doc:XR.fluor
C3262950|Guidance for biopsy.needle:Finding:Point in time:Chest>Pleura:Document:XR.fluor
C3262950|Chest Pleura Flr Bx needle guid
C3262950|Fluoroscopy Guidance for needle biopsy of Chest Pleura
C3262966|Knee-L XR AP+Lat Xtable
C3262966|Knee - left X-ray AP and lateral crosstable
C3262966|Views AP & lateral crosstable:Finding:Point in time:Knee.left:Document:XR
C3262966|Views AP & lateral crosstable:Find:Pt:Knee.left:Doc:XR
C3263083|Skull X-ray PA and lateral and Waters and Towne
C3263083|Skull XR PA+lateral+Waters+Towne
C3263083|Views PA & lateral & Waters & Towne:Find:Pt:Skull:Doc:XR
C3263083|Views PA & lateral & Waters & Towne:Finding:Point in time:Skull:Document:XR
C3263084|SB Flr W cntr via ileostomy
C3263084|Small bowel Fluoroscopy W contrast via ileostomy
C3263084|Views^W contrast via ileostomy:Find:Pt:Small bowel:Doc:XR.fluor
C3263084|Views^W contrast via ileostomy:Finding:Point in time:Small bowel:Document:XR.fluor
C3263097|Extremity artery - right US
C3263097|Extr a-R US
C3263097|Multisection:Finding:Point in time:Extremity artery.right:Document:Ultrasound
C3263097|Multisection:Find:Pt:Extremity artery.right:Doc:US
C3262888|Abd XR AP+Lat Xtable
C3262888|Abdomen X-ray AP and lateral crosstable
C3262888|Views AP & lateral crosstable:Find:Pt:Abdomen:Doc:XR
C3262888|Views AP & lateral crosstable:Finding:Point in time:Abdomen:Document:XR
C3262891|Brst-Bl Mam Needle local guid
C3262891|Mammogram Guidance for needle localization of Breast - bilateral
C3262891|Guidance for needle localization:Finding:Point in time:Breast.bilateral:Document:Mam
C3262891|Guidance for needle localization:Find:Pt:Breast.bilateral:Doc:Mam
C0944152|Views:Finding:Point in time:Pelvis:Narrative:XR
C0944152|Pelvis X-ray
C0944152|Pelvis XR
C0944152|Views:Find:Pt:Pelvis:Doc:XR
C0944152|Views:Finding:Point in time:Pelvis:Document:XR
C0942163|Ribs - right X-ray
C0942163|Ribs-R XR
C0942163|Views:Find:Pt:Ribs.right:Doc:XR
C0942163|Views:Finding:Point in time:Ribs.right:Document:XR
C0942172|Thumb-R XR
C0942172|Thumb - right X-ray
C0942172|Views:Find:Pt:Thumb.right:Doc:XR
C0942172|Views:Finding:Point in time:Thumb.right:Document:XR
C0945320|Extr-L CT W contr IV
C0945320|Extremity - left CT W contrast IV
C0945320|Multisection^W contrast IV:Find:Pt:Extremity.left:Doc:CT
C0945320|Multisection^W contrast Intravenous:Finding:Point in time:Extremity.left:Document:Computerized Tomography
C0942207|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder.left:Document:MRI
C0942207|Should-L MRI WO+W contr IV
C0942207|Multisection^WO & W contrast IV:Find:Pt:Shoulder.left:Doc:MRI
C0942207|Shoulder - left MRI WO and W contrast IV
C0942214|Ankle-R MRI
C0942214|Ankle - right MRI
C0942214|Multisection:Finding:Point in time:Ankle.right:Document:MRI
C0942214|Multisection:Find:Pt:Ankle.right:Doc:MRI
C2709262|Deprecated Thigh Right MRI Multisection
C2709262|Multisection:Find:Pt:Thigh.right:Nar:MRI
C2709262|Deprecated Thigh-R MRI
C2709262|Multisection:Finding:Point in time:Thigh.right:Narrative:MRI
C0942292|Vein-L XRA Stent plac guid
C0942292|Fluoroscopic angiogram Guidance for placement of stent in Vein - left
C0942292|Guidance for placement of stent:Find:Pt:Vein.left:Doc:XR.fluor.angio
C0942292|Guidance for placement of stent:Finding:Point in time:Vein.left:Document:XR.fluor.angio
C0882039|Neck Flr W contr intra Lary
C0882039|Neck Fluoroscopy W contrast intra larynx
C0882039|Views^W contrast intra larynx:Find:Pt:Neck:Doc:XR.fluor
C0882039|Views^W contrast intra larynx:Finding:Point in time:Neck:Document:XR.fluor
C0882101|Skull XR 3V
C0882101|Skull X-ray 3 views
C0882101|Views 3:Find:Pt:Skull:Doc:XR
C0882101|Views 3:Finding:Point in time:Skull:Document:XR
C0882108|Spine US
C0882108|Multisection:Finding:Point in time:Spine:Document:Ultrasound
C0882108|Multisection:Find:Pt:Spine:Doc:US
C0882554|C-spine XR AP+Lat
C0882554|Views AP & lateral:Find:Pt:Spine.cervical:Doc:XR
C0882554|Views AP & lateral:Finding:Point in time:Spine.cervical:Document:XR
C0882554|Cervical spine X-ray AP and lateral
C0882135|Fluoroscopy Guidance for aspiration of Spine Lumbar Space
C0882135|L-spine space Flr Asp guid
C0882135|Guidance for aspiration:Finding:Point in time:Spine.lumbar space:Document:XR.fluor
C0882135|Guidance for aspiration:Find:Pt:Spine.lumbar space:Doc:XR.fluor
C0942112|Scrotum+Test-L RI W Tc99mP IV
C0942112|Scrotum and Testicle - left Scan W Tc-99m pertechnetate IV
C0942112|Views^W Tc-99m pertechnetate Intravenous:Finding:Point in time:Scrotum+Testicle.left:Document:Radnuc
C0942112|Views^W Tc-99m pertechnetate IV:Find:Pt:Scrotum+Testicle.left:Doc:Radnuc
C0942137|Deprecated Views:Finding:Point in time:Femur.left:Narrative:XR.DEXA
C0942137|Deprecated Femur-L DEXA
C0942137|Views:Find:Pt:Femur.left:Nar:XR.DEXA
C0942137|Views:Finding:Point in time:Femur.left:Narrative:XR.DEXA
C0942137|Deprecated Femur- left DEXA Bone density
C0942148|AC joint-Bl XR
C0942148|Acromioclavicular joint - bilateral X-ray
C0942148|Views:Finding:Point in time:Acromioclavicular joint.bilateral:Document:XR
C0942148|Views:Find:Pt:Acromioclavicular joint.bilateral:Doc:XR
C0881803|Abdomen X-ray AP upright portable
C0881803|Abd XR AP Upr port
C0881803|View AP upright portable:Finding:Point in time:Abdomen:Document:XR
C0881803|View AP upright portable:Find:Pt:Abdomen:Doc:XR
C0881812|BDs+GB Flr in Surg W contr BD
C0881812|Biliary ducts and Gallbladder Fluoroscopy during surgery W contrast biliary duct
C0881812|Views^during surgery W contrast biliary duct:Finding:Point in time:Biliary ducts+Gallbladder:Document:XR.fluor
C0881812|Views^during surgery W contrast biliary duct:Find:Pt:Biliary ducts+Gallbladder:Doc:XR.fluor
C0881819|Brach a+Subclavian a XRA W contr IA
C0881819|Brachial artery and Subclavian artery Fluoroscopic angiogram W contrast IA
C0881819|Views^W contrast IA:Find:Pt:Brachial artery+Subclavian artery:Doc:XR.fluor.angio
C0881819|Views^W contrast Intra-arterial:Finding:Point in time:Brachial artery+Subclavian artery:Document:XR.fluor.angio
C0881832|Brst specimen US
C0881832|Breast specimen US
C0881832|Multisection:Finding:Point in time:Breast specimen:Document:Ultrasound
C0881832|Multisection:Find:Pt:Breast specimen:Doc:US
C0881849|Carotid artery US
C0881849|Carot a US
C0881849|Multisection:Finding:Point in time:Carotid artery:Document:Ultrasound
C0881849|Multisection:Find:Pt:Carotid artery:Doc:US
C0881858|Multisection:Finding:Point in time:Chest:Narrative:COMPUTERIZED TOMOGRAPHY
C0881858|Chest CT
C0881858|Multisection:Find:Pt:Chest:Doc:CT
C0881858|Multisection:Finding:Point in time:Chest:Document:Computerized Tomography
C0881911|LE XR
C0881911|Lower extremity X-ray
C0881911|Views:Finding:Point in time:Lower extremity:Document:XR
C0881911|Views:Find:Pt:Lower extremity:Doc:XR
C0881919|Face CT W contr IV
C0881919|Multisection^W contrast Intravenous:Finding:Point in time:Facial bones:Document:Computerized Tomography
C0881919|Multisection^W contrast IV:Find:Pt:Facial bones:Doc:CT
C0881919|Facial bones CT W contrast IV
C1114533|TMJ XRTomo
C1114533|Temporomandibular joint X-ray tomograph
C1114533|Multisection:Find:Pt:Temporomandibular joint:Doc:XR.tomo
C1114533|Multisection:Finding:Point in time:Temporomandibular joint:Document:XR.tomo
C2608009|Views portable:Finding:Point in time:Skull:Narrative:XR
C2608009|Skull XR port
C2608009|Skull X-ray portable
C2608009|Views portable:Find:Pt:Skull:Doc:XR
C2608009|Views portable:Finding:Point in time:Skull:Document:XR
C1114546|Chest XR R+L Obl port
C1114546|Chest X-ray right and left oblique portable
C1114546|Views R- & L-oblique portable:Find:Pt:Chest:Doc:XR
C1114546|Views R- & L-oblique portable:Finding:Point in time:Chest:Document:XR
C1116467|Chest XR PA+Lat+R-Obl+L-Obl port
C1116467|Chest X-ray PA and lateral and right oblique and left oblique portable
C1116467|Views PA & lateral & R-oblique & L-oblique portable:Find:Pt:Chest:Doc:XR
C1116467|Views PA & lateral & R-oblique & L-oblique portable:Finding:Point in time:Chest:Document:XR
C1114655|Head vessels MRI angiogram
C1114655|Head ves MRI.Angio
C1114655|Multisection:Finding:Point in time:Head vessels:Document:MRI.angio
C1114655|Multisection:Find:Pt:Head vessels:Doc:MRI.angio
C1114956|Ft ves MRI.Angio
C1114956|Foot vessels MRI angiogram
C1114956|Multisection:Find:Pt:Foot vessels:Doc:MRI.angio
C1114956|Multisection:Finding:Point in time:Foot vessels:Document:MRI.angio
C1114673|US Guidance for aspiration of Unspecified body region
C1114673|XXX US Asp guid
C1114673|Guidance for aspiration:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1114673|Guidance for aspiration:Find:Pt:XXX:Doc:US
C1114680|Pelvis.symphysis pubis XR
C1114680|Pelvis symphysis pubis X-ray
C1114680|Views:Finding:Point in time:Pelvis.symphysis pubis:Document:XR
C1114680|Views:Find:Pt:Pelvis.symphysis pubis:Doc:XR
C1114463|Fluoroscopy Guidance for injection of Hip
C1114463|Hip Flr Inj guid
C1114463|Guidance for injection:Find:Pt:Hip:Doc:XR.fluor
C1114463|Guidance for injection:Finding:Point in time:Hip:Document:XR.fluor
C1543766|Hrt RI PF W Tl-201 IV
C1543766|Heart Scan perfusion W Tl-201 IV
C1543766|Views perfusion^W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1543766|Views perfusion^W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542850|SPECT Guidance for localization of tumor limited
C1542850|SPECT Tum local guid Ltd W RNC IV
C1542850|Guidance for localization of tumor limited^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1542850|Guidance for localization of tumor limited^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543804|SPECT Guidance for localization of tumor
C1543804|SPECT Tum local guid W RNC IV
C1543804|Guidance for localization of tumor^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543804|Guidance for localization of tumor^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543857|Bone Scan static
C1543857|Bone RI Static W RNC IV
C1543857|Views static^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543857|Views static^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543869|RI for ETr WB W I-131 mIBG IV
C1543869|Scan for endocrine tumor whole body W I-131 MIBG IV
C1543869|Views for endocrine tumor whole body^W I-131 MIBG IV:Find:Pt:^Patient:Doc:Radnuc
C1543869|Views for endocrine tumor whole body^W I-131 MIBG Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542898|Views ventilation^W radionuclide gaseous IH:Find:Pt:Lung:Doc:Radnuc
C1542898|Lung Scan ventilation W radionuclide gaseous IH
C1542898|Views ventilation^W radionuclide gaseous Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1542898|Lung RI V W RNC Gas IH
C1543879|PV shunt RI for Pat W RNC IT
C1543879|Peritoneovenous shunt Scan for patency W radionuclide IT
C1543879|Views for shunt patency^W radionuclide IT:Find:Pt:Peritoneovenous shunt:Doc:Radnuc
C1543879|Views for shunt patency^W radionuclide Intrathecal:Finding:Point in time:Peritoneovenous shunt:Document:Radnuc
C1543886|Thyroid RI Flow W RNC IV
C1543886|Thyroid Scan flow
C1543886|Views flow^W radionuclide IV:Find:Pt:Thyroid:Doc:Radnuc
C1543886|Views flow^W radionuclide Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1542923|Hrt RI FP W Stress+W Tc99mMIBI IV
C1542923|Heart Scan first pass W stress and W Tc-99m Sestamibi IV
C1542923|Views first pass^W stress & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1542923|Views first pass^W stress & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542855|RI for Tumor Mul Areas W Ga-67 IV
C1542855|Views for tumor multiple areas^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542855|Views for tumor multiple areas^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1542855|Scan for tumor multiple areas W Ga-67 IV
C1543509|UE ves-L DOP
C1543509|Upper extremity vessels - left US.doppler
C1543509|Multisection:Find:Pt:Upper extremity vessels.left:Doc:US.doppler
C1543509|Multisection:Finding:Point in time:Upper extremity vessels.left:Document:Ultrasound.doppler
C1543510|Lower extremity artery US.doppler
C1543510|LE a DOP
C1543510|Multisection:Finding:Point in time:Lower extremity artery:Document:Ultrasound.doppler
C1543510|Multisection:Find:Pt:Lower extremity artery:Doc:US.doppler
C1543174|Ribs X-ray lateral
C1543174|Ribs XR Lat
C1543174|View lateral:Finding:Point in time:Ribs:Document:XR
C1543174|View lateral:Find:Pt:Ribs:Doc:XR
C1543592|Should XR Stryker Notch+ West Point
C1543592|Shoulder X-ray Stryker Notch and West Point
C1543592|View Stryker Notch & West Point:Find:Pt:Shoulder:Doc:XR
C1543592|View Stryker Notch & West Point:Finding:Point in time:Shoulder:Document:XR
C1543683|SPECT Guidance for abscess localization
C1543683|SPECT Abscess local guid W RNC IV
C1543683|Guidance for abscess localization^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543683|Guidance for abscess localization^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1524257|Should-R XR AP+Ax+Outlet+Zanca
C1524257|Shoulder - right X-ray AP and axillary and outlet and Zanca
C1524257|Views AP & axillary & outlet & Zanca:Find:Pt:Shoulder.right:Doc:XR
C1524257|Views AP & axillary & outlet & Zanca:Finding:Point in time:Shoulder.right:Document:XR
C1526754|Olecranon - right X-ray
C1526754|Olecranon-R XR
C1526754|Views:Find:Pt:Olecranon.right:Doc:XR
C1526754|Views:Finding:Point in time:Olecranon.right:Document:XR
C1526756|Ac arch+Subclavian a-R XRA W contr IA
C1526756|Aortic arch and Subclavian artery - right Fluoroscopic angiogram W contrast IA
C1526756|Views^W contrast IA:Find:Pt:Aortic arch+Subclavian artery.right:Doc:XR.fluor.angio
C1526756|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Subclavian artery.right:Document:XR.fluor.angio
C1543702|Brain SPECT W Tc99mDTPA IV
C1543702|Brain SPECT W Tc-99m DTPA IV
C1543702|Multisection^W Tc-99m DTPA Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1543702|Multisection^W Tc-99m DTPA IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1543703|Brain SPECT W Tc99mGHA IV
C1543703|Brain SPECT W Tc-99m glucoheptonate IV
C1543703|Multisection^W Tc-99m glucoheptonate IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1543703|Multisection^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1542969|GB RI W Tc99mDISIDA IV
C1542969|Gallbladder Scan W Tc-99m DISIDA IV
C1542969|Views^W Tc-99m DISIDA Intravenous:Finding:Point in time:Gallbladder:Document:Radnuc
C1542969|Views^W Tc-99m DISIDA IV:Find:Pt:Gallbladder:Doc:Radnuc
C1526813|Ribs - left X-ray lateral
C1526813|Ribs-L XR Lat
C1526813|View lateral:Finding:Point in time:Ribs.left:Document:XR
C1526813|View lateral:Find:Pt:Ribs.left:Doc:XR
C1526816|Wrist-L XR AP+Lat
C1526816|Wrist - left X-ray AP and lateral
C1526816|Views AP & lateral:Find:Pt:Wrist.left:Doc:XR
C1526816|Views AP & lateral:Finding:Point in time:Wrist.left:Document:XR
C1543407|Should XR AP(w IR+ER)+Ax
C1543407|Shoulder X-ray AP (W internal rotation and W external rotation) and axillary
C1543407|Views AP (W internal rotation & W external rotation) & axillary:Find:Pt:Shoulder:Doc:XR
C1543407|Views AP (W internal rotation & W external rotation) & axillary:Finding:Point in time:Shoulder:Document:XR
C1524177|Should-Bl CT
C1524177|Shoulder - bilateral CT
C1524177|Multisection:Finding:Point in time:Shoulder.bilateral:Document:Computerized Tomography
C1524177|Multisection:Find:Pt:Shoulder.bilateral:Doc:CT
C1524178|Shoulder - left CT
C1524178|Should-L CT
C1524178|Multisection:Find:Pt:Shoulder.left:Doc:CT
C1524178|Multisection:Finding:Point in time:Shoulder.left:Document:Computerized Tomography
C1524185|Scrotum+Test MRI
C1524185|Scrotum and Testicle MRI
C1524185|Multisection:Finding:Point in time:Scrotum+Testicle:Document:MRI
C1524185|Multisection:Find:Pt:Scrotum+Testicle:Doc:MRI
C1524193|Vena cava MRI angiogram
C1524193|VC MRI.Angio
C1524193|Multisection:Find:Pt:Vena cava:Doc:MRI.angio
C1524193|Multisection:Finding:Point in time:Vena cava:Document:MRI.angio
C1524841|Upper extremity - bilateral CT WO contrast
C1524841|UE-Bl CT WO contr
C1524841|Multisection^WO contrast:Finding:Point in time:Upper extremity.bilateral:Document:Computerized Tomography
C1524841|Multisection^WO contrast:Find:Pt:Upper extremity.bilateral:Doc:CT
C1525113|UE vv-R MRI.Angio
C1525113|Upper extremity veins - right MRI angiogram
C1525113|Multisection:Find:Pt:Upper extremity veins.right:Doc:MRI.angio
C1525113|Multisection:Finding:Point in time:Upper extremity veins.right:Document:MRI.angio
C1525117|Abdominal vessels MRI angiogram
C1525117|Abd ves MRI.Angio
C1525117|Multisection:Find:Pt:Abdominal vessels:Doc:MRI.angio
C1525117|Multisection:Finding:Point in time:Abdominal vessels:Document:MRI.angio
C1524195|IVC MRI
C1524195|Inferior vena cava MRI
C1524195|Multisection:Finding:Point in time:Vena cava.inferior:Document:MRI
C1524195|Multisection:Find:Pt:Vena cava.inferior:Doc:MRI
C1524456|T-spine MRI Ltd W contr IV
C1524456|Multisection limited^W contrast Intravenous:Finding:Point in time:Spine.thoracic:Document:MRI
C1524456|Multisection limited^W contrast IV:Find:Pt:Spine.thoracic:Doc:MRI
C1524456|Thoracic spine MRI limited W contrast IV
C1525291|Ribs-L XR AP 1V
C1525291|Ribs - left X-ray AP single view
C1525291|View AP:Finding:Point in time:Ribs.left:Document:XR
C1525291|View AP:Find:Pt:Ribs.left:Doc:XR
C1525299|Hand - left X-ray Brewerton
C1525299|Hand-L XR Brewerton
C1525299|View Brewerton:Find:Pt:Hand.left:Doc:XR
C1525299|View Brewerton:Finding:Point in time:Hand.left:Document:XR
C1525195|UE joint-R MRI W contr IV
C1525195|Upper extremity joint - right MRI W contrast IV
C1525195|Multisection^W contrast IV:Find:Pt:Upper extremity.joint.right:Doc:MRI
C1525195|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.joint.right:Document:MRI
C1525261|Abd CT Asp+Drain tube plac guid
C1525261|CT Guidance for aspiration and placement of drainage tube of Abdomen
C1525261|Guidance for aspiration & placement of drainage tube:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1525261|Guidance for aspiration & placement of drainage tube:Find:Pt:Abdomen:Doc:CT
C1525272|Deprecated Unspecified body region CT stereotactic
C1525272|Deprecated XXX CT Stereo
C1525272|Multisection stereotactic:Find:Pt:XXX:Doc:CT
C1525272|Multisection stereotactic:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1525275|Adrenal CT W contr IV
C1525275|Adrenal gland CT W contrast IV
C1525275|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen>Adrenal gland:Document:Computerized Tomography
C1525275|Multisection^W contrast IV:Find:Pt:Abdomen>Adrenal gland:Doc:CT
C1525340|Chest XR L-Obl
C1525340|Chest X-ray left oblique
C1525340|View L-oblique:Finding:Point in time:Chest:Document:XR
C1525340|View L-oblique:Find:Pt:Chest:Doc:XR
C1525341|L-spine XR L-Obl
C1525341|View L-oblique:Find:Pt:Spine.lumbar:Doc:XR
C1525341|View L-oblique:Finding:Point in time:Spine.lumbar:Document:XR
C1525341|Lumbar spine X-ray left oblique
C1525349|Knee - bilateral X-ray Sunrise
C1525349|Knee-Bl XR Sunrise
C1525349|View Sunrise:Finding:Point in time:Knee.bilateral:Document:XR
C1525349|View Sunrise:Find:Pt:Knee.bilateral:Doc:XR
C1525489|L-spine XR AP+Lat port
C1525489|Views AP & lateral portable:Finding:Point in time:Spine.lumbar:Document:XR
C1525489|Views AP & lateral portable:Find:Pt:Spine.lumbar:Doc:XR
C1525489|Lumbar spine X-ray AP and lateral portable
C1524251|C-spine XR AP+Lat+Odont
C1524251|Views AP & lateral & odontoid:Finding:Point in time:Spine.cervical:Document:XR
C1524251|Views AP & lateral & odontoid:Find:Pt:Spine.cervical:Doc:XR
C1524251|Cervical spine X-ray AP and lateral and odontoid
C1525508|Knee-L XR AP+Lat+Sunrise
C1525508|Knee - left X-ray AP and lateral and Sunrise
C1525508|Views AP & lateral & Sunrise:Finding:Point in time:Knee.left:Document:XR
C1525508|Views AP & lateral & Sunrise:Find:Pt:Knee.left:Doc:XR
C1525535|Should-L XR Lat+Y
C1525535|Shoulder - left X-ray lateral and Y
C1525535|Views lateral & Y:Finding:Point in time:Shoulder.left:Document:XR
C1525535|Views lateral & Y:Find:Pt:Shoulder.left:Doc:XR
C1525542|Chest XR PA+Lat+AP Lat-Decub
C1525542|Chest X-ray PA and lateral and AP lateral-decubitus
C1525542|Views PA & lateral & AP lateral-decubitus:Finding:Point in time:Chest:Document:XR
C1525542|Views PA & lateral & AP lateral-decubitus:Find:Pt:Chest:Doc:XR
C1525595|Chest Fluoroscopy W contrast PO
C1525595|Chest Flr W contr PO
C1525595|Views^W contrast PO:Find:Pt:Chest:Doc:XR.fluor
C1525595|Views^W contrast Oral:Finding:Point in time:Chest:Document:XR.fluor
C1525608|CT Guidance for biopsy of Epididymis
C1525608|Guidance for biopsy:Finding:Point in time:Scrotum+Testicle>Epididymis:Document:Computerized Tomography
C1525608|Guidance for biopsy:Find:Pt:Scrotum+Testicle>Epididymis:Doc:CT
C1525608|Scrot+Test Epid CT Bx guid
C1525621|TMJ CT
C1525621|Temporomandibular joint CT
C1525621|Multisection:Find:Pt:Temporomandibular joint:Doc:CT
C1525621|Multisection:Finding:Point in time:Temporomandibular joint:Document:Computerized Tomography
C1525684|Sternoclavicular joint - bilateral X-ray
C1525684|SC joint-Bl XR
C1525684|Views:Find:Pt:Sternoclavicular joint.bilateral:Doc:XR
C1525684|Views:Finding:Point in time:Sternoclavicular joint.bilateral:Document:XR
C1525736|Extr vv-Bl XRA W contr IV
C1525736|Extremity veins - bilateral Fluoroscopic angiogram W contrast IV
C1525736|Views^W contrast IV:Find:Pt:Extremity veins.bilateral:Doc:XR.fluor.angio
C1525736|Views^W contrast Intravenous:Finding:Point in time:Extremity veins.bilateral:Document:XR.fluor.angio
C1525748|Wrist - bilateral X-ray tomograph
C1525748|Wrist-Bl XRTomo
C1525748|Multisection:Find:Pt:Wrist.bilateral:Doc:XR.tomo
C1525748|Multisection:Finding:Point in time:Wrist.bilateral:Document:XR.tomo
C1524690|Wrist MRI W contrast IS
C1524690|Multisection^W contrast Intrasynovial:Finding:Point in time:Wrist:Document:MRI
C1524690|Multisection^W contrast IS:Find:Pt:Wrist:Doc:MRI
C1524690|Wrist MRI W contr IS
C1525776|Clavicle-Bl XR 45 Deg Ceph Angle
C1525776|Clavicle - bilateral X-ray 45 degree cephalic angle
C1525776|View 45 degree cephalic angle:Finding:Point in time:Clavicle.bilateral:Document:XR
C1525776|View 45 degree cephalic angle:Find:Pt:Clavicle.bilateral:Doc:XR
C1525789|Humerus XR AP+Transthoracic
C1525789|Humerus X-ray AP and transthoracic
C1525789|Views AP & transthoracic:Find:Pt:Humerus:Doc:XR
C1525789|Views AP & transthoracic:Finding:Point in time:Humerus:Document:XR
C1525856|Knee XR W Stress
C1525856|Knee X-ray W manual stress
C1525856|Views^W manual stress:Finding:Point in time:Knee:Document:XR
C1525856|Views^W manual stress:Find:Pt:Knee:Doc:XR
C1525894|Orbit - bilateral X-ray 4 views
C1525894|Orbit-Bl XR 4V
C1525894|Views 4:Find:Pt:Orbit.bilateral:Doc:XR
C1525894|Views 4:Finding:Point in time:Orbit.bilateral:Document:XR
C1525830|Great toe-Bl XR
C1525830|Great toe - bilateral X-ray
C1525830|Views:Find:Pt:Great toe.bilateral:Doc:XR
C1525830|Views:Finding:Point in time:Great toe.bilateral:Document:XR
C1526000|Elbow-R XR AP+Lat
C1526000|Elbow - right X-ray AP and lateral
C1526000|Views AP & lateral:Find:Pt:Elbow.right:Doc:XR
C1526000|Views AP & lateral:Finding:Point in time:Elbow.right:Document:XR
C1526011|Finger - right X-ray 3 views
C1526011|Finger-R XR 3V
C1526011|Views 3:Find:Pt:Finger.right:Doc:XR
C1526011|Views 3:Finding:Point in time:Finger.right:Document:XR
C1526013|Foot - right X-ray 2 views
C1526013|Ft-R XR 2V
C1526013|Views 2:Find:Pt:Foot.right:Doc:XR
C1526013|Views 2:Finding:Point in time:Foot.right:Document:XR
C1526043|Hip - right X-ray lateral crosstable
C1526043|Hip-R XR Lat Xtable
C1526043|Hip-R XR +Lat Xtable
C1526043|Hip - right X-ray and lateral crosstable
C1526043|Views & lateral crosstable:Find:Pt:Hip.right:Doc:XR
C1526043|View lateral crosstable:Find:Pt:Hip.right:Doc:XR
C1526043|View lateral crosstable:Finding:Point in time:Hip.right:Document:XR
C1526043|Views & lateral crosstable:Finding:Point in time:Hip.right:Document:XR
C1526069|Knee - right X-ray W manual stress
C1526069|Knee-R XR W Stress
C1526069|Views^W manual stress:Finding:Point in time:Knee.right:Document:XR
C1526069|Views^W manual stress:Find:Pt:Knee.right:Doc:XR
C1525130|Ribs - right X-ray 2 views
C1525130|Ribs-R XR 2V
C1525130|Views 2:Find:Pt:Ribs.right:Doc:XR
C1525130|Views 2:Finding:Point in time:Ribs.right:Document:XR
C1526100|Shoulder - right X-ray 5 views
C1526100|Should-R XR 5V
C1526100|Views 5:Find:Pt:Shoulder.right:Doc:XR
C1526100|Views 5:Finding:Point in time:Shoulder.right:Document:XR
C1526139|Should XR Y
C1526139|Shoulder X-ray Y
C1526139|View Y:Find:Pt:Shoulder:Doc:XR
C1526139|View Y:Finding:Point in time:Shoulder:Document:XR
C1526172|Thumb X-ray oblique single view
C1526172|Thumb XR Obl 1V
C1526172|View oblique:Finding:Point in time:Thumb:Document:XR
C1526172|View oblique:Find:Pt:Thumb:Doc:XR
C1526189|T-spine XR Lat Hyperext
C1526189|View lateral hyperextension:Finding:Point in time:Spine.thoracic:Document:XR
C1526189|View lateral hyperextension:Find:Pt:Spine.thoracic:Doc:XR
C1526189|Thoracic spine X-ray lateral hyperextension
C1524701|Upper extremity X-ray tomograph
C1524701|UE XRTomo
C1524701|Multisection:Finding:Point in time:Upper extremity:Document:XR.tomo
C1524701|Multisection:Find:Pt:Upper extremity:Doc:XR.tomo
C1524709|Wrist XR PA V1
C1524709|Wrist X-ray PA
C1524709|View PA:Find:Pt:Wrist:Doc:XR
C1524709|View PA:Finding:Point in time:Wrist:Document:XR
C1526217|Carotid artery.external - right Fluoroscopic angiogram W contrast IA
C1526217|Carot a.ext-R XRA W contr IA
C1526217|Views^W contrast IA:Find:Pt:Carotid artery.external.right:Doc:XR.fluor.angio
C1526217|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.external.right:Document:XR.fluor.angio
C1526225|Ribs lower - right X-ray
C1526225|Ribs.lower-R XR
C1526225|Views:Finding:Point in time:Ribs.lower.right:Document:XR
C1526225|Views:Find:Pt:Ribs.lower.right:Doc:XR
C1526249|Views Broden:Find:Pt:Calcaneus.left:Doc:XR
C1526249|Deprecated Heel-L XR Broden
C1526249|Views Broden:Finding:Point in time:Calcaneus.left:Document:XR
C1526249|Deprecated Calcaneus - left X-ray Broden
C1526255|Foot - left X-ray AP standing
C1526255|Ft-L XR AP stand
C1526255|Views AP^standing:Find:Pt:Foot.left:Doc:XR
C1526255|Views AP^standing:Finding:Point in time:Foot.left:Document:XR
C1526262|BDs+GB US
C1526262|Biliary ducts and Gallbladder US
C1526262|Multisection:Find:Pt:Biliary ducts+Gallbladder:Doc:US
C1526262|Multisection:Finding:Point in time:Biliary ducts+Gallbladder:Document:Ultrasound
C1527043|Kidney US
C1527043|Multisection:Finding:Point in time:Kidney:Narrative:Ultrasound
C1527043|Multisection:Finding:Point in time:Kidney:Document:Ultrasound
C1527043|Multisection:Find:Pt:Kidney:Doc:US
C1526277|Mediastinum US
C1526277|Multisection:Find:Pt:Mediastinum:Doc:US
C1526277|Multisection:Finding:Point in time:Mediastinum:Document:Ultrasound
C1526332|Neck XR 2V Lat
C1526332|Neck X-ray 2 views lateral
C1526332|Views 2 lateral:Find:Pt:Neck:Doc:XR
C1526332|Views 2 lateral:Finding:Point in time:Neck:Document:XR
C1525918|US Guidance for aspiration of cyst of Pancreas
C1525918|Pancreas US Cyst Asp guid
C1525918|Guidance for aspiration of cyst:Find:Pt:Pancreas:Doc:US
C1525918|Guidance for aspiration of cyst:Finding:Point in time:Pancreas:Document:Ultrasound
C1526339|Iliac ves-L US
C1526339|Iliac vessels - left US
C1526339|Multisection:Find:Pt:Iliac vessels.left:Doc:US
C1526339|Multisection:Finding:Point in time:Iliac vessels.left:Document:Ultrasound
C1526301|Ribs Ant-Bl XR
C1526301|Ribs anterior - bilateral X-ray
C1526301|Views:Finding:Point in time:Ribs.anterior.bilateral:Document:XR
C1526301|Views:Find:Pt:Ribs.anterior.bilateral:Doc:XR
C1526302|Ribs Ant-L XR
C1526302|Ribs anterior - left X-ray
C1526302|Views:Finding:Point in time:Ribs.anterior.left:Document:XR
C1526302|Views:Find:Pt:Ribs.anterior.left:Doc:XR
C1526314|Breast duct - left Mammogram W contrast intra duct
C1526314|Brst.duct-L Mam W contr intra Dct
C1526314|Views^W contrast intra duct:Finding:Point in time:Breast.duct.left:Document:Mam
C1526314|Views^W contrast intra duct:Find:Pt:Breast.duct.left:Doc:Mam
C1524880|Upper arm-R MRI WO contr
C1524880|Upper arm - right MRI WO contrast
C1524880|Multisection^WO contrast:Find:Pt:Upper arm.right:Doc:MRI
C1524880|Multisection^WO contrast:Finding:Point in time:Upper arm.right:Document:MRI
C1524915|Lower leg - left MRI WO contrast
C1524915|Lower leg-L MRI WO contr
C1524915|Multisection^WO contrast:Find:Pt:Lower leg.left:Doc:MRI
C1524915|Multisection^WO contrast:Finding:Point in time:Lower leg.left:Document:MRI
C1524569|Neck CT W contr IV
C1524569|Neck CT W contrast IV
C1524569|Multisection^W contrast IV:Find:Pt:Neck:Doc:CT
C1524569|Multisection^W contrast Intravenous:Finding:Point in time:Neck:Document:Computerized Tomography
C1524280|Extr a XRA Angpsty W contr IA
C1524280|Extremity artery Fluoroscopic angiogram Angioplasty W contrast IA
C1524280|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Extremity artery:Document:XR.fluor.angio
C1524280|Angioplasty^W contrast IA:Find:Pt:Extremity artery:Doc:XR.fluor.angio
C1524595|Lower leg-L MRI W contr IV
C1524595|Lower leg - left MRI W contrast IV
C1524595|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg.left:Document:MRI
C1524595|Multisection^W contrast IV:Find:Pt:Lower leg.left:Doc:MRI
C1524596|Lower leg-R CT W contr IV
C1524596|Lower leg - right CT W contrast IV
C1524596|Multisection^W contrast IV:Find:Pt:Lower leg.right:Doc:CT
C1524596|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg.right:Document:Computerized Tomography
C1524129|Multisection^WO & W contrast Intravenous:Finding:Point in time:Calcaneus.right:Document:Computerized Tomography
C1524129|Multisection^WO & W contrast IV:Find:Pt:Calcaneus.right:Doc:CT
C1524129|Deprecated Calcaneus - right CT WO and W contrast IV
C1524129|Deprecated Heel-R CT WO+W contr IV
C1524957|Femur X-ray oblique single view
C1524957|Femur XR Obl 1V
C1524957|View oblique:Find:Pt:Femur:Doc:XR
C1524957|View oblique:Finding:Point in time:Femur:Document:XR
C1524979|Pelvis+Hip-L XR
C1524979|Pelvis and Hip - left X-ray
C1524979|Views:Finding:Point in time:Pelvis+Hip.left:Document:XR
C1524979|Views:Find:Pt:Pelvis+Hip.left:Doc:XR
C1524320|CT Guidance for drainage of Pelvis
C1524320|Pelvis CT Drain guid
C1524320|Guidance for drainage:Find:Pt:Pelvis:Doc:CT
C1524320|Guidance for drainage:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1524349|Brst-L MRI
C1524349|Breast - left MRI
C1524349|Multisection:Finding:Point in time:Breast.left:Document:MRI
C1524349|Multisection:Find:Pt:Breast.left:Doc:MRI
C1524633|Foot - left X-ray 3 views
C1524633|Ft-L XR 3V
C1524633|Views 3:Finding:Point in time:Foot.left:Document:XR
C1524633|Views 3:Find:Pt:Foot.left:Doc:XR
C1524995|Coccyx XR 2V
C1524995|Coccyx X-ray 2 views
C1524995|Views 2:Find:Pt:Coccyx:Doc:XR
C1524995|Views 2:Finding:Point in time:Coccyx:Document:XR
C1524731|Foot - right CT WO and W contrast IV
C1524731|Ft-R CT WO+W contr IV
C1524731|Multisection^WO & W contrast Intravenous:Finding:Point in time:Foot.right:Document:Computerized Tomography
C1524731|Multisection^WO & W contrast IV:Find:Pt:Foot.right:Doc:CT
C1524393|Gallbladder X-ray tomograph
C1524393|GB XRTomo
C1524393|Multisection:Finding:Point in time:Gallbladder:Document:XR.tomo
C1524393|Multisection:Find:Pt:Gallbladder:Doc:XR.tomo
C1524394|Hand X-ray tomograph
C1524394|Hand XRTomo
C1524394|Multisection:Finding:Point in time:Hand:Document:XR.tomo
C1524394|Multisection:Find:Pt:Hand:Doc:XR.tomo
C1524405|Hip-Bl CT
C1524405|Hip - bilateral CT
C1524405|Multisection:Finding:Point in time:Hip.bilateral:Document:Computerized Tomography
C1524405|Multisection:Find:Pt:Hip.bilateral:Doc:CT
C1524425|Knee X-ray tomograph
C1524425|Knee XRTomo
C1524425|Multisection:Finding:Point in time:Knee:Document:XR.tomo
C1524425|Multisection:Find:Pt:Knee:Doc:XR.tomo
C1524771|Pancreas MRI WO and W contrast IV
C1524771|Pancreas MRI WO+W contr IV
C1524771|Multisection^WO & W contrast IV:Find:Pt:Pancreas:Doc:MRI
C1524771|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pancreas:Document:MRI
C1524787|Multisection^WO & W contrast IV:Find:Pt:Spine.lumbar:Doc:CT
C1524787|L-spine CT WO+W contr IV
C1524787|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1524787|Lumbar spine CT WO and W contrast IV
C1524807|Upper extremity vessels MRI angiogram WO and W contrast IV
C1524807|UE ves MRI.Angio WO+W contr IV
C1524807|Multisection^WO & W contrast IV:Find:Pt:Upper extremity vessels:Doc:MRI.angio
C1524807|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity vessels:Document:MRI.angio
C1525073|Knee-Bl XR Obl
C1525073|Knee - bilateral X-ray oblique
C1525073|Views oblique:Find:Pt:Knee.bilateral:Doc:XR
C1525073|Views oblique:Finding:Point in time:Knee.bilateral:Document:XR
C1830228|Chest CT W red contr vol IV
C1830228|Chest CT W reduced contrast volume IV
C1830228|Multisection^W reduced contrast volume IV:Find:Pt:Chest:Doc:CT
C1830228|Multisection^W reduced contrast volume Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C1830244|Wrist - right X-ray GE 3 views
C1830244|Wrist-R XR GE 3V
C1830244|Views GE 3:Finding:Point in time:Wrist.right:Document:XR
C1830244|Views GE 3:Find:Pt:Wrist.right:Doc:XR
C1830274|SPECT Guidance for superficial biopsy of Bone
C1830274|Bone SPECT Bx super guid W RNC IV
C1830274|Guidance for superficial biopsy^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1830274|Guidance for superficial biopsy^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1715467|Lung Flr PC Bx needle guid
C1715467|Fluoroscopy Guidance for percutaneous needle biopsy of Lung
C1715467|Guidance for percutaneous biopsy.needle:Find:Pt:Lung:Doc:XR.fluor
C1715467|Guidance for percutaneous biopsy.needle:Finding:Point in time:Lung:Document:XR.fluor
C1644153|LE a-L US
C1644153|Lower extremity artery - left US
C1644153|Multisection:Finding:Point in time:Lower extremity artery.left:Document:Ultrasound
C1644153|Multisection:Find:Pt:Lower extremity artery.left:Doc:US
C1632799|Ribs lower post-L XR
C1632799|Ribs lower posterior - left X-ray
C1632799|Views:Find:Pt:Ribs.lower.posterior.left:Doc:XR
C1632799|Views:Finding:Point in time:Ribs.lower.posterior.left:Document:XR
C1643612|Unspecified body region MRI cine for CSF flow
C1643612|XXX MRI Cine for CSF flow
C1643612|Multisection cine for CSF flow:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1643612|Multisection cine for CSF flow:Find:Pt:XXX:Doc:MRI
C1714792|Pulmonary system MRI
C1714792|Pulm MRI
C1714792|Multisection:Finding:Point in time:Pulmonary system:Document:MRI
C1714792|Multisection:Find:Pt:Pulmonary system:Doc:MRI
C1714800|Chest and Abdomen X-ray AP (supine and upright) and PA chest
C1714800|Chest+Abd XR AP (supine+Upr)+PA Chst
C1714800|Views AP (supine & upright) & PA chest:Find:Pt:Chest+Abdomen:Doc:XR
C1714800|Views AP (supine & upright) & PA chest:Finding:Point in time:Chest+Abdomen:Document:XR
C1714817|Joint XR W FE
C1714817|Joint X-ray W flexion and W extension
C1714817|Views^W flexion & W extension:Find:Pt:Joint:Doc:XR
C1714817|Views^W flexion & W extension:Finding:Point in time:Joint:Document:XR
C0882526|Views AP (R-lateral-decubitus & L-lateral-decubitus):Finding:Point in time:Chest:Narrative:XR
C0882526|Chest XR AP (R+L-Lat Decub)
C0882526|Deprecated Chest XR AP (R+L-Lat Decub)
C0882526|Views AP (R-lateral-decubitus & L-lateral-decubitus):Find:Pt:Chest:Nar:XR
C0882526|Deprecated Chest X-ray AP (R-lateral-decubitus & L-lateral-decubitus)
C0882526|Chest X-ray AP (right lateral-decubitus and left lateral-decubitus)
C0882526|Views AP (R-lateral-decubitus & L-lateral-decubitus):Find:Pt:Chest:Doc:XR
C0882526|Views AP (R-lateral-decubitus & L-lateral-decubitus):Finding:Point in time:Chest:Document:XR
C1705867|Deprecated Finger.3rd-R XR GE 3V
C1705867|Views GE 3:Find:Pt:Finger.third.right:Nar:XR
C1705867|Deprecated Finger third Right X-ray GE 3 views
C1705867|Views GE 3:Finding:Point in time:Finger.third.right:Narrative:XR
C1714942|Study observation.general:Imp:Pt:^Fetuses.twins:Nar:US
C1714942|Deprecated US Study Observation general
C1714942|Deprecated Study observation general of fetuses US
C1714942|Study observation.general:Impression/interpretation of study:Point in time:^Fetuses.twins:Narrative:Ultrasound
C1714948|Bladder+Urethra Flr W contr IB void
C1714948|Urinary Bladder and Urethra Fluoroscopy W contrast intra bladder during voiding
C1714948|Views^W contrast intra bladder during voiding:Finding:Point in time:Urinary bladder+Urethra:Document:XR.fluor
C1714948|Views^W contrast intra bladder during voiding:Find:Pt:Urinary bladder+Urethra:Doc:XR.fluor
C1715015|Foot sesamoid bones - left X-ray
C1715015|Ft.Sesamoids-L XR
C1715015|Views:Find:Pt:Foot.sesamoid bones.left:Doc:XR
C1715015|Views:Finding:Point in time:Foot.sesamoid bones.left:Document:XR
C1715019|Hrt RI for Infarct Ql+Qn W RNC IV
C1715019|Heart Scan for infarct qualitative and quantitative
C1715019|Views for infarct qualitative & quantitative^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1715019|Views for infarct qualitative & quantitative^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1715024|Liver+Spleen SPECT Flow W RNC IV
C1715024|Liver and Spleen SPECT flow
C1715024|Multisection flow^W radionuclide Intravenous:Finding:Point in time:Liver+Spleen:Document:Radnuc.SPECT
C1715024|Multisection flow^W radionuclide IV:Find:Pt:Liver+Spleen:Doc:Radnuc.SPECT
C1715036|Thyroid RI +Uptake W RNC IV
C1715036|Thyroid Scan and uptake
C1715036|Views & uptake^W radionuclide IV:Find:Pt:Thyroid:Doc:Radnuc
C1715036|Views & uptake^W radionuclide Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1637279|Ankle-L XR AP+Lat+Obl W Stress
C1637279|Ankle - left X-ray AP and lateral and oblique W manual stress
C1637279|Views AP & lateral & oblique^W manual stress:Find:Pt:Ankle.left:Doc:XR
C1637279|Views AP & lateral & oblique^W manual stress:Finding:Point in time:Ankle.left:Document:XR
C1635009|T+L-spine XR Scoli AP Stand+W+WO bending
C1635009|Spine Thoracic and Lumbar X-ray scoliosis AP standing and W right bending and W left bending and WO bending
C1635009|Views scoliosis AP^standing & W R-bending & W L-bending & WO bending:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1635009|Views scoliosis AP^standing & W R-bending & W L-bending & WO bending:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1646316|US Guidance for biopsy of Endomyocardium
C1646316|Endomyocardium US Bx guid
C1646316|Guidance for biopsy:Finding:Point in time:Endomyocardium:Document:Ultrasound
C1646316|Guidance for biopsy:Find:Pt:Endomyocardium:Doc:US
C1639532|UE ves graft-R DOP
C1639532|Upper extremity vessel graft - right US.doppler
C1639532|Multisection:Finding:Point in time:Upper extremity vessel graft.right:Document:Ultrasound.doppler
C1639532|Multisection:Find:Pt:Upper extremity vessel graft.right:Doc:US.doppler
C1639904|Deprecated Guidance for percutaneous biopsy.core needle:Find:Pt:Breast:Nar:Mam
C1639904|Deprecated Brst Mam PC Bx CN guid
C1639904|Deprecated Breast Mammogram Guidance for percutaneous biopsy.core needle
C1639904|Guidance for percutaneous biopsy.core needle:Find:Pt:Breast:Nar:Mam
C1639904|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast:Narrative:Mam
C1648947|Deprecated View AP portable:Finding:Point in time:Abdomen:Narrative:XR
C1648947|Deprecated Abdomen X-ray AP portable
C1648947|View AP portable:Find:Pt:Abdomen:Nar:XR
C1648947|Deprecated Abd XR AP port
C1648947|View AP portable:Finding:Point in time:Abdomen:Narrative:XR
C1977261|Breast duct - left Mammogram Single view W contrast intra duct
C1977261|Brst.duct-L Mam 1V W contr intra Dct
C1977261|View 1^W contrast intra duct:Find:Pt:Breast.duct.left:Doc:Mam
C1977261|View 1^W contrast intra duct:Finding:Point in time:Breast.duct.left:Document:Mam
C1953953|C-spine MRI W contr IT
C1953953|Multisection^W contrast IT:Find:Pt:Spine.cervical:Doc:MRI
C1953953|Multisection^W contrast Intrathecal:Finding:Point in time:Spine.cervical:Document:MRI
C1953953|Cervical spine MRI W contrast IT
C1953983|Breast implant - bilateral Mammogram diagnostic
C1953983|Brst implant-Bl Mam Dx
C1953983|Views diagnostic:Find:Pt:Breast implant.bilateral:Doc:Mam
C1953983|Views diagnostic:Finding:Point in time:Breast implant.bilateral:Document:Mam
C3262974|Should-L XR 3V+Y
C3262974|Shoulder - left X-ray 3 views and Y
C3262974|Views 3 & Y:Find:Pt:Shoulder.left:Doc:XR
C3262974|Views 3 & Y:Finding:Point in time:Shoulder.left:Document:XR
C3262976|Wrist - left X-ray lateral W flexion and W extension
C3262976|Wrist-L XR Lat W FE
C3262976|Views lateral^W flexion & W extension:Find:Pt:Wrist.left:Doc:XR
C3262976|Views lateral^W flexion & W extension:Finding:Point in time:Wrist.left:Document:XR
C3262985|Breast implant - bilateral MRI
C3262985|Brst implant-Bl MRI
C3262985|Multisection:Find:Pt:Breast implant.bilateral:Doc:MRI
C3262985|Multisection:Finding:Point in time:Breast implant.bilateral:Document:MRI
C3262987|Brst implant-Bl MRI W contr IV
C3262987|Breast implant - bilateral MRI W contrast IV
C3262987|Multisection^W contrast Intravenous:Finding:Point in time:Breast implant.bilateral:Document:MRI
C3262987|Multisection^W contrast IV:Find:Pt:Breast implant.bilateral:Doc:MRI
C3263000|Upper arm - bilateral MRI
C3263000|Upper arm-Bl MRI
C3263000|Multisection:Finding:Point in time:Upper arm.bilateral:Document:MRI
C3263000|Multisection:Find:Pt:Upper arm.bilateral:Doc:MRI
C3263004|Shoulder - bilateral MRI W contrast IV
C3263004|Should-Bl MRI W contr IV
C3263004|Multisection^W contrast IV:Find:Pt:Shoulder.bilateral:Doc:MRI
C3263004|Multisection^W contrast Intravenous:Finding:Point in time:Shoulder.bilateral:Document:MRI
C3483135|T-spine US CSF asp guid
C3483135|Guidance for CSF aspiration:Find:Pt:Spine.thoracic:Doc:US
C3483135|Guidance for CSF aspiration:Finding:Point in time:Spine.thoracic:Document:Ultrasound
C3483135|US Guidance for CSF aspiration of Thoracic spine
C3263013|Extr MRI
C3263013|Extremity MRI
C3263013|Multisection:Finding:Point in time:Extremity:Document:MRI
C3263013|Multisection:Find:Pt:Extremity:Doc:MRI
C3263047|Spleen SPECT W Tc-99m tagged RBC IV
C3263047|Spleen SPECT W Tc99mRBC IV
C3263047|Multisection^W Tc-99m tagged RBC IV:Find:Pt:Spleen:Doc:Radnuc.SPECT
C3263047|Multisection^W Tc-99m tagged RBC Intravenous:Finding:Point in time:Spleen:Document:Radnuc.SPECT
C3263052|Patella X-ray Sunrise
C3263052|Patella XR Sunrise
C3263052|View Sunrise:Finding:Point in time:Patella:Document:XR
C3263052|View Sunrise:Find:Pt:Patella:Doc:XR
C3263102|Wrist XR W clenched fist
C3263102|Wrist X-ray W clenched fist
C3263102|View^W clenched fist:Finding:Point in time:Wrist:Document:XR
C3263102|View^W clenched fist:Find:Pt:Wrist:Doc:XR
C3261470|View 1:Finding:Point in time:Calcaneus.left:Document:XR
C3261470|View 1:Find:Pt:Calcaneus.left:Doc:XR
C3261470|Deprecated Heel-R XR 1V
C3261470|Deprecated Calcaneus - right X-ray Single view
C3261470|Deprecated View 1:Find:Pt:Calcaneus.left:Doc:XR
C3262879|Aortic arch Fluoroscopic angiogram W contrast IA
C3262879|Ac arch XRA W contr IA
C3262879|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch:Document:XR.fluor.angio
C3262879|Views^W contrast IA:Find:Pt:Aortic arch:Doc:XR.fluor.angio
C0942151|Mastoid-Bl XR
C0942151|Mastoid - bilateral X-ray
C0942151|Views:Finding:Point in time:Mastoid.bilateral:Document:XR
C0942151|Views:Find:Pt:Mastoid.bilateral:Doc:XR
C0942164|Scapula - bilateral X-ray
C0942164|Scapula-Bl XR
C0942164|Views:Finding:Point in time:Scapula.bilateral:Document:XR
C0942164|Views:Find:Pt:Scapula.bilateral:Doc:XR
C0942175|Tib+Fib-R XR
C0942175|Tibia - right and Fibula - right X-ray
C0942175|Views:Find:Pt:Tibia.right+Fibula.right:Doc:XR
C0942175|Views:Finding:Point in time:Tibia.right+Fibula.right:Document:XR
C0942190|Extr-Bl CT W contr IV
C0942190|Extremity - bilateral CT W contrast IV
C0942190|Multisection^W contrast Intravenous:Finding:Point in time:Extremity.bilateral:Document:Computerized Tomography
C0942190|Multisection^W contrast IV:Find:Pt:Extremity.bilateral:Doc:CT
C0942201|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thigh.left:Document:MRI
C0942201|Multisection^WO & W contrast IV:Find:Pt:Thigh.left:Doc:MRI
C0942201|Thigh - left MRI WO and W contrast IV
C0942201|Thigh-L MRI WO+W contr IV
C0942209|Wrist - bilateral MRI WO and W contrast IV
C0942209|Wrist-Bl MRI WO+W contr IV
C0942209|Multisection^WO & W contrast IV:Find:Pt:Wrist.bilateral:Doc:MRI
C0942209|Multisection^WO & W contrast Intravenous:Finding:Point in time:Wrist.bilateral:Document:MRI
C0942216|Thoracic outlet - left MRI
C0942216|TO-L MRI
C0942216|Multisection:Finding:Point in time:Thoracic outlet.left:Document:MRI
C0942216|Multisection:Find:Pt:Thoracic outlet.left:Doc:MRI
C0942258|Popliteal space - left US
C0942258|Popliteal space-L US
C0942258|Multisection:Find:Pt:Popliteal space.left:Doc:US
C0942258|Multisection:Finding:Point in time:Popliteal space.left:Document:Ultrasound
C0942277|Knee - bilateral X-ray Merchants
C0942277|Knee-Bl XR Merchants
C0942277|View Merchants:Find:Pt:Knee.bilateral:Doc:XR
C0942277|View Merchants:Finding:Point in time:Knee.bilateral:Document:XR
C0942281|Breast - bilateral Mammogram limited
C0942281|Brst-Bl Mam Ltd
C0942281|Views limited:Finding:Point in time:Breast.bilateral:Document:Mam
C0942281|Views limited:Find:Pt:Breast.bilateral:Doc:Mam
C0942288|Cent v-L XRA Cath repos W contr IV
C0942288|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein - left-- W contrast IV
C0942288|Guidance for reposition of catheter^W contrast Intravenous:Finding:Point in time:Central vein.left:Document:XR.fluor.angio
C0942288|Guidance for reposition of catheter^W contrast IV:Find:Pt:Central vein.left:Doc:XR.fluor.angio
C0942291|Vein-Bl XRA Stent plac guid
C0942291|Fluoroscopic angiogram Guidance for placement of stent in Vein - bilateral
C0942291|Guidance for placement of stent:Find:Pt:Vein.bilateral:Doc:XR.fluor.angio
C0942291|Guidance for placement of stent:Finding:Point in time:Vein.bilateral:Document:XR.fluor.angio
C0942318|Cent v-Bl XRA CC change guid W contr IV
C0942318|Fluoroscopic angiogram Guidance for change of central catheter in Central vein - bilateral-- W contrast IV
C0942318|Guidance for change of central catheter^W contrast IV:Find:Pt:Central vein.bilateral:Doc:XR.fluor.angio
C0942318|Guidance for change of central catheter^W contrast Intravenous:Finding:Point in time:Central vein.bilateral:Document:XR.fluor.angio
C0942329|Brst-R Mam Cyst Asp guid
C0942329|Mammogram Guidance for aspiration of cyst of Breast - right
C0942329|Guidance for aspiration of cyst:Find:Pt:Breast.right:Doc:Mam
C0942329|Guidance for aspiration of cyst:Finding:Point in time:Breast.right:Document:Mam
C0945344|Knee - left X-ray AP single view standing
C0945344|Knee-L XR AP 1V stand
C0945344|View AP^standing:Finding:Point in time:Knee.left:Document:XR
C0945344|View AP^standing:Find:Pt:Knee.left:Doc:XR
C0942350|Iliac a-Bl XRA Angpsty W contr IA
C0942350|Iliac artery - bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C0942350|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Iliac artery.bilateral:Document:XR.fluor.angio
C0942350|Angioplasty^W contrast IA:Find:Pt:Iliac artery.bilateral:Doc:XR.fluor.angio
C0882063|Pelvis ves MRI.Angio W contr IV
C0882063|Pelvis vessels MRI angiogram W contrast IV
C0882063|Multisection^W contrast IV:Find:Pt:Pelvis vessels:Doc:MRI.angio
C0882063|Multisection^W contrast Intravenous:Finding:Point in time:Pelvis vessels:Document:MRI.angio
C0882069|Pituitary+ST MRI
C0882069|Pituitary and Sella turcica MRI
C0882069|Multisection:Finding:Point in time:Pituitary+Sella turcica:Document:MRI
C0882069|Multisection:Find:Pt:Pituitary+Sella turcica:Doc:MRI
C0882122|C-spine XR Swimmers
C0882122|View Swimmers:Find:Pt:Spine.cervical:Doc:XR
C0882122|View Swimmers:Finding:Point in time:Spine.cervical:Document:XR
C0882122|Cervical spine X-ray Swimmers
C0882127|L-spine CT W contr IV
C0882127|Multisection^W contrast IV:Find:Pt:Spine.lumbar:Doc:CT
C0882127|Multisection^W contrast Intravenous:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C0882127|Lumbar spine CT W contrast IV
C0882178|Uterus+FT Flr W contr IU
C0882178|Views^W contrast IU:Find:Pt:Uterus+Fallopian tubes:Doc:XR.fluor
C0882178|Views^W contrast Intrauterine:Finding:Point in time:Uterus+Fallopian tubes:Document:XR.fluor
C0882178|Uterus and Fallopian tubes Fluoroscopy W contrast IU
C0945314|Hip - right X-ray
C0945314|Hip-R XR
C0945314|Views:Find:Pt:Hip.right:Doc:XR
C0945314|Views:Finding:Point in time:Hip.right:Document:XR
C0942149|AC joint-L XR
C0942149|Acromioclavicular joint - left X-ray
C0942149|Views:Find:Pt:Acromioclavicular joint.left:Doc:XR
C0942149|Views:Finding:Point in time:Acromioclavicular joint.left:Document:XR
C0881776|Abdominal vessels US.doppler
C0881776|Abd ves DOP
C0881776|Multisection:Finding:Point in time:Abdominal vessels:Document:Ultrasound.doppler
C0881776|Multisection:Find:Pt:Abdominal vessels:Doc:US.doppler
C0881814|Urinary Bladder Aa XRA W contr IA
C0881814|Urinary bladder arteries Fluoroscopic angiogram W contrast IA
C0881814|Views^W contrast Intra-arterial:Finding:Point in time:Urinary bladder arteries:Document:XR.fluor.angio
C0881814|Views^W contrast IA:Find:Pt:Urinary bladder arteries:Doc:XR.fluor.angio
C0881828|Brain RI BD Protocol W Tc99mHMPAO IV
C0881828|Brain Scan brain death protocol W Tc-99m HMPAO IV
C0881828|Views brain death protocol^W Tc-99m HMPAO Intravenous:Finding:Point in time:Brain:Document:Radnuc
C0881828|Views brain death protocol^W Tc-99m HMPAO IV:Find:Pt:Brain:Doc:Radnuc
C0882521|Brst US Ltd
C0882521|Breast US limited
C0882521|Multisection limited:Finding:Point in time:Breast:Document:Ultrasound
C0882521|Multisection limited:Find:Pt:Breast:Doc:US
C0881847|Carotid artery extracranial Fluoroscopic angiogram Angioplasty W contrast IA
C0881847|Carot a.EC XRA Angpsty W contr IA
C0881847|Angioplasty^W contrast IA:Find:Pt:Carotid artery.extracranial:Doc:XR.fluor.angio
C0881847|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Carotid artery.extracranial:Document:XR.fluor.angio
C0881857|Centl v XRA Cath repos W contr IV
C0881857|Fluoroscopic angiogram Guidance for reposition of catheter in Central vein-- W contrast IV
C0881857|Guidance for reposition of catheter^W contrast IV:Find:Pt:Central vein:Doc:XR.fluor.angio
C0881857|Guidance for reposition of catheter^W contrast Intravenous:Finding:Point in time:Central vein:Document:XR.fluor.angio
C0881862|Unspecified body region Fluoroscopy Central vein catheter placement check
C0881862|XXX Flr CVC plac Ck
C0881862|Central vein catheter placement check:Find:Pt:XXX:Doc:XR.fluor
C0881862|Central vein catheter placement check:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C0881887|US Guidance for aspiration of Pleural space
C0881887|Pl space US Asp guid
C0881887|Guidance for aspiration:Find:Pt:Chest>Pleural space:Doc:US
C0881887|Guidance for aspiration:Finding:Point in time:Chest>Pleural space:Document:Ultrasound
C0881921|Fem a XRA Runoff W contr IA
C0881921|Femoral artery Fluoroscopic angiogram runoff W contrast IA
C0881921|View runoff^W contrast IA:Find:Pt:Femoral artery:Doc:XR.fluor.angio
C0881921|View runoff^W contrast Intra-arterial:Finding:Point in time:Femoral artery:Document:XR.fluor.angio
C0881932|Gallbladder X-ray 48 hours post contrast PO
C0881932|GB XR 48h p contr PO
C0881932|Views^48H post contrast Oral:Finding:Point in time:Gallbladder:Document:XR
C0881932|Views^48H post contrast PO:Find:Pt:Gallbladder:Doc:XR
C0881955|Petrous bone X-ray
C0881955|Petrous bone XR
C0881955|Views:Finding:Point in time:Petrous bone:Document:XR
C0881955|Views:Find:Pt:Petrous bone:Doc:XR
C0881960|Views^W 201 tl subtraction Tc-99m Intravenous:Finding:Point in time:Parathyroid:Narrative:Radnuc
C0881960|Parathyroid RI W TI201-Tc99mIV
C0881960|Views^W TI-201 subtraction Tc-99m IV:Find:Pt:Parathyroid:Doc:Radnuc
C0881960|Parathyroid Scan W TI-201 subtraction Tc-99m IV
C0881960|Views^W TI-201 subtraction Tc-99m Intravenous:Finding:Point in time:Parathyroid:Document:Radnuc
C0882536|VIEWS^W CONTRAST.XXX INTRA ARTICULAR:FINDING:POINT IN TIME:HIP:NARRATIVE:XR.FLUOR
C0882536|Views^W contrast IS:Find:Pt:Hip:Doc:XR.fluor
C0882536|Hip Fluoroscopy W contrast IS
C0882536|Hip Flr W contr IS
C0882536|Views^W contrast Intrasynovial:Finding:Point in time:Hip:Document:XR.fluor
C0881992|Abd XR AP+AP L-Lat Decub Port
C0881992|Abdomen X-ray AP and AP left lateral-decubitus portable
C0881992|Views AP & AP L-lateral-decubitus portable:Finding:Point in time:Abdomen:Document:XR
C0881992|Views AP & AP L-lateral-decubitus portable:Find:Pt:Abdomen:Doc:XR
C1114479|Brain MRI WO contr
C1114479|Brain MRI WO contrast
C1114479|Multisection^WO contrast:Find:Pt:Brain:Doc:MRI
C1114479|Multisection^WO contrast:Finding:Point in time:Brain:Document:MRI
C1114496|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pelvis:Document:MRI
C1114496|Multisection^WO & W contrast IV:Find:Pt:Pelvis:Doc:MRI
C1114496|Pelvis MRI WO and W contrast IV
C1114496|Pelvis MRI WO+W contr IV
C1114514|Scrotum+Test RI W RNC IV
C1114514|Scrotum and Testicle Scan
C1114514|Views^W radionuclide IV:Find:Pt:Scrotum+Testicle:Doc:Radnuc
C1114514|Views^W radionuclide Intravenous:Finding:Point in time:Scrotum+Testicle:Document:Radnuc
C1114519|Pericardial space US Asp guid
C1114519|US Guidance for aspiration of Pericardial space
C1114519|Guidance for aspiration:Find:Pt:Pericardial space:Doc:US
C1114519|Guidance for aspiration:Finding:Point in time:Pericardial space:Document:Ultrasound
C1114525|Hip US Devel joint assess
C1114525|Hip US developmental joint assessment
C1114525|Multisection^developmental joint assessment:Find:Pt:Hip:Doc:US
C1114525|Multisection^developmental joint assessment:Finding:Point in time:Hip:Document:Ultrasound
C1114548|Chest X-ray AP lateral-decubitus portable
C1114548|Chest XR AP Lat Decub Port
C1114548|View AP lateral-decubitus portable:Finding:Point in time:Chest:Document:XR
C1114548|View AP lateral-decubitus portable:Find:Pt:Chest:Doc:XR
C1114600|Breast - bilateral MRI
C1114600|Brst-Bl MRI
C1114600|Multisection:Find:Pt:Breast.bilateral:Doc:MRI
C1114600|Multisection:Finding:Point in time:Breast.bilateral:Document:MRI
C1114628|Brachial artery Fluoroscopic angiogram W contrast IA
C1114628|Brach a XRA W contr IA
C1114628|Views^W contrast Intra-arterial:Finding:Point in time:Brachial artery:Document:XR.fluor.angio
C1114628|Views^W contrast IA:Find:Pt:Brachial artery:Doc:XR.fluor.angio
C1114646|Renal v XRA W contr IV
C1114646|Renal vein Fluoroscopic angiogram W contrast IV
C1114646|Views^W contrast Intravenous:Finding:Point in time:Renal vein:Document:XR.fluor.angio
C1114646|Views^W contrast IV:Find:Pt:Renal vein:Doc:XR.fluor.angio
C1114646|VIEWS^W CONTRAST.XXX INTRAVENOUS:FINDING:POINT IN TIME:VEIN.RENAL:NARRATIVE:XR.FLUOR.ANGIO
C1114663|Lumbar plexus MRI
C1114663|Multisection:Finding:Point in time:Lumbar plexus:Document:MRI
C1114663|Multisection:Find:Pt:Lumbar plexus:Doc:MRI
C1114672|KD-Bl+Renal ves RI W RNC IV
C1114672|Kidney - bilateral and Renal vessels Scan
C1114672|Views^W radionuclide IV:Find:Pt:Kidney.bilateral+Renal vessels:Doc:Radnuc
C1114672|Views^W radionuclide Intravenous:Finding:Point in time:Kidney.bilateral+Renal vessels:Document:Radnuc
C1114927|Diaphragm Fluoroscopy Motion
C1114927|Diaphragm Flr Motion
C1114927|Motion:Find:Pt:Diaphragm:Doc:XR.fluor
C1114927|Motion:Finding:Point in time:Diaphragm:Document:XR.fluor
C1114471|Periph a XRA Add'l Angpsty W contr IA
C1114471|Peripheral artery Fluoroscopic angiogram Additional angioplasty W contrast IA
C1114471|Angioplasty.additional^W contrast IA:Find:Pt:Peripheral artery:Doc:XR.fluor.angio
C1114471|Angioplasty.additional^W contrast Intra-arterial:Finding:Point in time:Peripheral artery:Document:XR.fluor.angio
C1543481|Sinuses X-ray 3 views and submentovertex
C1543481|Sinuses XR 3V+SMV
C1543481|Views 3 & submentovertex:Find:Pt:Sinuses:Doc:XR
C1543481|Views 3 & submentovertex:Finding:Point in time:Sinuses:Document:XR
C1542849|Scan Guidance for localization of tumor of Breast
C1542849|Brst RI Tum local guid W RNC IV
C1542849|Guidance for localization of tumor^W radionuclide Intravenous:Finding:Point in time:Breast:Document:Radnuc
C1542849|Guidance for localization of tumor^W radionuclide IV:Find:Pt:Breast:Doc:Radnuc
C1543861|Bone Scan delayed
C1543861|Bone RI Delayed W RNC IV
C1543861|Views delayed^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543861|Views delayed^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1542907|RI WB W In-111 Satmb IV
C1542907|Scan whole body W In-111 Satumomab IV
C1542907|Views whole body^W In-111 Satumomab IV:Find:Pt:^Patient:Doc:Radnuc
C1542907|Views whole body^W In-111 Satumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543908|Hrt RI FP+WM Rest+W RNC IV
C1543908|Heart Scan first pass and wall motion at rest and W radionuclide IV
C1543908|Views first pass & wall motion^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543908|Views first pass & wall motion^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543940|Hrt SPECT Gated+WM W RNC IV
C1543940|Heart SPECT gated and wall motion
C1543940|Multisection gated & wall motion^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543940|Multisection gated & wall motion^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543508|Lower extremity vein - left US.doppler
C1543508|LE v-L DOP
C1543508|Multisection:Find:Pt:Lower extremity vein.left:Doc:US.doppler
C1543508|Multisection:Finding:Point in time:Lower extremity vein.left:Document:Ultrasound.doppler
C1543513|Multisection:Finding:Point in time:Carotid artery.right:Narrative:ULTRASOUND.doppler
C1543513|Carot a-R DOP
C1543513|Carotid artery - right US.doppler
C1543513|Multisection:Finding:Point in time:Carotid artery.right:Document:Ultrasound.doppler
C1543513|Multisection:Find:Pt:Carotid artery.right:Doc:US.doppler
C1543526|Gastrointestine US W contrast PO
C1543526|GI US W contr PO
C1543526|Multisection^W contrast PO:Find:Pt:Gastrointestine:Doc:US
C1543526|Multisection^W contrast Oral:Finding:Point in time:Gastrointestine:Document:Ultrasound
C1543566|Femur+Tib-R XR Leg Length
C1543566|Femur - right and Tibia - right X-ray for leg length
C1543566|Views for leg length:Finding:Point in time:Femur.right+Tibia.right:Document:XR
C1543566|Views for leg length:Find:Pt:Femur.right+Tibia.right:Doc:XR
C1543582|Upper extremity artery - right US.doppler
C1543582|UE a-R DOP
C1543582|Multisection:Find:Pt:Upper extremity artery.right:Doc:US.doppler
C1543582|Multisection:Finding:Point in time:Upper extremity artery.right:Document:Ultrasound.doppler
C1526351|Bone density:Mass Aeric:Point in time:Calcaneus:Quantitative:XR.DXA
C1526351|Bone density:MAric:Pt:Calcaneus:Qn:XR.DXA
C1526351|Deprecated Calcaneus DXA Bone density
C1526351|Deprecated Heel DXA BDM
C1543192|Knee XR AP+Lat+Merchants
C1543192|Knee X-ray AP and lateral and Merchants
C1543192|Views AP & lateral & Merchants:Find:Pt:Knee:Doc:XR
C1543192|Views AP & lateral & Merchants:Finding:Point in time:Knee:Document:XR
C1525169|Lower extremity vessels - right MRI angiogram WO contrast
C1525169|LE ves-R MRI.Angio WO contr
C1525169|Multisection^WO contrast:Find:Pt:Lower extremity vessels.right:Doc:MRI.angio
C1525169|Multisection^WO contrast:Finding:Point in time:Lower extremity vessels.right:Document:MRI.angio
C1542864|Breast FFD mammogram screening
C1542864|Brst FFDM Screening
C1542864|Views screening:Find:Pt:Breast:Doc:Mam.FFD
C1542864|Views screening:Finding:Point in time:Breast:Document:Mam.FFD
C1543696|Brain RI Static Ltd W RNC IV
C1543696|Brain Scan static limited
C1543696|Views static limited ^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc
C1543696|Views static limited^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1524264|Should-R XR Grashey+Ax+ Y
C1524264|Shoulder - right X-ray Grashey and axillary and Y
C1524264|Views Grashey & axillary & Y:Finding:Point in time:Shoulder.right:Document:XR
C1524264|Views Grashey & axillary & Y:Find:Pt:Shoulder.right:Doc:XR
C1526772|Views Grashey^WO & W weight:Finding:Point in time:Shoulder.right:Document:XR
C1526772|Shoulder - right X-ray Grashey WO and W weight
C1526772|Views Grashey^WO & W weight:Find:Pt:Shoulder.right:Doc:XR
C1526772|Should-R XR Grashey WO+W Wt
C1526773|Breast implant - right MRI WO contrast
C1526773|Brst implant-R MRI WO contr
C1526773|Multisection^WO contrast:Find:Pt:Breast implant.right:Doc:MRI
C1526773|Multisection^WO contrast:Finding:Point in time:Breast implant.right:Document:MRI
C3484383|Brst RI W RNC IV
C3484383|Breast Scan
C3484383|Views^W radionuclide IV:Find:Pt:Breast:Doc:Radnuc
C3484383|Views^W radionuclide Intravenous:Finding:Point in time:Breast:Document:Radnuc
C1526809|Lower extremity vessels - left Fluoroscopic angiogram W contrast
C1526809|LE ves-L XRA W contr
C1526809|Views^W contrast:Finding:Point in time:Lower extremity vessels.left:Document:XR.fluor.angio
C1526809|Views^W contrast:Find:Pt:Lower extremity vessels.left:Doc:XR.fluor.angio
C1524837|Lower extremity - left CT WO contrast
C1524837|LE-L CT WO contr
C1524837|Multisection^WO contrast:Finding:Point in time:Lower extremity.left:Document:Computerized Tomography
C1524837|Multisection^WO contrast:Find:Pt:Lower extremity.left:Doc:CT
C1525315|Hip - left X-ray Judet
C1525315|Hip-L XR Judet
C1525315|View Judet:Finding:Point in time:Hip.left:Document:XR
C1525315|View Judet:Find:Pt:Hip.left:Doc:XR
C1525197|Orbit-R MRI W contr IV
C1525197|Orbit - right MRI W contrast IV
C1525197|Multisection^W contrast IV:Find:Pt:Orbit.right:Doc:MRI
C1525197|Multisection^W contrast Intravenous:Finding:Point in time:Orbit.right:Document:MRI
C1525221|Head vv MRI.Angio WO+W contr IV
C1525221|Multisection^WO & W contrast IV:Find:Pt:Head veins:Doc:MRI.angio
C1525221|Head veins MRI angiogram WO and W contrast IV
C1525221|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head veins:Document:MRI.angio
C1525256|Pelvis ves MRI.Angio WO contr
C1525256|Pelvis vessels MRI angiogram WO contrast
C1525256|Multisection^WO contrast:Find:Pt:Pelvis vessels:Doc:MRI.angio
C1525256|Multisection^WO contrast:Finding:Point in time:Pelvis vessels:Document:MRI.angio
C1525259|Mastoid XR Ltd
C1525259|Mastoid X-ray limited
C1525259|Views limited:Finding:Point in time:Mastoid:Document:XR
C1525259|Views limited:Find:Pt:Mastoid:Doc:XR
C1525268|Brain MRI Bx Str Guid
C1525268|MRI Guidance for stereotactic biopsy of Brain
C1525268|Guidance for stereotactic biopsy:Finding:Point in time:Brain:Document:MRI
C1525268|Guidance for stereotactic biopsy:Find:Pt:Brain:Doc:MRI
C1525331|Knee-Bl XR Lat Hyperext
C1525331|Knee - bilateral X-ray lateral hyperextension
C1525331|View lateral hyperextension:Finding:Point in time:Knee.bilateral:Document:XR
C1525331|View lateral hyperextension:Find:Pt:Knee.bilateral:Doc:XR
C1525332|Knee-L XR Lat Hyperext
C1525332|Knee - left X-ray lateral hyperextension
C1525332|View lateral hyperextension:Finding:Point in time:Knee.left:Document:XR
C1525332|View lateral hyperextension:Find:Pt:Knee.left:Doc:XR
C1525343|L-spine XR R-Obl
C1525343|View R-oblique:Find:Pt:Spine.lumbar:Doc:XR
C1525343|View R-oblique:Finding:Point in time:Spine.lumbar:Document:XR
C1525343|Lumbar spine X-ray right oblique
C1525488|Hip XR AP+Lat Xtable port
C1525488|Hip X-ray AP and lateral crosstable portable
C1525488|Views AP & lateral crosstable portable:Find:Pt:Hip:Doc:XR
C1525488|Views AP & lateral crosstable portable:Finding:Point in time:Hip:Document:XR
C1525541|Hand-Bl XR PA+Lat+Ball Catcher
C1525541|Hand - bilateral X-ray PA and lateral and Ball Catcher
C1525541|Views PA & lateral & Ball Catcher:Find:Pt:Hand.bilateral:Doc:XR
C1525541|Views PA & lateral & Ball Catcher:Finding:Point in time:Hand.bilateral:Document:XR
C1525631|Sinus tract CT W contrast intra sinus tract
C1525631|Sinus tr CT W contr intra ST
C1525631|Multisection^W contrast intra sinus tract:Finding:Point in time:Sinus tract:Document:Computerized Tomography
C1525631|Multisection^W contrast intra sinus tract:Find:Pt:Sinus tract:Doc:CT
C1525668|Temporomandibular joint - left MRI WO contrast
C1525668|TMJ-L MRI WO contr
C1525668|Multisection^WO contrast:Finding:Point in time:Temporomandibular joint.left:Document:MRI
C1525668|Multisection^WO contrast:Find:Pt:Temporomandibular joint.left:Doc:MRI
C1525674|Abd+Fetus XR 1V for FTA
C1525674|Abdomen and Fetus X-ray View for fetal age
C1525674|View for fetal age:Finding:Point in time:Abdomen+Fetus:Document:XR
C1525674|View for fetal age:Find:Pt:Abdomen+Fetus:Doc:XR
C1525798|Fluoroscopy Guidance for injection of Tendon
C1525798|Tendon Flr Inj guid
C1525798|Guidance for injection:Find:Pt:XXX tendon:Doc:XR.fluor
C1525798|Guidance for injection:Finding:Point in time:To be specified in another part of the message tendon:Document:XR.fluor
C1525843|Wrist-Bl XR PA+Lat
C1525843|Wrist - bilateral X-ray PA and lateral
C1525843|Views PA & lateral:Find:Pt:Wrist.bilateral:Doc:XR
C1525843|Views PA & lateral:Finding:Point in time:Wrist.bilateral:Document:XR
C1524142|Ext lymphr-L Flr W contr IL
C1524142|Extremity lymphatics - left Fluoroscopy W contrast intra lymphatic
C1524142|Views^W contrast intra lymphatic:Finding:Point in time:Extremity lymphatics.left:Document:XR.fluor
C1524142|Views^W contrast intra lymphatic:Find:Pt:Extremity lymphatics.left:Doc:XR.fluor
C1525892|Optic foramen XR 4V
C1525892|Optic foramen X-ray 4 views
C1525892|Views 4:Find:Pt:Optic foramen:Doc:XR
C1525892|Views 4:Finding:Point in time:Optic foramen:Document:XR
C1525981|Ankle - right X-ray 3 views
C1525981|Ankle-R XR 3V
C1525981|Views 3:Find:Pt:Ankle.right:Doc:XR
C1525981|Views 3:Finding:Point in time:Ankle.right:Document:XR
C1525987|Ankle - right X-ray Mortise W manual stress
C1525987|Ankle-R XR Mortise W Stress
C1525987|View Mortise^W manual stress:Find:Pt:Ankle.right:Doc:XR
C1525987|View Mortise^W manual stress:Finding:Point in time:Ankle.right:Document:XR
C1525988|Ankle - right X-ray 2 views W manual stress
C1525988|Ankle-R XR 2V W Stress
C1525988|Views 2^W manual stress:Finding:Point in time:Ankle.right:Document:XR
C1525988|Views 2^W manual stress:Find:Pt:Ankle.right:Doc:XR
C1526141|Shoulder X-ray axillary
C1526141|Should XR Ax
C1526141|View axillary:Find:Pt:Shoulder:Doc:XR
C1526141|View axillary:Finding:Point in time:Shoulder:Document:XR
C1526175|Tib+Fib XR 2V
C1526175|Tibia and Fibula X-ray 2 views
C1526175|Views 2:Find:Pt:Tibia+Fibula:Doc:XR
C1526175|Views 2:Finding:Point in time:Tibia+Fibula:Document:XR
C1526187|T-spine XR 4V
C1526187|Views 4:Find:Pt:Spine.thoracic:Doc:XR
C1526187|Views 4:Finding:Point in time:Spine.thoracic:Document:XR
C1526187|Thoracic spine X-ray 4 views
C1526251|Elbow - bilateral X-ray radial head capitellar
C1526251|Elbow-Bl XR Radial Head Capitellar
C1526251|View radial head capitellar:Finding:Point in time:Elbow.bilateral:Document:XR
C1526251|View radial head capitellar:Find:Pt:Elbow.bilateral:Doc:XR
C1525132|Elbow-R XR Radial Head Capitellar
C1525132|Elbow - right X-ray radial head capitellar
C1525132|View radial head capitellar:Find:Pt:Elbow.right:Doc:XR
C1525132|View radial head capitellar:Finding:Point in time:Elbow.right:Document:XR
C1526258|US Guidance for fine needle aspiration of Prostate
C1526258|Prostate US FNA Asp
C1526258|Guidance for aspiration.fine needle:Find:Pt:Prostate:Doc:US
C1526258|Guidance for aspiration.fine needle:Finding:Point in time:Prostate:Document:Ultrasound
C1526260|Thyroid US FNA Asp
C1526260|US Guidance for fine needle aspiration of Thyroid
C1526260|Guidance for aspiration.fine needle:Find:Pt:Thyroid:Doc:US
C1526260|Guidance for aspiration.fine needle:Finding:Point in time:Thyroid:Document:Ultrasound
C1526265|US Guidance for core needle biopsy of Unspecified body region
C1526265|XXX US Bx CN guid
C1526265|Guidance for biopsy.core needle:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1526265|Guidance for biopsy.core needle:Find:Pt:XXX:Doc:US
C1526270|US Guidance for needle biopsy of Chest
C1526270|Chest US Bx needle guid
C1526270|Guidance for biopsy.needle:Find:Pt:Chest:Doc:US
C1526270|Guidance for biopsy.needle:Finding:Point in time:Chest:Document:Ultrasound
C1526297|Chest X-ray right anterior oblique
C1526297|Chest XR R-Ant Obl
C1526297|View R-anterior oblique:Find:Pt:Chest:Doc:XR
C1526297|View R-anterior oblique:Finding:Point in time:Chest:Document:XR
C1524858|Forearm-L CT WO contr
C1524858|Forearm - left CT WO contrast
C1524858|Multisection^WO contrast:Finding:Point in time:Forearm.left:Document:Computerized Tomography
C1524858|Multisection^WO contrast:Find:Pt:Forearm.left:Doc:CT
C1524870|Hip - bilateral CT WO contrast
C1524870|Hip-Bl CT WO contr
C1524870|Multisection^WO contrast:Find:Pt:Hip.bilateral:Doc:CT
C1524870|Multisection^WO contrast:Finding:Point in time:Hip.bilateral:Document:Computerized Tomography
C1524889|Kidney - bilateral MRI WO contrast
C1524889|Multisection^WO contrast:Finding:Point in time:Kidney.bilateral:Document:MRI
C1524889|Multisection^WO contrast:Find:Pt:Kidney.bilateral:Doc:MRI
C1524889|Kdny-Bl MRI WO contr
C1524515|UE-R MRI W contr IV
C1524515|Upper extremity - right MRI W contrast IV
C1524515|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.right:Document:MRI
C1524515|Multisection^W contrast IV:Find:Pt:Upper extremity.right:Doc:MRI
C1524921|Inferior vena cava MRI WO contrast
C1524921|IVC MRI WO contr
C1524921|Multisection^WO contrast:Finding:Point in time:Vena cava.inferior:Document:MRI
C1524921|Multisection^WO contrast:Find:Pt:Vena cava.inferior:Doc:MRI
C1524550|UE joint MRI W contr IV
C1524550|Multisection^W contrast IV:Find:Pt:Upper extremity.joint:Doc:MRI
C1524550|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.joint:Document:MRI
C1524550|Upper extremity.joint MRI W contrast IV
C1524573|TO MRI W contr IV
C1524573|Thoracic outlet MRI W contrast IV
C1524573|Multisection^W contrast Intravenous:Finding:Point in time:Thoracic outlet:Document:MRI
C1524573|Multisection^W contrast IV:Find:Pt:Thoracic outlet:Doc:MRI
C1524580|Sacrum MRI W contr IV
C1524580|Sacrum MRI W contrast IV
C1524580|Multisection^W contrast Intravenous:Finding:Point in time:Sacrum:Document:MRI
C1524580|Multisection^W contrast IV:Find:Pt:Sacrum:Doc:MRI
C1524295|CT Guidance for biopsy of Lower extremity
C1524295|LE CT Bx guid
C1524295|Guidance for biopsy:Finding:Point in time:Lower extremity:Document:Computerized Tomography
C1524295|Guidance for biopsy:Find:Pt:Lower extremity:Doc:CT
C1524593|Lower leg MRI W contr IV
C1524593|Lower leg MRI W contrast IV
C1524593|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg:Document:MRI
C1524593|Multisection^W contrast IV:Find:Pt:Lower leg:Doc:MRI
C1524611|Elbow CT WO+W contr IV
C1524611|Multisection^WO & W contrast Intravenous:Finding:Point in time:Elbow:Document:Computerized Tomography
C1524611|Elbow CT WO and W contrast IV
C1524611|Multisection^WO & W contrast IV:Find:Pt:Elbow:Doc:CT
C1524314|Appendix CT Drain guid
C1524314|CT Guidance for drainage of Appendix
C1524314|Guidance for drainage:Find:Pt:Abdomen+Pelvis>Appendix:Doc:CT
C1524314|Guidance for drainage:Finding:Point in time:Abdomen+Pelvis>Appendix:Document:Computerized Tomography
C1524326|Fluoroscopy Guidance for injection of Sacroiliac Joint
C1524326|SIJ Flr Inj guid
C1524326|Guidance for injection:Finding:Point in time:Sacroiliac joint:Document:XR.fluor
C1524326|Guidance for injection:Find:Pt:Sacroiliac joint:Doc:XR.fluor
C1524644|Face XR 4V
C1524644|Facial bones X-ray 4 views
C1524644|Views 4:Find:Pt:Facial bones:Doc:XR
C1524644|Views 4:Finding:Point in time:Facial bones:Document:XR
C1524991|Chest X-ray 2 views
C1524991|Chest XR 2V
C1524991|Views 2:Finding:Point in time:Chest:Document:XR
C1524991|Views 2:Find:Pt:Chest:Doc:XR
C1524160|Views 2:Find:Pt:Calcaneus.left:Doc:XR
C1524160|Views 2:Finding:Point in time:Calcaneus.left:Document:XR
C1524160|Deprecated Heel-L XR 2V
C1524160|Deprecated Calcaneus - left X-ray 2 views
C1524378|Femur CT
C1524378|Multisection:Find:Pt:Femur:Doc:CT
C1524378|Multisection:Finding:Point in time:Femur:Document:Computerized Tomography
C1525057|Tib+Fib-L XR AP+Lat
C1525057|Tibia - left and Fibula - left X-ray AP and lateral
C1525057|Views AP & lateral:Finding:Point in time:Tibia.left+Fibula.left:Document:XR
C1525057|Views AP & lateral:Find:Pt:Tibia.left+Fibula.left:Doc:XR
C1525060|Ankle-L XR AP+Lat+Obl
C1525060|Ankle - left X-ray AP and lateral and oblique
C1525060|Views AP & lateral & oblique:Finding:Point in time:Ankle.left:Document:XR
C1525060|Views AP & lateral & oblique:Find:Pt:Ankle.left:Doc:XR
C1524402|Multisection:Finding:Point in time:Calcaneus:Document:XR.tomo
C1524402|Multisection:Find:Pt:Calcaneus:Doc:XR.tomo
C1524402|Deprecated Heel XRTomo
C1524402|Deprecated Calcaneus X-ray tomograph
C1524422|Kidney - bilateral MRI
C1524422|Multisection:Find:Pt:Kidney.bilateral:Doc:MRI
C1524422|Multisection:Finding:Point in time:Kidney.bilateral:Document:MRI
C1524422|Kdny-Bl MRI
C1524426|Knee-Bl XRTomo
C1524426|Knee - bilateral X-ray tomograph
C1524426|Multisection:Find:Pt:Knee.bilateral:Doc:XR.tomo
C1524426|Multisection:Finding:Point in time:Knee.bilateral:Document:XR.tomo
C1524769|Mandible CT WO+W contr IV
C1524769|Multisection^WO & W contrast IV:Find:Pt:Mandible:Doc:CT
C1524769|Mandible CT WO and W contrast IV
C1524769|Multisection^WO & W contrast Intravenous:Finding:Point in time:Mandible:Document:Computerized Tomography
C1524780|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder:Document:Computerized Tomography
C1524780|Shoulder CT WO and W contrast IV
C1524780|Should CT WO+W contr IV
C1524780|Multisection^WO & W contrast IV:Find:Pt:Shoulder:Doc:CT
C1524782|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder.right:Document:Computerized Tomography
C1524782|Multisection^WO & W contrast IV:Find:Pt:Shoulder.right:Doc:CT
C1524782|Shoulder - right CT WO and W contrast IV
C1524782|Should-R CT WO+W contr IV
C1524804|Multisection^WO & W contrast IV:Find:Pt:Vena cava.superior:Doc:MRI
C1524804|Superior vena cava MRI WO and W contrast IV
C1524804|Multisection^WO & W contrast Intravenous:Finding:Point in time:Vena cava.superior:Document:MRI
C1524804|SVC MRI WO+W contr IV
C1524670|Knee-Bl XR AP+Lat+Obl
C1524670|Knee - bilateral X-ray AP and lateral and oblique
C1524670|Views AP & lateral & oblique:Finding:Point in time:Knee.bilateral:Document:XR
C1524670|Views AP & lateral & oblique:Find:Pt:Knee.bilateral:Doc:XR
C1830186|Thyroid US Bx CN guid
C1830186|US Guidance for core needle biopsy of Thyroid
C1830186|Guidance for biopsy.core needle:Finding:Point in time:Thyroid:Document:Ultrasound
C1830186|Guidance for biopsy.core needle:Find:Pt:Thyroid:Doc:US
C1830230|Pelvis CT W red contr vol IV
C1830230|Pelvis CT W reduced contrast volume IV
C1830230|Multisection^W reduced contrast volume IV:Find:Pt:Pelvis:Doc:CT
C1830230|Multisection^W reduced contrast volume Intravenous:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1830085|X-ray Guidance for change of percutaneous tube in Unspecified body region-- W contrast
C1830085|XXX XR PC tube change guid W contr
C1830085|Guidance for change of percutaneous tube^W contrast:Find:Pt:XXX:Doc:XR
C1830085|Guidance for change of percutaneous tube^W contrast:Finding:Point in time:To be specified in another part of the message:Document:XR
C1830086|BDs Flr PC drain guid
C1830086|Fluoroscopy Guidance for percutaneous drainage of Biliary ducts
C1830086|Guidance for percutaneous drainage:Finding:Point in time:Biliary ducts:Document:XR.fluor
C1830086|Guidance for percutaneous drainage:Find:Pt:Biliary ducts:Doc:XR.fluor
C1830090|Views^W contrast antegrade:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C1830090|Kidney - bilateral Fluoroscopy W contrast antegrade
C1830090|Views^W contrast antegrade:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C1830090|Kdny-Bl Flr W contr Ante
C1830092|Knee-Bl XR PA Stand+W Flx
C1830092|Knee - bilateral X-ray PA standing and W flexion
C1830092|Views PA^standing & W flexion:Find:Pt:Knee.bilateral:Doc:XR
C1830092|Views PA^standing & W flexion:Finding:Point in time:Knee.bilateral:Document:XR
C1830271|Hand ves DOP
C1830271|Hand vessels US.doppler
C1830271|Multisection:Finding:Point in time:Hand vessels:Document:Ultrasound.doppler
C1830271|Multisection:Find:Pt:Hand vessels:Doc:US.doppler
C1715391|Multisection:Find:Pt:Colon:Doc:CT
C1715391|Deprecated Colon CT
C1715391|Multisection:Finding:Point in time:Colon:Document:Computerized Tomography
C1715418|Brain RI Static W Tc99mBicisate IV
C1715418|Brain Scan static W Tc-99m bicisate IV
C1715418|Views static^W Tc-99m bicisate Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1715418|Views static^W Tc-99m bicisate IV:Find:Pt:Brain:Doc:Radnuc
C1715425|US Guidance for fine needle aspiration of Pancreas
C1715425|Pancreas US FNA Asp
C1715425|Guidance for aspiration.fine needle:Finding:Point in time:Pancreas:Document:Ultrasound
C1715425|Guidance for aspiration.fine needle:Find:Pt:Pancreas:Doc:US
C1715497|Ribs-Ul+chest XR GE 3V+PA Chst Port
C1715497|Ribs - unilateral and Chest X-ray Ge 3 and PA Chest Portable views
C1715497|Views GE 3 & PA chest portable:Finding:Point in time:Ribs.unilateral+Chest:Document:XR
C1715497|Views GE 3 & PA chest portable:Find:Pt:Ribs.unilateral+Chest:Doc:XR
C1644645|Abdomen CT
C1644645|Abd CT
C1644645|Multisection:Finding:Point in time:Abdomen:Narrative:Computerized Tomography
C1644645|Multisection:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1644645|Multisection:Find:Pt:Abdomen:Doc:CT
C1649483|Wrist - left X-ray portable
C1649483|Wrist-L XR port
C1649483|Views portable:Finding:Point in time:Wrist.left:Document:XR
C1649483|Views portable:Find:Pt:Wrist.left:Doc:XR
C1627420|Brain MRI cine for CSF flow
C1627420|Multisection cine for CSF flow:Find:Pt:Brain:Doc:MRI
C1627420|Multisection cine for CSF flow:Finding:Point in time:Brain:Document:MRI
C1627371|Wrist X-ray scaphoid single view
C1627371|Wrist XR Scaphoid 1V
C1627371|View scaphoid:Finding:Point in time:Wrist:Document:XR
C1627371|View scaphoid:Find:Pt:Wrist:Doc:XR
C1717224|Kidney XR in Surg W contr retro
C1717224|Views^during surgery W contrast retrograde:Find:Pt:Kidney:Doc:XR
C1717224|Kidney X-ray during surgery W contrast retrograde
C1717224|Views^during surgery W contrast retrograde:Finding:Point in time:Kidney:Document:XR
C1714917|Wrist Ves-R MRI.Angio WO contr
C1714917|Wrist vessels - right MRI angiogram WO contrast
C1714917|Multisection^WO contrast:Finding:Point in time:Wrist vessels.right:Document:MRI.angio
C1714917|Multisection^WO contrast:Find:Pt:Wrist vessels.right:Doc:MRI.angio
C1714932|Deprecated Mandible-L XR 4V
C1714932|Deprecated Mandible - left X-ray 4 views
C1714932|Views 4:Find:Pt:Mandible.left:Doc:XR
C1714932|Views 4:Finding:Point in time:Mandible.left:Document:XR
C1714958|Guidance for biopsy.needle:Find:Pt:Soft bone:Doc:CT
C1714958|Deprecated Soft Bone CT Bx needle guid
C1714958|Guidance for biopsy.needle:Finding:Point in time:Soft bone:Document:Computerized Tomography
C1714958|Deprecated CT Guidance for needle biopsy of Soft bone
C1717269|Lung Scan perfusion quantitative
C1717269|Lung RI PF Qn W RNC IV
C1717269|Views perfusion quantitative^W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1717269|Views perfusion quantitative^W radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1715028|Lung RI Qn W RNC IV
C1715028|Lung Scan quantitative
C1715028|Views quantitative^W radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1715028|Views quantitative^W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1715030|Hrt SPECT PF Ql Rest+W RNC IV
C1715030|Heart SPECT perfusion qualitative at rest and W radionuclide IV
C1715030|Multisection perfusion qualitative^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1715030|Multisection perfusion qualitative^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1714496|Renal ves SPECT Flow W Tc99mGHA IV
C1714496|Renal vessels SPECT flow W Tc-99m glucoheptonate IV
C1714496|Multisection flow^W Tc-99m glucoheptonate IV:Find:Pt:Renal vessels:Doc:Radnuc.SPECT
C1714496|Multisection flow^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Renal vessels:Document:Radnuc.SPECT
C1715098|Kidney CT WO contr
C1715098|Kidney CT WO contrast
C1715098|Multisection^WO contrast:Find:Pt:Kidney:Doc:CT
C1715098|Multisection^WO contrast:Finding:Point in time:Kidney:Document:Computerized Tomography
C1715104|Chest X-ray AP supine portable
C1715104|Chest XR AP supine port
C1715104|View AP supine portable:Find:Pt:Chest:Doc:XR
C1715104|View AP supine portable:Finding:Point in time:Chest:Document:XR
C1715114|Tube Flr for Pat W contr via tb
C1715114|Tube Fluoroscopy for patency W contrast via tube
C1715114|Views for patency^W contrast via tube:Find:Pt:XXX tube:Doc:XR.fluor
C1715114|Views for patency^W contrast via tube:Finding:Point in time:To be specified in another part of the message tube:Document:XR.fluor
C1633470|ST XRTomo
C1633470|Sella turcica X-ray tomograph
C1633470|Multisection:Find:Pt:Sella turcica:Doc:XR.tomo
C1633470|Multisection:Finding:Point in time:Sella turcica:Document:XR.tomo
C1623094|Deprecated Neck XR Lat
C1623094|Deprecated Neck X-ray lateral
C1623094|View lateral:Find:Pt:Neck:Nar:XR
C1623094|View lateral:Finding:Point in time:Neck:Narrative:XR
C1644657|Deprecated Views^W water soluble contrast Rectal:Finding:Point in time:Colon:Narrative:XR.fluor
C1644657|Views^W water soluble contrast PR:Find:Pt:Colon:Nar:XR.fluor
C1644657|Deprecated Colon X-ray fluoroscopy W water soluble contrast PR
C1644657|Deprecated Colon Flr W H2O sol contr PR
C1644657|Views^W water soluble contrast Rectal:Finding:Point in time:Colon:Narrative:XR.fluor
C1638280|UGI+GB Flr W contr PO
C1638280|Gastrointestine upper and Gallbladder Fluoroscopy W contrast PO
C1638280|View^W contrast PO:Find:Pt:Gastrointestine.upper+Gallbladder:Doc:XR.fluor
C1638280|View^W contrast Oral:Finding:Point in time:Gastrointestine.upper+Gallbladder:Document:XR.fluor
C1639907|Vessels Fluoroscopic angiogram W contrast IA
C1639907|Vesl XRA W contr IA
C1639907|Views^W contrast Intra-arterial:Finding:Point in time:Vessels:Document:XR.fluor.angio
C1639907|Views^W contrast IA:Find:Pt:Vessels:Doc:XR.fluor.angio
C1627301|Deprecated Views portable:Finding:Point in time:Tibia.right+Fibula.right:Narrative:XR
C1627301|Deprecated Tib+Fib-R XR port
C1627301|Views portable:Find:Pt:Tibia.right+Fibula.right:Nar:XR
C1627301|Deprecated Tibia Right & Fibula Right X-ray
C1627301|Views portable:Finding:Point in time:Tibia.right+Fibula.right:Narrative:XR
C1649480|Chest XR in Surg
C1649480|Chest X-ray during surgery
C1649480|View^during surgery:Finding:Point in time:Chest:Document:XR
C1649480|View^during surgery:Find:Pt:Chest:Doc:XR
C1644665|Kidney SPECT W RNC IV
C1644665|Kidney SPECT
C1644665|Multisection^W radionuclide IV:Find:Pt:Kidney:Doc:Radnuc.SPECT
C1644665|Multisection^W radionuclide Intravenous:Finding:Point in time:Kidney:Document:Radnuc.SPECT
C1623597|CT Guidance for localization of placenta of Uterus
C1623597|Uterus CT Placenta local guid
C1623597|Guidance for localization of placenta:Find:Pt:Uterus:Doc:CT
C1623597|Guidance for localization of placenta:Finding:Point in time:Uterus:Document:Computerized Tomography
C1623599|Hrt US Ltd
C1623599|Heart US limited
C1623599|Multisection limited:Finding:Point in time:Heart:Document:Ultrasound
C1623599|Multisection limited:Find:Pt:Heart:Doc:US
C1624135|RI WB W In-111 WBC IV
C1624135|Scan whole body W In-111 tagged WBC IV
C1624135|Views whole body^W In-111 tagged WBC Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1624135|Views whole body^W In-111 tagged WBC IV:Find:Pt:^Patient:Doc:Radnuc
C1978438|Wrist+Hand-R XR
C1978438|Wrist - right and Hand - right X-ray
C1978438|Views:Finding:Point in time:Wrist.right+Hand.right:Document:XR
C1978438|Views:Find:Pt:Wrist.right+Hand.right:Doc:XR
C1977262|Fem a XRA Runoff WO+W contr IA
C1977262|View runoff^WO & W contrast IA:Find:Pt:Femoral artery:Doc:XR.fluor.angio
C1977262|View runoff^WO & W contrast Intra-arterial:Finding:Point in time:Femoral artery:Document:XR.fluor.angio
C1977262|Femoral artery Fluoroscopic angiogram runoff WO and W contrast IA
C1953942|L-spine MRI W contr IT
C1953942|Multisection^W contrast Intrathecal:Finding:Point in time:Spine.lumbar:Document:MRI
C1953942|Multisection^W contrast IT:Find:Pt:Spine.lumbar:Doc:MRI
C1953942|Lumbar spine MRI W contrast IT
C1953992|Ribs-R+Chest XR GE 3V+PA Chst
C1953992|Ribs - right and Chest X-ray GE 3 and PA Chest views
C1953992|Views GE 3 & PA chest:Find:Pt:Ribs.right+Chest:Doc:XR
C1953992|Views GE 3 & PA chest:Finding:Point in time:Ribs.right+Chest:Document:XR
C1952653|Skull X-ray GE 4 views
C1952653|Skull XR GE 4V
C1952653|Views GE 4:Finding:Point in time:Skull:Document:XR
C1952653|Views GE 4:Find:Pt:Skull:Doc:XR
C3169529|Extr-L US Ltd
C3169529|Extremity - left US limited
C3169529|Multisection limited:Find:Pt:Extremity.left:Doc:US
C3169529|Multisection limited:Finding:Point in time:Extremity.left:Document:Ultrasound
C3262936|Kidney - right CT
C3262936|Kidney-R CT
C3262936|Multisection:Finding:Point in time:Kidney.right:Document:Computerized Tomography
C3262936|Multisection:Find:Pt:Kidney.right:Doc:CT
C3262942|TA CT.Angio WO contr
C3262942|Multisection^WO contrast:Finding:Point in time:Chest>Aorta.thoracic:Document:Computerized Tomography.angio
C3262942|Multisection^WO contrast:Find:Pt:Chest>Aorta.thoracic:Doc:CT.angio
C3262942|Thoracic Aorta CT angiogram WO contrast
C3263006|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.bilateral:Document:MRI
C3263006|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.bilateral:Doc:MRI
C3263006|Upper extremity - bilateral MRI WO and W contrast IV
C3263006|UE-Bl MRI WO+W contr IV
C3263016|Finger MRI WO contrast
C3263016|Finger MRI WO contr
C3263016|Multisection^WO contrast:Finding:Point in time:Finger:Document:MRI
C3263016|Multisection^WO contrast:Find:Pt:Finger:Doc:MRI
C3263026|MRI Guidance for biopsy of Breast - right
C3263026|Brst-R MRI Bx guid
C3263026|Guidance for biopsy:Find:Pt:Breast.right:Doc:MRI
C3263026|Guidance for biopsy:Finding:Point in time:Breast.right:Document:MRI
C3263037|Abd Flr Bx needle guid
C3263037|Fluoroscopy Guidance for needle biopsy of Abdomen
C3263037|Guidance for biopsy.needle:Find:Pt:Abdomen:Doc:XR.fluor
C3263037|Guidance for biopsy.needle:Finding:Point in time:Abdomen:Document:XR.fluor
C3263054|Fluoroscopy Guidance for percutaneous drainage of abscess of Abdomen
C3263054|Abd Flr PC Abscess Drain guid
C3263054|Guidance for percutaneous drainage of abscess:Find:Pt:Abdomen:Doc:XR.fluor
C3263054|Guidance for percutaneous drainage of abscess:Finding:Point in time:Abdomen:Document:XR.fluor
C3263055|Fluoroscopy Guidance for percutaneous drainage of abscess of Appendix
C3263055|Appendix Flr PC Abscess Drain guid
C3263055|Guidance for percutaneous drainage of abscess:Finding:Point in time:Appendix:Document:XR.fluor
C3263055|Guidance for percutaneous drainage of abscess:Find:Pt:Appendix:Doc:XR.fluor
C3261711|Ab Ao US
C3261711|Aorta abdominal US
C3261711|Multisection:Find:Pt:Aorta.abdominal:Doc:US
C3261711|Multisection:Finding:Point in time:Aorta.abdominal:Document:Ultrasound
C3261713|US Guidance for aspiration of Breast - bilateral
C3261713|Brst-Bl US Asp guid
C3261713|Guidance for aspiration:Find:Pt:Breast.bilateral:Doc:US
C3261713|Guidance for aspiration:Finding:Point in time:Breast.bilateral:Document:Ultrasound
C3263103|Wrist X-ray ulnar deviation and radial deviation
C3263103|Wrist XR Ulnar+Radial Deviation
C3263103|Views ulnar deviation & radial deviation:Find:Pt:Wrist:Doc:XR
C3263103|Views ulnar deviation & radial deviation:Finding:Point in time:Wrist:Document:XR
C0942185|Brst-L Mam Screening
C0942185|Breast - left Mammogram screening
C0942185|Views screening:Finding:Point in time:Breast.left:Document:Mam
C0942185|Views screening:Find:Pt:Breast.left:Doc:Mam
C0942270|Multisection:Finding:Point in time:Thigh.right:Narrative:MRI
C0942270|Thigh - right MRI
C0942270|Thigh-R MRI
C0942270|Multisection:Finding:Point in time:Thigh.right:Document:MRI
C0942270|Multisection:Find:Pt:Thigh.right:Doc:MRI
C0945330|Hip-L US
C0945330|Hip - left US
C0945330|Multisection:Finding:Point in time:Hip.left:Document:Ultrasound
C0945330|Multisection:Find:Pt:Hip.left:Doc:US
C0942247|Hip - right US
C0942247|Hip-R US
C0942247|Multisection:Finding:Point in time:Hip.right:Document:Ultrasound
C0942247|Multisection:Find:Pt:Hip.right:Doc:US
C0942361|Shoulder - bilateral X-ray 3 views
C0942361|Should-Bl XR 3V
C0942361|Views 3:Finding:Point in time:Shoulder.bilateral:Document:XR
C0942361|Views 3:Find:Pt:Shoulder.bilateral:Doc:XR
C0942375|Patella - right X-ray 2 views
C0942375|Patella-R XR 2V
C0942375|Views 2:Finding:Point in time:Patella.right:Document:XR
C0942375|Views 2:Find:Pt:Patella.right:Doc:XR
C0882037|Neck XR Lat
C0882037|Neck X-ray lateral
C0882037|View lateral:Find:Pt:Neck:Doc:XR
C0882037|View lateral:Finding:Point in time:Neck:Document:XR
C0882544|Pelvis CT W contr IV
C0882544|Pelvis CT W contrast IV
C0882544|Multisection^W contrast Intravenous:Finding:Point in time:Pelvis:Document:Computerized Tomography
C0882544|Multisection^W contrast IV:Find:Pt:Pelvis:Doc:CT
C0882093|Views^W contrast IS:Find:Pt:Shoulder:Doc:XR.fluor
C0882093|Views^W contrast Intrasynovial:Finding:Point in time:Shoulder:Document:XR.fluor
C0882093|Should Flr W contr IS
C0882093|Shoulder Fluoroscopy W contrast IS
C0882111|T+L-spine XR Scoli
C0882111|Spine Thoracic and Lumbar X-ray scoliosis
C0882111|Views scoliosis:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C0882111|Views scoliosis:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C0882121|C-spine XR Lat
C0882121|View lateral:Find:Pt:Spine.cervical:Doc:XR
C0882121|View lateral:Finding:Point in time:Spine.cervical:Document:XR
C0882121|Cervical spine X-ray lateral
C0882142|T-spine MRI W contr IV
C0882142|Multisection^W contrast IV:Find:Pt:Spine.thoracic:Doc:MRI
C0882142|Multisection^W contrast Intravenous:Finding:Point in time:Spine.thoracic:Document:MRI
C0882142|Thoracic spine MRI W contrast IV
C0882159|TMJ MRI
C0882159|Temporomandibular joint MRI
C0882159|Multisection:Finding:Point in time:Temporomandibular joint:Document:MRI
C0882159|Multisection:Find:Pt:Temporomandibular joint:Doc:MRI
C0882165|Views:Finding:Point in time:Thumb:Narrative:XR
C0882165|Thumb X-ray
C0882165|Thumb XR
C0882165|Views:Finding:Point in time:Thumb:Document:XR
C0882165|Views:Find:Pt:Thumb:Doc:XR
C0882172|Upper GI tract Replacement of percutaneous gastrojejunostomy
C0882172|Upr GI Tract Replac of PGJ
C0882172|Replacement of percutaneous gastrojejunostomy:Find:Pt:Upper GI tract:Doc
C0882172|Replacement of percutaneous gastrojejunostomy:Finding:Point in time:Upper GI tract:Document
C0882181|VC XRA W contr IV
C0882181|Vena cava Fluoroscopic angiogram W contrast IV
C0882181|Views^W contrast Intravenous:Finding:Point in time:Vena cava:Document:XR.fluor.angio
C0882181|Views^W contrast IV:Find:Pt:Vena cava:Doc:XR.fluor.angio
C0882185|Fluoroscopic angiogram Guidance for placement of catheter for vasoconstrictor infusion in Vessels
C0882185|Vesl XRA Cath plac guidfor VC inf
C0882185|Guidance for placement of catheter for vasoconstrictor infusion:Find:Pt:Vessels:Doc:XR.fluor.angio
C0882185|Guidance for placement of catheter for vasoconstrictor infusion:Finding:Point in time:Vessels:Document:XR.fluor.angio
C0882205|Multisection sagittal & coronal disarticulation:Find:Pt:XXX:Doc:CT.3D
C0882205|Multisection sagittal & coronal disarticulation:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography.3D
C0882205|Deprecated Unspecified body region CT 3D sagittal and coronal disarticulation
C0882205|Deprecated XXX CT.3D Sagittal+Coronal di
C0942109|Knee - bilateral Scan
C0942109|Knee-Bl RI W RNC IV
C0942109|Views^W radionuclide IV:Find:Pt:Knee.bilateral:Doc:Radnuc
C0942109|Views^W radionuclide Intravenous:Finding:Point in time:Knee.bilateral:Document:Radnuc
C0942131|Lower extremity - left X-ray
C0942131|LE-L XR
C0942131|Views:Finding:Point in time:Lower extremity.left:Document:XR
C0942131|Views:Find:Pt:Lower extremity.left:Doc:XR
C0881775|Abd ves MRI.Angio W contr IV
C0881775|Abdominal vessels MRI angiogram W contrast IV
C0881775|Multisection^W contrast Intravenous:Finding:Point in time:Abdominal vessels:Document:MRI.angio
C0881775|Multisection^W contrast IV:Find:Pt:Abdominal vessels:Doc:MRI.angio
C0881806|Deprecated Abd>Retroperitoneum CT W cont
C0881806|Multisection^W contrast:Find:Pt:Abdomen>Retroperitoneum:Doc:CT
C0881806|Multisection^W contrast:Finding:Point in time:Abdomen>Retroperitoneum:Document:Computerized Tomography
C0881806|Deprecated Abdomen>Retroperitoneum CT W contrast
C0881865|Chest XR PA Upr W insp+exp
C0881865|Chest X-ray PA upright W inspiration and expiration
C0881865|Views PA upright^W inspiration & expiration:Find:Pt:Chest:Doc:XR
C0881865|Views PA upright^W inspiration & expiration:Finding:Point in time:Chest:Document:XR
C0881873|Chest XR PA+R-Lat+R-Obl+L-Obl Upr
C0881873|Chest X-ray PA and right lateral and right oblique and left oblique upright
C0881873|Views PA & R-lateral & R-oblique & L-oblique upright:Find:Pt:Chest:Doc:XR
C0881873|Views PA & R-lateral & R-oblique & L-oblique upright:Finding:Point in time:Chest:Document:XR
C0881916|Extr US
C0881916|Extremity US
C0881916|Multisection:Find:Pt:Extremity:Doc:US
C0881916|Multisection:Finding:Point in time:Extremity:Document:Ultrasound
C0881923|Femur DXA Bone density
C0881923|Bone density:Mass Aeric:Point in time:Femur:Quantitative:XR.DXA
C0881923|Bone density:MAric:Pt:Femur:Qn:XR.DXA
C0881923|Femur DXA BDM
C0881942|Wrist+Hand XR Bone Age
C0881942|Wrist and Hand X-ray bone age
C0881942|Views bone age:Finding:Point in time:Wrist+Hand:Document:XR
C0881942|Views bone age:Find:Pt:Wrist+Hand:Doc:XR
C0882007|Knee XR AP+PA stand
C0882007|Knee X-ray AP and PA standing
C0882007|Views AP & PA^standing:Find:Pt:Knee:Doc:XR
C0882007|Views AP & PA^standing:Finding:Point in time:Knee:Document:XR
C1114477|Head.cistern MRI
C1114477|Head Cistern MRI
C1114477|Multisection:Finding:Point in time:Head.cistern:Document:MRI
C1114477|Multisection:Find:Pt:Head.cistern:Doc:MRI
C1114544|Zygomatic arch-Bl XR port
C1114544|Zygomatic arch - bilateral X-ray portable
C1114544|Views portable:Finding:Point in time:Zygomatic arch.bilateral:Document:XR
C1114544|Views portable:Find:Pt:Zygomatic arch.bilateral:Doc:XR
C1114556|Chest XR PA+Lat+R-or-L-Obl
C1114556|Chest X-ray PA and lateral and right or-left oblique
C1114556|Views PA & lateral & R-or-L-oblique:Find:Pt:Chest:Doc:XR
C1114556|Views PA & lateral & R-or-L-oblique:Finding:Point in time:Chest:Document:XR
C1114584|Ankle XR AP+Lat
C1114584|Ankle X-ray AP and lateral
C1114584|Views AP & lateral:Find:Pt:Ankle:Doc:XR
C1114584|Views AP & lateral:Finding:Point in time:Ankle:Document:XR
C1114597|Patella X-ray portable
C1114597|Patella XR port
C1114597|Views portable:Finding:Point in time:Patella:Document:XR
C1114597|Views portable:Find:Pt:Patella:Doc:XR
C1114950|Lung-Bl XR W contr IB
C1114950|Lung - bilateral X-ray W contrast intrabronchial
C1114950|Views^W contrast intrabronchial:Find:Pt:Lung.bilateral:Doc:XR
C1114950|Views^W contrast intrabronchial:Finding:Point in time:Lung.bilateral:Document:XR
C1114615|Fluoroscopy Guidance for injection of Spine Thoracic Facet Joint
C1114615|T-spine facet joint Flr Inj guid
C1114615|Guidance for injection:Find:Pt:Spine.thoracic facet joint:Doc:XR.fluor
C1114615|Guidance for injection:Finding:Point in time:Spine.thoracic facet joint:Document:XR.fluor
C1114684|Temporomandibular joint - left X-ray
C1114684|TMJ-L XR
C1114684|Views:Finding:Point in time:Temporomandibular joint.left:Document:XR
C1114684|Views:Find:Pt:Temporomandibular joint.left:Doc:XR
C1543438|Ribs upper post-L XR
C1543438|Ribs upper posterior - left X-ray
C1543438|Views:Finding:Point in time:Ribs.upper.posterior.left:Document:XR
C1543438|Views:Find:Pt:Ribs.upper.posterior.left:Doc:XR
C1543777|Hrt SPECT PF Rest+W ADE+Tl201 IV
C1543777|Heart SPECT perfusion at rest and W adenosine and W Tl-201 IV
C1543777|Multisection perfusion^at rest & W adenosine & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543777|Multisection perfusion^at rest & W adenosine & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543487|T-spine XR AP 1V W L-bending
C1543487|View AP^W L-bending:Find:Pt:Spine.thoracic:Doc:XR
C1543487|View AP^W L-bending:Finding:Point in time:Spine.thoracic:Document:XR
C1543487|Thoracic spine X-ray AP single view W left bending
C1543791|Pancreas RI W RNC IV
C1543791|Pancreas Scan
C1543791|Views^W radionuclide IV:Find:Pt:Pancreas:Doc:Radnuc
C1543791|Views^W radionuclide Intravenous:Finding:Point in time:Pancreas:Document:Radnuc
C1543870|RI for ETr WB W In-111-P IV
C1543870|Scan for endocrine tumor whole body W In-111 pentetreotide IV
C1543870|Views for endocrine tumor whole body^W In-111 pentetreotide IV:Find:Pt:^Patient:Doc:Radnuc
C1543870|Views for endocrine tumor whole body^W In-111 pentetreotide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543909|Hrt RI FP+EF Rest+W RNC IV
C1543909|Heart Scan first pass and ejection fraction at rest and W radionuclide IV
C1543909|Views first pass & ejection fraction^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543909|Views first pass & ejection fraction^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543916|Heart Scan static for shunt detection
C1543916|Hrt RI Static for Shunt Det W RNC IV
C1543916|Views static for shunt detection^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543916|Views static for shunt detection^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543183|Ribs X-ray 3 views
C1543183|Ribs XR 3V
C1543183|Views 3:Find:Pt:Ribs:Doc:XR
C1543183|Views 3:Finding:Point in time:Ribs:Document:XR
C1543262|BM MRI for Blood Flow
C1543262|Bone marrow MRI for blood flow
C1543262|Multisection for blood flow:Finding:Point in time:Bone marrow:Document:MRI
C1543262|Multisection for blood flow:Find:Pt:Bone marrow:Doc:MRI
C1543686|Adrenal RI W I-131 NP59 IV
C1543686|Adrenal gland Scan W I-131 NP59 IV
C1543686|Views^W I-131 NP59 IV:Find:Pt:Adrenal gland:Doc:Radnuc
C1543686|Views^W I-131 NP59 Intravenous:Finding:Point in time:Adrenal gland:Document:Radnuc
C1543713|Hrt RI W ADE+Tl-201 IV
C1543713|Heart Scan W adenosine and W Tl-201 IV
C1543713|Views^W adenosine & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543713|Views^W adenosine & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1542966|Rectum Scan W radionuclide PO
C1542966|Rectum RI W RNC PO
C1542966|Views^W radionuclide PO:Find:Pt:Rectum:Doc:Radnuc
C1542966|Views^W radionuclide Oral:Finding:Point in time:Rectum:Document:Radnuc
C1542967|Esophagus Scan for motility W radionuclide PO
C1542967|Esoph RI for Motility W RNC PO
C1542967|Views for motility^W radionuclide PO:Find:Pt:Esophagus:Doc:Radnuc
C1542967|Views for motility^W radionuclide Oral:Finding:Point in time:Esophagus:Document:Radnuc
C1526777|Brst Specimen-R Mam
C1526777|Breast specimen - right Mammogram
C1526777|Views:Finding:Point in time:Breast specimen.right:Document:Mam
C1526777|Views:Find:Pt:Breast specimen.right:Doc:Mam
C1526778|Should-R XR AP+Transthoracic
C1526778|Shoulder - right X-ray AP and transthoracic
C1526778|Views AP & transthoracic:Finding:Point in time:Shoulder.right:Document:XR
C1526778|Views AP & transthoracic:Find:Pt:Shoulder.right:Doc:XR
C1526803|Hand-L XR AP+Lat
C1526803|Hand - left X-ray AP and lateral
C1526803|Views AP & lateral:Finding:Point in time:Hand.left:Document:XR
C1526803|Views AP & lateral:Find:Pt:Hand.left:Doc:XR
C1526815|UE vv-L XRA W contr IV
C1526815|Upper extremity veins - left Fluoroscopic angiogram W contrast IV
C1526815|Views^W contrast IV:Find:Pt:Upper extremity veins.left:Doc:XR.fluor.angio
C1526815|Views^W contrast Intravenous:Finding:Point in time:Upper extremity veins.left:Document:XR.fluor.angio
C1524183|Sternum CT
C1524183|Multisection:Find:Pt:Sternum:Doc:CT
C1524183|Multisection:Finding:Point in time:Sternum:Document:Computerized Tomography
C1524847|Femur - left CT WO contrast
C1524847|Femur-L CT WO contr
C1524847|Multisection^WO contrast:Finding:Point in time:Femur.left:Document:Computerized Tomography
C1524847|Multisection^WO contrast:Find:Pt:Femur.left:Doc:CT
C1525098|BDs+GB CT Drain guid
C1525098|CT Guidance for drainage of Biliary ducts and Gallbladder
C1525098|Guidance for drainage:Find:Pt:Abdomen>Biliary ducts+Gallbladder:Doc:CT
C1525098|Guidance for drainage:Finding:Point in time:Abdomen>Biliary ducts+Gallbladder:Document:Computerized Tomography
C1525105|Orbit-R MRI
C1525105|Orbit - right MRI
C1525105|Multisection:Finding:Point in time:Orbit.right:Document:MRI
C1525105|Multisection:Find:Pt:Orbit.right:Doc:MRI
C1525108|Subclavian a MRI.Angio
C1525108|Subclavian artery MRI angiogram
C1525108|Multisection:Find:Pt:Subclavian artery:Doc:MRI.angio
C1525108|Multisection:Finding:Point in time:Subclavian artery:Document:MRI.angio
C1525211|Deprecated Temporal bones MRI W & WO contrast IV
C1525211|Deprecated Temporal bones MRI W+WO contr
C1525211|Multisection^W & WO contrast IV:Find:Pt:Temporal bone:Nar:MRI
C1525211|Multisection^W & WO contrast Intravenous:Finding:Point in time:Temporal bone:Narrative:MRI
C1525245|Joint MRI WO contrast
C1525245|Joint MRI WO contr
C1525245|Multisection^WO contrast:Find:Pt:Joint:Doc:MRI
C1525245|Multisection^WO contrast:Finding:Point in time:Joint:Document:MRI
C1525246|Orbit-L MRI WO contr
C1525246|Orbit - left MRI WO contrast
C1525246|Multisection^WO contrast:Find:Pt:Orbit.left:Doc:MRI
C1525246|Multisection^WO contrast:Finding:Point in time:Orbit.left:Document:MRI
C1525247|Orbit-R MRI WO contr
C1525247|Orbit - right MRI WO contrast
C1525247|Multisection^WO contrast:Finding:Point in time:Orbit.right:Document:MRI
C1525247|Multisection^WO contrast:Find:Pt:Orbit.right:Doc:MRI
C1525251|Abd ves MRI.Angio WO contr
C1525251|Abdominal vessels MRI angiogram WO contrast
C1525251|Multisection^WO contrast:Finding:Point in time:Abdominal vessels:Document:MRI.angio
C1525251|Multisection^WO contrast:Find:Pt:Abdominal vessels:Doc:MRI.angio
C1525253|Carot ves MRI.Angio WO contr
C1525253|Carotid vessel MRI angiogram WO contrast
C1525253|Multisection^WO contrast:Find:Pt:Carotid vessel:Doc:MRI.angio
C1525253|Multisection^WO contrast:Finding:Point in time:Carotid vessel:Document:MRI.angio
C1525456|Brst-Bl Mam Tangential
C1525456|Breast - bilateral Mammogram tangential
C1525456|View tangential:Find:Pt:Breast.bilateral:Doc:Mam
C1525456|View tangential:Finding:Point in time:Breast.bilateral:Document:Mam
C1525462|Shoulder - bilateral X-ray Grashey
C1525462|Should-Bl XR Grashey
C1525462|View Grashey:Find:Pt:Shoulder.bilateral:Doc:XR
C1525462|View Grashey:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525470|Wrist - left X-ray ulnar deviation
C1525470|Wrist-L XR Ulnar Deviation
C1525470|View ulnar deviation:Finding:Point in time:Wrist.left:Document:XR
C1525470|View ulnar deviation:Find:Pt:Wrist.left:Doc:XR
C1525536|Kidney XR Ltd W contr IV
C1525536|Views limited^W contrast IV:Find:Pt:Kidney:Doc:XR
C1525536|Kidney X-ray limited W contrast IV
C1525536|Views limited^W contrast Intravenous:Finding:Point in time:Kidney:Document:XR
C1525547|Mandible XR PA+Lat+Obl+Towne
C1525547|Mandible X-ray PA and lateral and oblique and Towne
C1525547|Views PA & lateral & oblique & Towne:Finding:Point in time:Mandible:Document:XR
C1525547|Views PA & lateral & oblique & Towne:Find:Pt:Mandible:Doc:XR
C1525605|Toes-L XR stand
C1525605|Toes - left X-ray standing
C1525605|Views^standing:Find:Pt:Toes.left:Doc:XR
C1525605|Views^standing:Finding:Point in time:Toes.left:Document:XR
C1525612|Deprecated Aorta.endograft CT
C1525612|Multisection:Finding:Point in time:Aorta.endograft:Document:Computerized Tomography
C1525612|Multisection:Find:Pt:Aorta.endograft:Doc:CT
C1525682|Humerus bicipital groove - left X-ray
C1525682|Humerus bicipital groove-L XR
C1525682|Views:Find:Pt:Humerus.bicipital groove.left:Doc:XR
C1525682|Views:Finding:Point in time:Humerus.bicipital groove.left:Document:XR
C1525696|L-spine+Sacrum XR 5V
C1525696|Spine Lumbar and Sacrum X-ray 5 views
C1525696|Views 5:Finding:Point in time:Spine.lumbar+Sacrum:Document:XR
C1525696|Views 5:Find:Pt:Spine.lumbar+Sacrum:Doc:XR
C1525697|L-spine+Sacrum+Coccyx XR 5V
C1525697|Spine Lumbar and Sacrum and Coccyx X-ray 5 views
C1525697|Views 5:Find:Pt:Spine.lumbar+Sacrum+Coccyx:Doc:XR
C1525697|Views 5:Finding:Point in time:Spine.lumbar+Sacrum+Coccyx:Document:XR
C1524700|Wrist - bilateral X-ray 3 views
C1524700|Wrist-Bl XR 3V
C1524700|Views 3:Find:Pt:Wrist.bilateral:Doc:XR
C1524700|Views 3:Finding:Point in time:Wrist.bilateral:Document:XR
C1525778|Hand - bilateral X-ray Bora
C1525778|Hand-Bl XR Bora
C1525778|View Bora:Find:Pt:Hand.bilateral:Doc:XR
C1525778|View Bora:Finding:Point in time:Hand.bilateral:Document:XR
C1525857|Knee-Bl XR W Stress
C1525857|Knee - bilateral X-ray W manual stress
C1525857|Views^W manual stress:Find:Pt:Knee.bilateral:Doc:XR
C1525857|Views^W manual stress:Finding:Point in time:Knee.bilateral:Document:XR
C1525873|Acromioclavicular Joint X-ray W weight
C1525873|AC joint XR W Wt
C1525873|Views^W weight:Finding:Point in time:Acromioclavicular joint:Document:XR
C1525873|Views^W weight:Find:Pt:Acromioclavicular joint:Doc:XR
C1525891|Eye US FB local guid
C1525891|US Guidance for localization of foreign body of Eye
C1525891|Guidance for localization of foreign body:Finding:Point in time:Eye:Document:Ultrasound
C1525891|Guidance for localization of foreign body:Find:Pt:Eye:Doc:US
C1525943|Pelvis XR Ferguson
C1525943|Pelvis X-ray Ferguson
C1525943|View Ferguson:Finding:Point in time:Pelvis:Document:XR
C1525943|View Ferguson:Find:Pt:Pelvis:Doc:XR
C1525839|Brst-Bl Mam Mag
C1525839|Breast - bilateral Mammogram magnification
C1525839|Views magnification:Find:Pt:Breast.bilateral:Doc:Mam
C1525839|Views magnification:Finding:Point in time:Breast.bilateral:Document:Mam
C1525963|Sacroiliac Joint X-ray limited
C1525963|SIJ XR Ltd
C1525963|Views limited:Find:Pt:Sacroiliac joint:Doc:XR
C1525963|Views limited:Finding:Point in time:Sacroiliac joint:Document:XR
C1525972|Scapula X-ray 2 views
C1525972|Scapula XR 2V
C1525972|Views 2:Finding:Point in time:Scapula:Document:XR
C1525972|Views 2:Find:Pt:Scapula:Doc:XR
C1526005|Femur-R XR 1V
C1526005|Femur - right X-ray Single view
C1526005|View 1:Find:Pt:Femur.right:Doc:XR
C1526005|View 1:Finding:Point in time:Femur.right:Document:XR
C1526115|Acromioclavicular joint - right X-ray Zanca
C1526115|AC joint-R XR Zanca
C1526115|View Zanca:Finding:Point in time:Acromioclavicular joint.right:Document:XR
C1526115|View Zanca:Find:Pt:Acromioclavicular joint.right:Doc:XR
C1525903|Wrist - right X-ray lateral W extension
C1525903|Wrist-R XR Lat W Ext
C1525903|View lateral^W extension:Finding:Point in time:Wrist.right:Document:XR
C1525903|View lateral^W extension:Find:Pt:Wrist.right:Doc:XR
C1525904|Wrist - right X-ray lateral W flexion
C1525904|Wrist-R XR Lat W Flx
C1525904|View lateral^W flexion:Finding:Point in time:Wrist.right:Document:XR
C1525904|View lateral^W flexion:Find:Pt:Wrist.right:Doc:XR
C1526033|Hand-R XRTomo
C1526033|Hand - right X-ray tomograph
C1526033|Multisection:Find:Pt:Hand.right:Doc:XR.tomo
C1526033|Multisection:Finding:Point in time:Hand.right:Document:XR.tomo
C1526097|Should-R XR 1V
C1526097|Shoulder - right X-ray Single view
C1526097|View 1:Find:Pt:Shoulder.right:Doc:XR
C1526097|View 1:Finding:Point in time:Shoulder.right:Document:XR
C1526198|US Guidance for biopsy of Neck
C1526198|Neck US Bx guid
C1526198|Guidance for biopsy:Find:Pt:Neck:Doc:US
C1526198|Guidance for biopsy:Finding:Point in time:Neck:Document:Ultrasound
C1526228|Ribs anterior - right X-ray
C1526228|Ribs Ant-R XR
C1526228|Views:Finding:Point in time:Ribs.anterior.right:Document:XR
C1526228|Views:Find:Pt:Ribs.anterior.right:Doc:XR
C1526245|Visceral vessels Fluoroscopic angiogram W contrast
C1526245|Visceral ves XRA W contr
C1526245|Views^W contrast:Find:Pt:Visceral vessels:Doc:XR.fluor.angio
C1526245|Views^W contrast:Finding:Point in time:Visceral vessels:Document:XR.fluor.angio
C1526285|UE-R US
C1526285|Upper extremity - right US
C1526285|Multisection:Finding:Point in time:Upper extremity.right:Document:Ultrasound
C1526285|Multisection:Find:Pt:Upper extremity.right:Doc:US
C1524485|Multisection^W contrast IV:Find:Pt:Chest+Abdomen>Aorta:Doc:CT.angio
C1524485|Multisection^W contrast Intravenous:Finding:Point in time:Chest+Abdomen>Aorta:Document:Computerized Tomography.angio
C1524485|Chest+Abd Aorta CT.Angio W contr IV
C1524485|Chest and Abdomen Aorta CT angiogram W contrast IV
C1524488|Aortic arch CT angiogram W contrast IV
C1524488|Multisection^W contrast IV:Find:Pt:Chest>Aortic arch:Doc:CT.angio
C1524488|Multisection^W contrast Intravenous:Finding:Point in time:Chest>Aortic arch:Document:Computerized Tomography.angio
C1524488|Ao arch CT.Angio W contr IV
C1524856|Foot - right MRI WO contrast
C1524856|Ft-R MRI WO contr
C1524856|Multisection^WO contrast:Find:Pt:Foot.right:Doc:MRI
C1524856|Multisection^WO contrast:Finding:Point in time:Foot.right:Document:MRI
C1524535|Hand CT W contr IV
C1524535|Hand CT W contrast IV
C1524535|Multisection^W contrast Intravenous:Finding:Point in time:Hand:Document:Computerized Tomography
C1524535|Multisection^W contrast IV:Find:Pt:Hand:Doc:CT
C1524907|Spine MRI WO contr
C1524907|Spine MRI WO contrast
C1524907|Multisection^WO contrast:Find:Pt:Spine:Doc:MRI
C1524907|Multisection^WO contrast:Finding:Point in time:Spine:Document:MRI
C1524908|T-spine MRI WO contr
C1524908|Multisection^WO contrast:Find:Pt:Spine.thoracic:Doc:MRI
C1524908|Multisection^WO contrast:Finding:Point in time:Spine.thoracic:Document:MRI
C1524908|Thoracic spine MRI WO contrast
C1524559|Knee-L CT W contr IV
C1524559|Knee - left CT W contrast IV
C1524559|Multisection^W contrast Intravenous:Finding:Point in time:Knee.left:Document:Computerized Tomography
C1524559|Multisection^W contrast IV:Find:Pt:Knee.left:Doc:CT
C1524218|View AP portable:Finding:Point in time:Abdomen:Narrative:XR
C1524218|Abdomen X-ray AP portable single view
C1524218|Abd XR AP V1 port
C1524218|View AP portable:Find:Pt:Abdomen:Doc:XR
C1524218|View AP portable:Finding:Point in time:Abdomen:Document:XR
C1524283|Guidance for drainage of abscess:Find:Pt:Abdomen:Doc:CT
C1524283|Abd CT Abscess drain guid
C1524283|CT Guidance for drainage of abscess of Abdomen
C1524283|Guidance for drainage of abscess:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524302|Prostate CT Bx guid
C1524302|CT Guidance for biopsy of Prostate
C1524302|Guidance for biopsy:Find:Pt:Prostate:Doc:CT
C1524302|Guidance for biopsy:Finding:Point in time:Prostate:Document:Computerized Tomography
C1524950|Hip X-ray lateral
C1524950|Hip XR Lat
C1524950|View lateral:Find:Pt:Hip:Doc:XR
C1524950|View lateral:Finding:Point in time:Hip:Document:XR
C1524315|CT Guidance for drainage of Chest
C1524315|Chest CT Drain guid
C1524315|Guidance for drainage:Find:Pt:Chest:Doc:CT
C1524315|Guidance for drainage:Finding:Point in time:Chest:Document:Computerized Tomography
C1524316|CT Guidance for drainage of Gallbladder
C1524316|Abd GB CT Drain guid
C1524316|Guidance for drainage:Find:Pt:Abdomen>Gallbladder:Doc:CT
C1524316|Guidance for drainage:Finding:Point in time:Abdomen>Gallbladder:Document:Computerized Tomography
C1524343|Aorta MRI.Angio
C1524343|Aorta MRI angiogram
C1524343|Multisection:Find:Pt:Aorta:Doc:MRI.angio
C1524343|Multisection:Finding:Point in time:Aorta:Document:MRI.angio
C1524346|Aortic arch MRI angiogram
C1524346|Ac arch MRI.Angio
C1524346|Multisection:Find:Pt:Aortic arch:Doc:MRI.angio
C1524346|Multisection:Finding:Point in time:Aortic arch:Document:MRI.angio
C1524626|Elbow-Bl XR 3V
C1524626|Elbow - bilateral X-ray 3 views
C1524626|Views 3:Find:Pt:Elbow.bilateral:Doc:XR
C1524626|Views 3:Finding:Point in time:Elbow.bilateral:Document:XR
C1524661|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.left:Document:Computerized Tomography
C1524661|Upper extremity - left CT WO and W contrast IV
C1524661|UE-L CT WO+W contr IV
C1524661|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.left:Doc:CT
C1524992|Chest Fluoroscopy 2 views
C1524992|Chest Flr 2V
C1524992|Views 2:Finding:Point in time:Chest:Document:XR.fluor
C1524992|Views 2:Find:Pt:Chest:Doc:XR.fluor
C1525004|Acromioclavicular joint - left X-ray 2 views
C1525004|AC joint-L XR 2V
C1525004|Views 2:Find:Pt:Acromioclavicular joint.left:Doc:XR
C1525004|Views 2:Finding:Point in time:Acromioclavicular joint.left:Document:XR
C1524733|Forearm CT WO and W contrast IV
C1524733|Forearm CT WO+W contr IV
C1524733|Multisection^WO & W contrast Intravenous:Finding:Point in time:Forearm:Document:Computerized Tomography
C1524733|Multisection^WO & W contrast IV:Find:Pt:Forearm:Doc:CT
C1524766|Knee - left CT WO and W contrast IV
C1524766|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee.left:Document:Computerized Tomography
C1524766|Knee-L CT WO+W contr IV
C1524766|Multisection^WO & W contrast IV:Find:Pt:Knee.left:Doc:CT
C1525048|Knee XR AP+Lat
C1525048|Knee X-ray AP and lateral
C1525048|Views AP & lateral:Find:Pt:Knee:Doc:XR
C1525048|Views AP & lateral:Finding:Point in time:Knee:Document:XR
C1525049|Knee-L XR AP+Lat
C1525049|Knee - left X-ray AP and lateral
C1525049|Views AP & lateral:Finding:Point in time:Knee.left:Document:XR
C1525049|Views AP & lateral:Find:Pt:Knee.left:Doc:XR
C1524776|Sacrum MRI WO+W contr IV
C1524776|Sacrum MRI WO and W contrast IV
C1524776|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sacrum:Document:MRI
C1524776|Multisection^WO & W contrast IV:Find:Pt:Sacrum:Doc:MRI
C1524794|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower leg.left:Document:Computerized Tomography
C1524794|Multisection^WO & W contrast IV:Find:Pt:Lower leg.left:Doc:CT
C1524794|Lower leg - left CT WO and W contrast IV
C1524794|Lower leg-L CT WO+W contr IV
C1525082|Mandible XR PA+Lat
C1525082|Mandible X-ray PA and lateral
C1525082|Views PA & lateral:Find:Pt:Mandible:Doc:XR
C1525082|Views PA & lateral:Finding:Point in time:Mandible:Document:XR
C1830198|Multisection^W radionuclide Intravenous:Finding:Point in time:^Patient:Narrative:Radnuc.SPECT
C1830198|SPECT W RNC IV
C1830198|SPECT
C1830198|Multisection^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1830198|Multisection^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1830256|Breast - left FFD mammogram screening
C1830256|Views screening:Find:Pt:Breast.left:Doc:Mam.FFD
C1830256|Views screening:Finding:Point in time:Breast.left:Document:Mam.FFD
C1830256|Brst-L FFDM Screening
C1830261|Ac arch MRI.Angio WO+W contr IV
C1830261|Multisection^WO & W contrast Intravenous:Finding:Point in time:Aortic arch:Document:MRI.angio
C1830261|Multisection^WO & W contrast IV:Find:Pt:Aortic arch:Doc:MRI.angio
C1830261|Aortic arch MRI angiogram WO and W contrast IV
C1831071|Knee-L XR 1V or 2V
C1831071|Knee - left X-ray 1 or 2 views
C1831071|Views 1 or 2:Finding:Point in time:Knee.left:Document:XR
C1831071|Views 1 or 2:Find:Pt:Knee.left:Doc:XR
C1830075|Mastoid X-ray GE 3 views
C1830075|Mastoid XR GE 3V
C1830075|Views GE 3:Find:Pt:Mastoid:Doc:XR
C1830075|Views GE 3:Finding:Point in time:Mastoid:Document:XR
C1715382|CT Guidance for needle localization of Breast
C1715382|Brst CT Needle local guid
C1715382|Guidance for needle localization:Find:Pt:Breast:Doc:CT
C1715382|Guidance for needle localization:Finding:Point in time:Breast:Document:Computerized Tomography
C1715402|Aorta MRI angiogram WO contrast
C1715402|Aorta MRI.Angio WO contr
C1715402|Multisection^WO contrast:Find:Pt:Aorta:Doc:MRI.angio
C1715402|Multisection^WO contrast:Finding:Point in time:Aorta:Document:MRI.angio
C1715469|Orbit XR for FB
C1715469|Orbit X-ray for foreign body
C1715469|Views for foreign body:Find:Pt:Orbit:Doc:XR
C1715469|Views for foreign body:Finding:Point in time:Orbit:Document:XR
C1715481|Fluoroscopy Guidance for deep aspiration.fine needle of Tissue
C1715481|Guidance for deep aspiration.fine needle:Finding:Point in time:Tissue:Document:XR.fluor
C1715481|tiss Flr Guide for deep FNA
C1715481|Guidance for deep aspiration.fine needle:Find:Pt:Tissue:Doc:XR.fluor
C1639406|Fluoroscopy Guidance for biopsy of Prostate
C1639406|Prostate Flr Bx guid
C1639406|Guidance for biopsy:Find:Pt:Prostate:Doc:XR.fluor
C1639406|Guidance for biopsy:Finding:Point in time:Prostate:Document:XR.fluor
C1635071|Pulm CT W 133Xe IH
C1635071|Multisection^W Xe-133 IH:Find:Pt:Pulmonary system:Doc:CT
C1635071|Pulmonary system CT W Xe-133 IH
C1635071|Multisection^W Xe-133 Inhalation:Finding:Point in time:Pulmonary system:Document:Computerized Tomography
C1714904|Deprecated Aorta and Lower extremity vessels CT angiogram W contrast IV
C1714904|Multisection^W contrast Intravenous:Finding:Point in time:Aorta+Lower extremity vessels:Document:Computerized Tomography.angio
C1714904|Deprecated Aorta+LE ves CT.Angio W contr
C1714904|Multisection^W contrast IV:Find:Pt:Aorta+Lower extremity vessels:Doc:CT.angio
C1714910|Multisection^WO & W contrast IV:Find:Pt:Axilla.left:Doc:MRI
C1714910|Axilla - left MRI WO and W contrast IV
C1714910|Multisection^WO & W contrast Intravenous:Finding:Point in time:Axilla.left:Document:MRI
C1714910|Axilla-L MRI WO+W contr IV
C1714934|L-spine XRVideo
C1714934|Views:Finding:Point in time:Spine.lumbar:Document:XR.fluor.video
C1714934|Views:Find:Pt:Spine.lumbar:Doc:XR.fluor.video
C1714934|Lumbar spine Fluoroscopy video
C1714936|C-spine XR 2V or 3V
C1714936|Views 2 or 3:Find:Pt:Spine.cervical:Doc:XR
C1714936|Views 2 or 3:Finding:Point in time:Spine.cervical:Document:XR
C1714936|Cervical spine X-ray 2 or 3 views
C1714943|ves-L XRA W contr IV
C1714943|Views^W contrast Intravenous:Finding:Point in time:Vessels.left:Document:XR.fluor.angio
C1714943|Views^W contrast IV:Find:Pt:Vessels.left:Doc:XR.fluor.angio
C1714943|Vessels - left Fluoroscopic angiogram W contrast IV
C1714952|US Guidance for biopsy of Superficial muscle
C1714952|Superf Muscle US Bx guid
C1714952|Guidance for biopsy:Find:Pt:Superficial muscle:Doc:US
C1714952|Guidance for biopsy:Finding:Point in time:Superficial muscle:Document:Ultrasound
C1717268|Heart Scan for infarct quantitative
C1717268|Hrt RI for Infarct Qn W RNC IV
C1717268|Views for infarct quantitative^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1717268|Views for infarct quantitative^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1643611|Chest X-ray 2 views and apical
C1643611|Chest XR 2V+Apical
C1643611|Views 2 & apical:Finding:Point in time:Chest:Document:XR
C1643611|Views 2 & apical:Find:Pt:Chest:Doc:XR
C1634500|C-spine CT Needle local guid
C1634500|Guidance for needle localization:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C1634500|Guidance for needle localization:Find:Pt:Spine.cervical:Doc:CT
C1634500|CT Guidance for needle localization of Cervical spine
C1627296|Guidance for drainage of abscess:Finding:Point in time:Liver:Document:Ultrasound
C1627296|Liver US Abscess drain guid
C1627296|US Guidance for drainage of abscess of Liver
C1627296|Guidance for drainage of abscess:Find:Pt:Liver:Doc:US
C1638886|US Guidance for percutaneous biopsy of Muscle
C1638886|Muscle US PC Bx guid
C1638886|Guidance for percutaneous biopsy:Find:Pt:Muscle:Doc:US
C1638886|Guidance for percutaneous biopsy:Finding:Point in time:Muscle:Document:Ultrasound
C1648937|Views^W Tc-99m DMSA IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1648937|Kidney - bilateral Scan W Tc-99m DMSA IV
C1648937|Views^W Tc-99m DMSA Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1648937|Kdny-Bl RI W Tc99mDMCA IV
C1633402|Views & AP KUB^W air contrast PO:Find:Pt:Gastrointestine.upper:Nar:XR.fluor
C1633402|Deprecated UGI Flr +AP W contr PO
C1633402|Deprecated Gastrointestine upper Fluoroscopy & AP W contrast PO
C1633402|Views & AP KUB^W air contrast Oral:Finding:Point in time:Gastrointestine.upper:Narrative:XR.fluor
C1631260|Pancreas CT Drain guid
C1631260|CT Guidance for drainage of Pancreas
C1631260|Guidance for drainage:Find:Pt:Abdomen>Pancreas:Doc:CT
C1631260|Guidance for drainage:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C1978444|Wrist+Hand-L XR
C1978444|Wrist - left and Hand - left X-ray
C1978444|Views:Finding:Point in time:Wrist.left+Hand.left:Document:XR
C1978444|Views:Find:Pt:Wrist.left+Hand.left:Doc:XR
C1954154|Gastric emptying time^post 100 mg sodium acetate PO:Time:Pt:Exhl gas:Qn:Radnuc
C1954154|Exhaled gas Scan Gastric emptying time post 100 mg sodium acetate PO
C1954154|ExG RI GE time p 100mg Na acetate PO
C1954154|Gastric emptying time^post 100 mg sodium acetate Oral:Time:Point in time:Exhaled gas (breath):Quantitative:Radnuc
C1954310|Submandibular gland - right Fluoroscopy W contrast intra salivary duct
C1954310|Submandib gland-R Flr W contr intra SD
C1954310|Views^W contrast intra salivary duct:Find:Pt:Submandibular gland.right:Doc:XR.fluor
C1954310|Views^W contrast intra salivary duct:Finding:Point in time:Submandibular gland.right:Document:XR.fluor
C1953973|SIJ XR 1V or 2V
C1953973|Sacroiliac Joint X-ray 1 or 2 views
C1953973|Views 1 or 2:Find:Pt:Sacroiliac joint:Doc:XR
C1953973|Views 1 or 2:Finding:Point in time:Sacroiliac joint:Document:XR
C1953974|Ribs - bilateral and Chest X-ray 2 views and PA chest
C1953974|Views 2 & PA chest:Finding:Point in time:Ribs.bilateral+Chest:Document:XR
C1953974|Views 2 & PA chest:Find:Pt:Ribs.bilateral+Chest:Doc:XR
C1953974|Ribs-Bl+Chest XR 2V+PA Chst
C3533555|Fluoroscopy Guidance for removal of CVA device obstruction from Central vein
C3533555|Centl v Flr CVA dev obs rem guid
C3533555|Guidance for removal of CVA device obstruction:Find:Pt:Central vein:Doc:XR.fluor
C3533555|Guidance for removal of CVA device obstruction:Finding:Point in time:Central vein:Document:XR.fluor
C3533802|Multisection^W contrast Intravenous:Finding:Point in time:Toes.left:Document:MRI
C3533802|Toes-L MRI W contr IV
C3533802|Multisection^W contrast IV:Find:Pt:Toes.left:Doc:MRI
C3533802|Toes - left MRI W contrast IV
C3262947|Guidance for superficial aspiration.fine needle:Find:Pt:Tiss:Doc:XR.fluor
C3262947|Tiss Flr Sup FNA guid
C3262947|Guidance for superficial aspiration.fine needle:Finding:Point in time:Tissue, unspecified:Document:XR.fluor
C3262947|Fluoroscopy Guidance for superficial aspiration.fine needle of Tissue
C3262983|Ankle-Bl MRI W contr IV
C3262983|Ankle - bilateral MRI W contrast IV
C3262983|Multisection^W contrast Intravenous:Finding:Point in time:Ankle.bilateral:Document:MRI
C3262983|Multisection^W contrast IV:Find:Pt:Ankle.bilateral:Doc:MRI
C3262992|Femur - bilateral MRI W contrast IV
C3262992|Femur-Bl MRI W contr IV
C3262992|Multisection^W contrast IV:Find:Pt:Femur.bilateral:Doc:MRI
C3262992|Multisection^W contrast Intravenous:Finding:Point in time:Femur.bilateral:Document:MRI
C3262996|Forearm - bilateral MRI WO contrast
C3262996|Forearm-Bl MRI WO contr
C3262996|Multisection^WO contrast:Find:Pt:Forearm.bilateral:Doc:MRI
C3262996|Multisection^WO contrast:Finding:Point in time:Forearm.bilateral:Document:MRI
C3263040|Deprecated Fluoroscopy Guidance for needle biopsy of Pleura
C3263040|Deprecated
C3263040|Guidance for biopsy.needle:Find:Pt:Pleura:Doc:XR.fluor
C3263040|Guidance for biopsy.needle:Finding:Point in time:Pleura:Document:XR.fluor
C3203436|Ft-L XR 1V
C3203436|Foot - left X-ray Single view
C3203436|View 1:Finding:Point in time:Foot.left:Document:XR
C3203436|View 1:Find:Pt:Foot.left:Doc:XR
C3263202|Lower extremity veins - bilateral US
C3263202|LE vv-Bl US
C3263202|Multisection:Find:Pt:Lower extremity veins.bilateral:Doc:US
C3263202|Multisection:Finding:Point in time:Lower extremity veins.bilateral:Document:Ultrasound
C3262926|Multisection^W contrast Intrasynovial:Finding:Point in time:Elbow.left:Document:Computerized Tomography
C3262926|Multisection^W contrast IS:Find:Pt:Elbow.left:Doc:CT
C3262926|Elbow - left CT W contrast IS
C3262926|Elbow-L CT W contr IS
C0942157|Radius+Ulna-Bl XR
C0942157|Radius - bilateral and Ulna - bilateral X-ray
C0942157|Views:Finding:Point in time:Radius.bilateral+Ulna.bilateral:Document:XR
C0942157|Views:Find:Pt:Radius.bilateral+Ulna.bilateral:Doc:XR
C0942173|Tib+Fib-Bl XR
C0942173|Tibia - bilateral and Fibula - bilateral X-ray
C0942173|Views:Find:Pt:Tibia.bilateral+Fibula.bilateral:Doc:XR
C0942173|Views:Finding:Point in time:Tibia.bilateral+Fibula.bilateral:Document:XR
C0942309|Spine facet joint-Bl Flr Inj guid
C0942309|Fluoroscopy Guidance for injection of Spine facet joint - bilateral
C0942309|Guidance for injection:Find:Pt:Spine facet joint.bilateral:Doc:XR.fluor
C0942309|Guidance for injection:Finding:Point in time:Spine facet joint.bilateral:Document:XR.fluor
C0942315|US Guidance for drainage of Kidney - bilateral
C0942315|Guidance for drainage:Find:Pt:Kidney.bilateral:Doc:US
C0942315|Guidance for drainage:Finding:Point in time:Kidney.bilateral:Document:Ultrasound
C0942315|Kdny-Bl US Drain guid
C0942326|US Guidance for biopsy of Kidney - left
C0942326|Kidney-L US Bx guid
C0942326|Guidance for biopsy:Finding:Point in time:Kidney.left:Document:Ultrasound
C0942326|Guidance for biopsy:Find:Pt:Kidney.left:Doc:US
C0942330|Breast - bilateral Mammogram diagnostic
C0942330|Brst-Bl Mam Dx
C0942330|Views diagnostic:Find:Pt:Breast.bilateral:Doc:Mam
C0942330|Views diagnostic:Finding:Point in time:Breast.bilateral:Document:Mam
C0945341|Brst-Bl Mam Dx Ltd
C0945341|Breast - bilateral Mammogram diagnostic limited
C0945341|Views diagnostic limited:Find:Pt:Breast.bilateral:Doc:Mam
C0945341|Views diagnostic limited:Finding:Point in time:Breast.bilateral:Document:Mam
C0942373|Knee - right X-ray 2 views
C0942373|Knee-R XR 2V
C0942373|Views 2:Find:Pt:Knee.right:Doc:XR
C0942373|Views 2:Finding:Point in time:Knee.right:Document:XR
C0882048|Oropharynx Fluoroscopy video
C0882048|Oropharynx XRVideo
C0882048|Views:Finding:Point in time:Oropharynx:Document:XR.fluor.video
C0882048|Views:Find:Pt:Oropharynx:Doc:XR.fluor.video
C0882058|Pelvis MRI
C0882058|Multisection:Finding:Point in time:Pelvis:Narrative:MRI
C0882058|Multisection:Finding:Point in time:Pelvis:Document:MRI
C0882058|Multisection:Find:Pt:Pelvis:Doc:MRI
C0882076|Pylorus US for pyloric stenosis
C0882076|Multisection for pyloric stenosis:Find:Pt:Pylorus:Doc:US
C0882076|Multisection for pyloric stenosis:Finding:Point in time:Pylorus:Document:Ultrasound
C0882082|Views:Finding:Point in time:Ribs:Narrative:XR
C0882082|Ribs XR
C0882082|Ribs X-ray
C0882082|Views:Find:Pt:Ribs:Doc:XR
C0882082|Views:Finding:Point in time:Ribs:Document:XR
C0882103|Skull XR Lat
C0882103|Skull X-ray lateral
C0882103|View lateral:Finding:Point in time:Skull:Document:XR
C0882103|View lateral:Find:Pt:Skull:Doc:XR
C0882555|C-spine Flr W contr IT
C0882555|Views^W contrast IT:Find:Pt:Spine.cervical:Doc:XR.fluor
C0882555|Views^W contrast Intrathecal:Finding:Point in time:Spine.cervical:Document:XR.fluor
C0882555|Cervical spine Fluoroscopy W contrast IT
C0882556|L-spine CT W contr IT
C0882556|Multisection^W contrast Intrathecal:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C0882556|Multisection^W contrast IT:Find:Pt:Spine.lumbar:Doc:CT
C0882556|Lumbar spine CT W contrast IT
C0882167|Thyroid RI +Uptake W I-131 IV
C0882167|Thyroid Scan and uptake W I-131 IV
C0882167|Views & uptake^W I-131 IV:Find:Pt:Thyroid:Doc:Radnuc
C0882167|Views & uptake^W I-131 Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C0882203|Unspecified body region CT W conscious sedation
C0882203|XXX CT W conscious sedation
C0882203|Multisection^W conscious sedation:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882203|Multisection^W conscious sedation:Find:Pt:XXX:Doc:CT
C0882211|XXX US Bx guid
C0882211|US Guidance for biopsy of Unspecified body region
C0882211|Guidance for biopsy:Find:Pt:XXX:Doc:US
C0882211|Guidance for biopsy:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C0882214|Unspecified body region X-ray Comparison view
C0882214|XXX XR Comparison
C0882214|Comparison view.XXX:Find:Pt:XXX:Doc:XR
C0882214|Comparison view.XXX:Finding:Point in time:To be specified in another part of the message:Document:XR
C0942121|Deprecated Calcaneus - left X-ray
C0942121|Views:Find:Pt:Calcaneus.left:Doc:XR
C0942121|Views:Finding:Point in time:Calcaneus.left:Document:XR
C0942121|Deprecated Heel-L XR
C0881780|Multisection^WO & W contrast IV:Find:Pt:Ankle:Doc:MRI
C0881780|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ankle:Document:MRI
C0881780|Ankle MRI WO and W contrast IV
C0881780|Ankle MRI WO+W contr IV
C0881811|BDs+GB XR W contr IV
C0881811|Biliary ducts and Gallbladder X-ray W contrast IV
C0881811|Views^W contrast IV:Find:Pt:Biliary ducts+Gallbladder:Doc:XR
C0881811|Views^W contrast Intravenous:Finding:Point in time:Biliary ducts+Gallbladder:Document:XR
C0881888|Head.cistern RI W RNC IT
C0881888|Head Cistern Scan W radionuclide IT
C0881888|Views^W radionuclide IT:Find:Pt:Head.cistern:Doc:Radnuc
C0881888|Views^W radionuclide Intrathecal:Finding:Point in time:Head.cistern:Document:Radnuc
C0881900|Multisection^WO & W contrast IV:Find:Pt:Elbow:Doc:MRI
C0881900|Elbow MRI WO+W contr IV
C0881900|Elbow MRI WO and W contrast IV
C0881900|Multisection^WO & W contrast Intravenous:Finding:Point in time:Elbow:Document:MRI
C0881935|GI Flr Decompr tube plac guid
C0881935|Fluoroscopy Guidance for placement of decompression tube in Gastrointestine
C0881935|Guidance for placement of decompression tube:Finding:Point in time:Gastrointestine:Document:XR.fluor
C0881935|Guidance for placement of decompression tube:Find:Pt:Gastrointestine:Doc:XR.fluor
C0881969|Iliac artery Fluoroscopic angiogram Angioplasty W contrast IA
C0881969|Iliac a XRA Angpsty W contr IA
C0881969|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Iliac artery:Document:XR.fluor.angio
C0881969|Angioplasty^W contrast IA:Find:Pt:Iliac artery:Doc:XR.fluor.angio
C0882009|Liver CT Asp guid
C0882009|CT Guidance for aspiration of Liver
C0882009|Guidance for aspiration:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C0882009|Guidance for aspiration:Find:Pt:Abdomen>Liver:Doc:CT
C1114510|Knee MRI WO contr
C1114510|Knee MRI WO contrast
C1114510|Multisection^WO contrast:Find:Pt:Knee:Doc:MRI
C1114510|Multisection^WO contrast:Finding:Point in time:Knee:Document:MRI
C1114518|US Guidance for injection of Thyroid
C1114518|Thyroid US Inj guid
C1114518|Guidance for injection:Finding:Point in time:Thyroid:Document:Ultrasound
C1114518|Guidance for injection:Find:Pt:Thyroid:Doc:US
C1114530|T+L-spine XR Scoli Lat
C1114530|Views scoliosis lateral:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1114530|Spine Thoracic and Lumbar X-ray scoliosis lateral
C1114530|Views scoliosis lateral:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1114567|T-spine XR Lat Port
C1114567|View lateral portable:Finding:Point in time:Spine.thoracic:Document:XR
C1114567|View lateral portable:Find:Pt:Spine.thoracic:Doc:XR
C1114567|Thoracic spine X-ray lateral portable
C1114631|Adrenal artery Fluoroscopic angiogram W contrast IA
C1114631|Adrenal a XRA W contr IA
C1114631|Views^W contrast Intra-arterial:Finding:Point in time:Adrenal artery:Document:XR.fluor.angio
C1114631|Views^W contrast IA:Find:Pt:Adrenal artery:Doc:XR.fluor.angio
C1114641|Views^W contrast transhepatic & W hemodynamics:Finding:Point in time:Portal vein:Narrative:XR.fluor.angio
C1114641|Portal v XRA W contr TH+hemodyn
C1114641|Portal vein Fluoroscopic angiogram W contrast transhepatic and W hemodynamics
C1114641|Views^W contrast transhepatic & W hemodynamics:Finding:Point in time:Portal vein:Document:XR.fluor.angio
C1114641|Views^W contrast transhepatic & W hemodynamics:Find:Pt:Portal vein:Doc:XR.fluor.angio
C1114652|Brst.duct US W contr intra Dct
C1114652|Breast duct US W contrast intra duct
C1114652|Multisection^W contrast intra duct:Find:Pt:Breast.duct:Doc:US
C1114652|Multisection^W contrast intra duct:Finding:Point in time:Breast.duct:Document:Ultrasound
C1114656|Nerves cranial MRI
C1114656|Nerves.cranial MRI
C1114656|Multisection:Find:Pt:Nerves.cranial:Doc:MRI
C1114656|Multisection:Finding:Point in time:Nerves.cranial:Document:MRI
C1114431|CT Guidance for fine needle aspiration of Liver
C1114431|Liver CT FNA Asp
C1114431|Guidance for aspiration.fine needle:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1114431|Guidance for aspiration.fine needle:Find:Pt:Abdomen>Liver:Doc:CT
C1114438|CT Guidance for fine needle aspiration of Spleen
C1114438|Spleen CT FNA Asp
C1114438|Guidance for aspiration.fine needle:Find:Pt:Abdomen>Spleen:Doc:CT
C1114438|Guidance for aspiration.fine needle:Finding:Point in time:Abdomen>Spleen:Document:Computerized Tomography
C1114439|Liver CT WO contrast
C1114439|Liver CT WO contr
C1114439|Multisection^WO contrast:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1114439|Multisection^WO contrast:Find:Pt:Abdomen>Liver:Doc:CT
C1543435|Should-Bl XR Grashey+Outlet+Serendipity
C1543435|Shoulder - bilateral X-ray Grashey and outlet and Serendipity
C1543435|Views Grashey & outlet & Serendipity:Find:Pt:Shoulder.bilateral:Doc:XR
C1543435|Views Grashey & outlet & Serendipity:Finding:Point in time:Shoulder.bilateral:Document:XR
C1543456|Ankle-R XR +Mortise
C1543456|Ankle - right X-ray and Mortise
C1543456|Views & Mortise:Find:Pt:Ankle.right:Doc:XR
C1543456|Views & Mortise:Finding:Point in time:Ankle.right:Document:XR
C1543743|Liver SPECT W Tc99mRBC IV
C1543743|Liver SPECT W Tc-99m tagged RBC IV
C1543743|Multisection^W Tc-99m tagged RBC IV:Find:Pt:Liver:Doc:Radnuc.SPECT
C1543743|Multisection^W Tc-99m tagged RBC Intravenous:Finding:Point in time:Liver:Document:Radnuc.SPECT
C1543745|Views^W radionuclide Intravenous:Finding:Point in time:Liver:Narrative:Radnuc
C1543745|Liver RI W RNC IV
C1543745|Liver Scan
C1543745|Views^W radionuclide IV:Find:Pt:Liver:Doc:Radnuc
C1543745|Views^W radionuclide Intravenous:Finding:Point in time:Liver:Document:Radnuc
C1543462|Knee - right X-ray 2 views and tunnel standing
C1543462|Knee-R XR 2V+Tunnel stand
C1543462|Views 2 & tunnel^standing:Find:Pt:Knee.right:Doc:XR
C1543462|Views 2 & tunnel^standing:Finding:Point in time:Knee.right:Document:XR
C1543468|Knee-R XR AP+Lat+R-Obl+L-Obl
C1543468|Knee - right X-ray AP and lateral and right oblique and left oblique
C1543468|Views AP & lateral & R-oblique & L-oblique:Find:Pt:Knee.right:Doc:XR
C1543468|Views AP & lateral & R-oblique & L-oblique:Finding:Point in time:Knee.right:Document:XR
C1543482|Sternum XR Lat+R-Obl+L-Obl
C1543482|Sternum X-ray lateral and right oblique and left oblique
C1543482|Views lateral & R-oblique & L-oblique:Find:Pt:Sternum:Doc:XR
C1543482|Views lateral & R-oblique & L-oblique:Finding:Point in time:Sternum:Document:XR
C1543793|Parathyroid Scan delayed
C1543793|Parathyroid RI Delayed W RNC IV
C1543793|Views delayed^W radionuclide IV:Find:Pt:Parathyroid:Doc:Radnuc
C1543793|Views delayed^W radionuclide Intravenous:Finding:Point in time:Parathyroid:Document:Radnuc
C1543794|Views^W radionuclide Intravenous:Finding:Point in time:Parathyroid:Narrative:Radnuc
C1543794|Parathyroid Scan
C1543794|Parathyroid RI W RNC IV
C1543794|Views^W radionuclide IV:Find:Pt:Parathyroid:Doc:Radnuc
C1543794|Views^W radionuclide Intravenous:Finding:Point in time:Parathyroid:Document:Radnuc
C1543875|Views perfusion^W radionuclide gaseous IH:Find:Pt:Lung:Doc:Radnuc
C1543875|Lung RI PF W RNC Gas IH
C1543875|Lung Scan perfusion W radionuclide gaseous IH
C1543875|Views perfusion^W radionuclide gaseous Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1542899|Lung RI V W RNC IH
C1542899|Views ventilation^W radionuclide Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1542899|Lung Scan ventilation W radionuclide IH
C1542899|Views ventilation^W radionuclide IH:Find:Pt:Lung:Doc:Radnuc
C1543937|Hrt RI Gated W RNC IV
C1543937|Heart Scan gated
C1543937|Views gated^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543937|Views gated^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543581|LE a-R DOP
C1543581|Lower extremity artery - right US.doppler
C1543581|Multisection:Finding:Point in time:Lower extremity artery.right:Document:Ultrasound.doppler
C1543581|Multisection:Find:Pt:Lower extremity artery.right:Doc:US.doppler
C1543178|PA XRA W contr IA
C1543178|Pulmonary artery Fluoroscopic angiogram W contrast IA
C1543178|Views^W contrast IA:Find:Pt:Pulmonary artery:Doc:XR.fluor.angio
C1543178|Views^W contrast Intra-arterial:Finding:Point in time:Pulmonary artery:Document:XR.fluor.angio
C1543199|Finger XR PA+Lat+Obl
C1543199|Finger X-ray PA and lateral and oblique
C1543199|Views PA & lateral & oblique:Finding:Point in time:Finger:Document:XR
C1543199|Views PA & lateral & oblique:Find:Pt:Finger:Doc:XR
C1543263|Head CT perfusion W contrast IV
C1543263|Multisection^W contrast IV:Find:Pt:Head:Doc:CT.perfusion
C1543263|Head CT.perfusion W contr IV
C1543263|Multisection^W contrast Intravenous:Finding:Point in time:Head:Document:Computerized Tomography.perfusion
C1543685|RI Abscess local guid WB W RNC IV
C1543685|Scan Guidance for abscess localization whole body
C1543685|Guidance for abscess localization whole body^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543685|Guidance for abscess localization whole body^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C1543699|Brain SPECT flow
C1543699|Brain SPECT Flow W RNC IV
C1543699|Multisection flow^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1543699|Multisection flow^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1543701|Brain SPECT W Tl-201 IV
C1543701|Multisection^W Tl-201 IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1543701|Multisection^W Tl-201 Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1526798|Wrist-L XR V1 tunnel.carpal
C1526798|Wrist - left X-ray tunnel.carpal
C1526798|View tunnel.carpal:Find:Pt:Wrist.left:Doc:XR
C1526798|View tunnel.carpal:Finding:Point in time:Wrist.left:Document:XR
C1543411|Should-L XR AP(w IR)+Grashey+Ax+Outlet
C1543411|Shoulder - left X-ray AP (W internal rotation) and Grashey and axillary and outlet
C1543411|Views AP (W internal rotation) & Grashey & axillary & outlet:Find:Pt:Shoulder.left:Doc:XR
C1543411|Views AP (W internal rotation) & Grashey & axillary & outlet:Finding:Point in time:Shoulder.left:Document:XR
C1524434|Maxi+Mand CT
C1524434|Maxilla and Mandible CT
C1524434|Multisection:Find:Pt:Maxilla+Mandible:Doc:CT
C1524434|Multisection:Finding:Point in time:Maxilla+Mandible:Document:Computerized Tomography
C1524846|Thigh MRI WO contrast
C1524846|Thigh MRI WO contr
C1524846|Multisection^WO contrast:Find:Pt:Thigh:Doc:MRI
C1524846|Multisection^WO contrast:Finding:Point in time:Thigh:Document:MRI
C1525212|Multisection^WO & W contrast IV:Find:Pt:Temporal bone:Doc:CT
C1525212|Temporal bone CT WO+W contr IV
C1525212|Multisection^WO & W contrast Intravenous:Finding:Point in time:Temporal bone:Document:Computerized Tomography
C1525212|Temporal bone CT WO and W contrast IV
C1525233|LE ves-R MRI.Angio WO+W contr IV
C1525233|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity vessels.right:Document:MRI.angio
C1525233|Lower extremity vessels - right MRI angiogram WO and W contrast IV
C1525233|Multisection^WO & W contrast IV:Find:Pt:Lower extremity vessels.right:Doc:MRI.angio
C1525243|UE joint-L MRI WO contr
C1525243|Upper extremity joint - left MRI WO contrast
C1525243|Multisection^WO contrast:Finding:Point in time:Upper extremity.joint.left:Document:MRI
C1525243|Multisection^WO contrast:Find:Pt:Upper extremity.joint.left:Doc:MRI
C1525255|LE ves-L MRI.Angio WO contr
C1525255|Lower extremity vessels - left MRI angiogram WO contrast
C1525255|Multisection^WO contrast:Find:Pt:Lower extremity vessels.left:Doc:MRI.angio
C1525255|Multisection^WO contrast:Finding:Point in time:Lower extremity vessels.left:Document:MRI.angio
C1526993|Adrenal CT
C1526993|Adrenal gland CT
C1526993|Multisection:Finding:Point in time:Adrenal gland:Narrative:Computerized Tomography
C1526993|Multisection:Find:Pt:Abdomen>Adrenal gland:Doc:CT
C1526993|Multisection:Finding:Point in time:Abdomen>Adrenal gland:Document:Computerized Tomography
C1524227|Brst-Bl Mam XCCL
C1524227|Breast - bilateral Mammogram XCCL
C1524227|View XCCL:Finding:Point in time:Breast.bilateral:Document:Mam
C1524227|View XCCL:Find:Pt:Breast.bilateral:Doc:Mam
C1524254|Knee XR AP+Lat+Sunrise
C1524254|Knee X-ray AP and lateral and Sunrise
C1524254|Views AP & lateral & Sunrise:Finding:Point in time:Knee:Document:XR
C1524254|Views AP & lateral & Sunrise:Find:Pt:Knee:Doc:XR
C1525524|Scapula-L XR AP+Y
C1525524|Scapula - left X-ray AP and Y
C1525524|Views AP & Y:Finding:Point in time:Scapula.left:Document:XR
C1525524|Views AP & Y:Find:Pt:Scapula.left:Doc:XR
C1114538|Views portable:Finding:Point in time:Spine.cervical:Narrative:XR
C1114538|C-spine XR port
C1114538|Views portable:Finding:Point in time:Spine.cervical:Document:XR
C1114538|Views portable:Find:Pt:Spine.cervical:Doc:XR
C1114538|Cervical spine X-ray portable
C1525580|Views^W contrast Intrasynovial:Finding:Point in time:Ankle:Document:XR.fluor
C1525580|Ankle Flr W contr IS
C1525580|Ankle Fluoroscopy W contrast IS
C1525580|Views^W contrast IS:Find:Pt:Ankle:Doc:XR.fluor
C1525596|Chest X-ray W contrast PO
C1525596|Chest XR W contr PO
C1525596|Views^W contrast Oral:Finding:Point in time:Chest:Document:XR
C1525596|Views^W contrast PO:Find:Pt:Chest:Doc:XR
C1525609|Guidance for biopsy:Find:Pt:Chest>Mediastinum:Doc:CT
C1525609|Guidance for biopsy:Finding:Point in time:Chest>Mediastinum:Document:Computerized Tomography
C1525609|Chest medias CT Bx guid
C1525609|CT Guidance for biopsy of Chest Mediastinum
C1525678|Wrist - left X-ray scaphoid
C1525678|Wrist-L XR Scaphoid
C1525678|Views scaphoid:Find:Pt:Wrist.left:Doc:XR
C1525678|Views scaphoid:Finding:Point in time:Wrist.left:Document:XR
C1525758|Lung parenchyma CT
C1525758|Multisection:Finding:Point in time:Chest>Lung parenchyma:Document:Computerized Tomography
C1525758|Multisection:Find:Pt:Chest>Lung parenchyma:Doc:CT
C1525762|Multisection spectroscopy:Finding:Point in time:To be specified in another part of the message:Narrative:MRI
C1525762|Unspecified body region MRI spectroscopy
C1525762|XXX MRI Spectro
C1525762|Multisection spectroscopy:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1525762|Multisection spectroscopy:Find:Pt:XXX:Doc:MRI
C1524697|Wrist-L MRI W contr IV
C1524697|Wrist - left MRI W contrast IV
C1524697|Multisection^W contrast Intravenous:Finding:Point in time:Wrist.left:Document:MRI
C1524697|Multisection^W contrast IV:Find:Pt:Wrist.left:Doc:MRI
C1525845|Wrist-Bl XR PA+Lat+Obl
C1525845|Wrist - bilateral X-ray PA and lateral and oblique
C1525845|Views PA & lateral & oblique:Finding:Point in time:Wrist.bilateral:Document:XR
C1525845|Views PA & lateral & oblique:Find:Pt:Wrist.bilateral:Doc:XR
C1525801|Spine vessels MRI angiogram
C1525801|Spine ves MRI.Angio
C1525801|Multisection:Find:Pt:Spine vessels:Doc:MRI.angio
C1525801|Multisection:Finding:Point in time:Spine vessels:Document:MRI.angio
C1525804|Spine ves MRI.Angio W contr IV
C1525804|Spine vessels MRI angiogram W contrast IV
C1525804|Multisection^W contrast IV:Find:Pt:Spine vessels:Doc:MRI.angio
C1525804|Multisection^W contrast Intravenous:Finding:Point in time:Spine vessels:Document:MRI.angio
C1525973|Scapula XR Y
C1525973|Scapula X-ray Y
C1525973|View Y:Find:Pt:Scapula:Doc:XR
C1525973|View Y:Finding:Point in time:Scapula:Document:XR
C1526107|Shoulder - right X-ray outlet
C1526107|Should-R XR Outlet
C1526107|View outlet:Finding:Point in time:Shoulder.right:Document:XR
C1526107|View outlet:Find:Pt:Shoulder.right:Doc:XR
C1526108|Should-R XR Lat+Y
C1526108|Shoulder - right X-ray lateral and Y
C1526108|Views lateral & Y:Find:Pt:Shoulder.right:Doc:XR
C1526108|Views lateral & Y:Finding:Point in time:Shoulder.right:Document:XR
C1526049|Lower extremity - right X-ray AP single view standing
C1526049|LE-R XR AP 1V stand
C1526049|View AP^standing:Finding:Point in time:Lower extremity.right:Document:XR
C1526049|View AP^standing:Find:Pt:Lower extremity.right:Doc:XR
C1526056|Knee-R XR AP+Lat+Sunrise+Tunnel
C1526056|Knee - right X-ray AP and lateral and Sunrise and tunnel
C1526056|Views AP & lateral & Sunrise & tunnel:Finding:Point in time:Knee.right:Document:XR
C1526056|Views AP & lateral & Sunrise & tunnel:Find:Pt:Knee.right:Doc:XR
C1526070|Knee-R XR Lat stand
C1526070|Knee - right X-ray lateral standing
C1526070|View lateral^standing:Finding:Point in time:Knee.right:Document:XR
C1526070|View lateral^standing:Find:Pt:Knee.right:Doc:XR
C1526085|Brst-R Mam Mag+Spot
C1526085|Breast - right Mammogram magnification and spot
C1526085|Views magnification & spot:Finding:Point in time:Breast.right:Document:Mam
C1526085|Views magnification & spot:Find:Pt:Breast.right:Doc:Mam
C1526167|Spine X-ray Single view
C1526167|Spine XR 1V
C1526167|View 1:Finding:Point in time:Spine:Document:XR
C1526167|View 1:Find:Pt:Spine:Doc:XR
C1526168|Spine X-ray 4 views
C1526168|Spine XR 4V
C1526168|Views 4:Find:Pt:Spine:Doc:XR
C1526168|Views 4:Finding:Point in time:Spine:Document:XR
C1524270|Sternoclavicular Joint X-ray 3 views
C1524270|SC joint XR 3V
C1524270|Views 3:Find:Pt:Sternoclavicular joint:Doc:XR
C1524270|Views 3:Finding:Point in time:Sternoclavicular joint:Document:XR
C1526242|Upper extremity arteries Fluoroscopic angiogram W contrast IA
C1526242|UE aa XRA W contr IA
C1526242|Views^W contrast Intra-arterial:Finding:Point in time:Upper extremity arteries:Document:XR.fluor.angio
C1526242|Views^W contrast IA:Find:Pt:Upper extremity arteries:Doc:XR.fluor.angio
C1525134|C+T+L-spine XR
C1525134|Spine Cervical and Thoracic and Lumbar X-ray
C1525134|Views:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:XR
C1525134|Views:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:XR
C1526257|Chest wall US
C1526257|Multisection:Find:Pt:Chest wall:Doc:US
C1526257|Multisection:Finding:Point in time:Chest wall:Document:Ultrasound
C1526266|US Guidance for core needle percutaneous biopsy of Breast - right
C1526266|Brst-R US PC Bx CN guid
C1526266|Guidance for percutaneous biopsy.core needle:Find:Pt:Breast.right:Doc:US
C1526266|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast.right:Document:Ultrasound
C1524716|LE-L US
C1524716|Lower extremity - left US
C1524716|Multisection:Find:Pt:Lower extremity.left:Doc:US
C1524716|Multisection:Finding:Point in time:Lower extremity.left:Document:Ultrasound
C1526283|Lower extremity - right US limited
C1526283|LE-R US Ltd
C1526283|Multisection limited:Find:Pt:Lower extremity.right:Doc:US
C1526283|Multisection limited:Finding:Point in time:Lower extremity.right:Document:Ultrasound
C1508083|Abdomen X-ray left posterior oblique
C1508083|Abd XR L-Post Obl
C1508083|View L-posterior oblique:Find:Pt:Abdomen:Doc:XR
C1508083|View L-posterior oblique:Finding:Point in time:Abdomen:Document:XR
C1526324|Wrist XR Scaphoid
C1526324|Wrist X-ray scaphoid
C1526324|Views scaphoid:Finding:Point in time:Wrist:Document:XR
C1526324|Views scaphoid:Find:Pt:Wrist:Doc:XR
C1524484|Ankle-R MRI W contr IV
C1524484|Ankle - right MRI W contrast IV
C1524484|Multisection^W contrast IV:Find:Pt:Ankle.right:Doc:MRI
C1524484|Multisection^W contrast Intravenous:Finding:Point in time:Ankle.right:Document:MRI
C1524879|Upper arm - right CT WO contrast
C1524879|Upper arm-R CT WO contr
C1524879|Multisection^WO contrast:Find:Pt:Upper arm.right:Doc:CT
C1524879|Multisection^WO contrast:Finding:Point in time:Upper arm.right:Document:Computerized Tomography
C1524885|UE joint MRI WO contr
C1524885|Multisection^WO contrast:Find:Pt:Upper extremity.joint:Doc:MRI
C1524885|Multisection^WO contrast:Finding:Point in time:Upper extremity.joint:Document:MRI
C1524885|Upper extremity.joint MRI WO contrast
C1524534|Forearm-R MRI W contr IV
C1524534|Forearm - right MRI W contrast IV
C1524534|Multisection^W contrast Intravenous:Finding:Point in time:Forearm.right:Document:MRI
C1524534|Multisection^W contrast IV:Find:Pt:Forearm.right:Doc:MRI
C1524538|Hand-L MRI W contr IV
C1524538|Hand - left MRI W contrast IV
C1524538|Multisection^W contrast IV:Find:Pt:Hand.left:Doc:MRI
C1524538|Multisection^W contrast Intravenous:Finding:Point in time:Hand.left:Document:MRI
C1524539|Hand-R CT W contr IV
C1524539|Hand - right CT W contrast IV
C1524539|Multisection^W contrast Intravenous:Finding:Point in time:Hand.right:Document:Computerized Tomography
C1524539|Multisection^W contrast IV:Find:Pt:Hand.right:Doc:CT
C1524170|Hip-L MRI W contr IV
C1524170|Hip - left MRI W contrast IV
C1524170|Multisection^W contrast IV:Find:Pt:Hip.left:Doc:MRI
C1524170|Multisection^W contrast Intravenous:Finding:Point in time:Hip.left:Document:MRI
C1524896|Larynx CT WO contr
C1524896|Larynx CT WO contrast
C1524896|Multisection^WO contrast:Finding:Point in time:Neck>Larynx:Document:Computerized Tomography
C1524896|Multisection^WO contrast:Find:Pt:Neck>Larynx:Doc:CT
C1524899|Neck CT WO contrast
C1524899|Neck CT WO contr
C1524899|Multisection^WO contrast:Find:Pt:Neck:Doc:CT
C1524899|Multisection^WO contrast:Finding:Point in time:Neck:Document:Computerized Tomography
C1524902|Post fossa CT WO contr
C1524902|Posterior fossa CT WO contrast
C1524902|Multisection^WO contrast:Find:Pt:Posterior fossa:Doc:CT
C1524902|Multisection^WO contrast:Finding:Point in time:Posterior fossa:Document:Computerized Tomography
C1524943|Finger fourth X-ray lateral
C1524943|Finger.4th XR Lat
C1524943|View lateral:Finding:Point in time:Finger.fourth:Document:XR
C1524943|View lateral:Find:Pt:Finger.fourth:Doc:XR
C1524296|UE CT Bx guid
C1524296|CT Guidance for biopsy of Upper extremity
C1524296|Guidance for biopsy:Find:Pt:Upper extremity:Doc:CT
C1524296|Guidance for biopsy:Finding:Point in time:Upper extremity:Document:Computerized Tomography
C1524603|Ankle-L CT WO+W contr IV
C1524603|Ankle - left CT WO and W contrast IV
C1524603|Multisection^WO & W contrast IV:Find:Pt:Ankle.left:Doc:CT
C1524603|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ankle.left:Document:Computerized Tomography
C1524127|Multisection^WO & W contrast IV:Find:Pt:Breast.right:Doc:MRI
C1524127|Breast - right MRI WO and W contrast IV
C1524127|Brst-R MRI WO+W contr IV
C1524127|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast.right:Document:MRI
C1524964|Hand X-ray oblique single view
C1524964|Hand XR Obl 1V
C1524964|View oblique:Finding:Point in time:Hand:Document:XR
C1524964|View oblique:Find:Pt:Hand:Doc:XR
C1524981|SIJ-Bl XR
C1524981|Sacroiliac joint - bilateral X-ray
C1524981|Views:Find:Pt:Sacroiliac joint.bilateral:Doc:XR
C1524981|Views:Finding:Point in time:Sacroiliac joint.bilateral:Document:XR
C1524989|Abdomen X-ray 2 views
C1524989|Abd XR 2V
C1524989|Views 2:Finding:Point in time:Abdomen:Document:XR
C1524989|Views 2:Find:Pt:Abdomen:Doc:XR
C1524333|L-spine CT PC Vertebroplasty guid
C1524333|Guidance for percutaneous vertebroplasty:Find:Pt:Spine.lumbar:Doc:CT
C1524333|Guidance for percutaneous vertebroplasty:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1524333|CT Guidance for percutaneous vertebroplasty of Lumbar spine
C1524336|CT Guidance for placement of radiation therapy fields in Unspecified body region
C1524336|XXX CT RT fields plac guid
C1524336|Guidance for placement of radiation therapy fields:Find:Pt:XXX:Doc:CT
C1524336|Guidance for placement of radiation therapy fields:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1524627|Elbow-L XR 3V
C1524627|Elbow - left X-ray 3 views
C1524627|Views 3:Find:Pt:Elbow.left:Doc:XR
C1524627|Views 3:Finding:Point in time:Elbow.left:Document:XR
C1524640|Ribs - left X-ray 3 views
C1524640|Ribs-L XR 3V
C1524640|Views 3:Finding:Point in time:Ribs.left:Document:XR
C1524640|Views 3:Find:Pt:Ribs.left:Doc:XR
C1524996|Elbow X-ray 2 views
C1524996|Elbow XR 2V
C1524996|Views 2:Finding:Point in time:Elbow:Document:XR
C1524996|Views 2:Find:Pt:Elbow:Doc:XR
C1524999|Lower extremity X-ray 2 views
C1524999|LE XR 2V
C1524999|Views 2:Find:Pt:Lower extremity:Doc:XR
C1524999|Views 2:Finding:Point in time:Lower extremity:Document:XR
C1524158|Radius+Ulna-L XR 2V
C1524158|Radius - left and Ulna.left X-ray 2 views
C1524158|Views 2:Finding:Point in time:Radius.left+Ulna.left:Document:XR
C1524158|Views 2:Find:Pt:Radius.left+Ulna.left:Doc:XR
C1524367|Lower extremity - bilateral CT
C1524367|LE-Bl CT
C1524367|Multisection:Find:Pt:Lower extremity.bilateral:Doc:CT
C1524367|Multisection:Finding:Point in time:Lower extremity.bilateral:Document:Computerized Tomography
C1524732|Ft-R MRI WO+W contr IV
C1524732|Foot - right MRI WO and W contrast IV
C1524732|Multisection^WO & W contrast Intravenous:Finding:Point in time:Foot.right:Document:MRI
C1524732|Multisection^WO & W contrast IV:Find:Pt:Foot.right:Doc:MRI
C1525027|Coccyx XR AP+Lat
C1525027|Coccyx X-ray AP and lateral
C1525027|Views AP & lateral:Finding:Point in time:Coccyx:Document:XR
C1525027|Views AP & lateral:Find:Pt:Coccyx:Doc:XR
C1525062|Elbow-Bl XR AP+Lat+Obl
C1525062|Elbow - bilateral X-ray AP and lateral and oblique
C1525062|Views AP & lateral & oblique:Find:Pt:Elbow.bilateral:Doc:XR
C1525062|Views AP & lateral & oblique:Finding:Point in time:Elbow.bilateral:Document:XR
C1527039|Hand CT
C1527039|Multisection:Find:Pt:Hand:Doc:CT
C1527039|Multisection:Finding:Point in time:Hand:Document:Computerized Tomography
C1524400|Hrt MRI.Angio
C1524400|Heart MRI angiogram
C1524400|Multisection:Find:Pt:Heart:Doc:MRI.angio
C1524400|Multisection:Finding:Point in time:Heart:Document:MRI.angio
C1524421|Kidney XRTomo
C1524421|Kidney X-ray tomograph
C1524421|Multisection:Find:Pt:Kidney:Doc:XR.tomo
C1524421|Multisection:Finding:Point in time:Kidney:Document:XR.tomo
C1525070|Radius+Ulna-Bl XR Obl
C1525070|Radius - bilateral and Ulna - bilateral X-ray oblique
C1525070|Views oblique:Find:Pt:Radius.bilateral+Ulna.bilateral:Doc:XR
C1525070|Views oblique:Finding:Point in time:Radius.bilateral+Ulna.bilateral:Document:XR
C1525075|Mandible X-ray oblique
C1525075|Mandible XR Obl
C1525075|Views oblique:Find:Pt:Mandible:Doc:XR
C1525075|Views oblique:Finding:Point in time:Mandible:Document:XR
C1525084|Hand-Bl XR PA+Lat+Obl
C1525084|Hand - bilateral X-ray PA and lateral and oblique
C1525084|Views PA & lateral & oblique:Find:Pt:Hand.bilateral:Doc:XR
C1525084|Views PA & lateral & oblique:Finding:Point in time:Hand.bilateral:Document:XR
C1525085|Hand-L XR PA+Lat+Obl
C1525085|Hand - left X-ray PA and lateral and oblique
C1525085|Views PA & lateral & oblique:Find:Pt:Hand.left:Doc:XR
C1525085|Views PA & lateral & oblique:Finding:Point in time:Hand.left:Document:XR
C1525092|Fem ves+Popliteal a XRA Atherect W contr
C1525092|Femoral vessel and Popliteal artery Fluoroscopic angiogram Atherectomy W contrast
C1525092|Atherectomy^W contrast:Finding:Point in time:Femoral vessel+Popliteal artery:Document:XR.fluor.angio
C1525092|Atherectomy^W contrast:Find:Pt:Femoral vessel+Popliteal artery:Doc:XR.fluor.angio
C1830204|Upper extremity vessels US.doppler limited
C1830204|UE ves DOP Ltd
C1830204|Multisection limited:Find:Pt:Upper extremity vessels:Doc:US.doppler
C1830204|Multisection limited:Finding:Point in time:Upper extremity vessels:Document:Ultrasound.doppler
C1830251|Breast - unilateral Mammogram diagnostic
C1830251|Brst-UL Mam Dx
C1830251|Views diagnostic:Find:Pt:Breast.unilateral:Doc:Mam
C1830251|Views diagnostic:Finding:Point in time:Breast.unilateral:Document:Mam
C1831069|Hand - right X-ray GE 3 views
C1831069|Hand-R XR GE 3V
C1831069|Views GE 3:Find:Pt:Hand.right:Doc:XR
C1831069|Views GE 3:Finding:Point in time:Hand.right:Document:XR
C1715417|PV shunt RI for Pat W Tc99mMAA Inj
C1715417|Peritoneovenous shunt Scan for patency W Tc-99m MAA inj
C1715417|Views for shunt patency^W Tc-99m MAA inj:Find:Pt:Peritoneovenous shunt:Doc:Radnuc
C1715417|Views for shunt patency^W Tc-99m MAA inj:Finding:Point in time:Peritoneovenous shunt:Document:Radnuc
C1715495|Upper extremity vessel graft - bilateral US.doppler
C1715495|UE ves graft-Bl DOP
C1715495|Multisection:Find:Pt:Upper extremity vessel graft.bilateral:Doc:US.doppler
C1715495|Multisection:Finding:Point in time:Upper extremity vessel graft.bilateral:Document:Ultrasound.doppler
C1635662|Prostate MRI W endorectal coil
C1635662|Multisection^W endorectal coil:Finding:Point in time:Prostate:Document:MRI
C1635662|Multisection^W endorectal coil:Find:Pt:Prostate:Doc:MRI
C1635007|Kney XR (AP stand)+(Lat hyperext)
C1635007|Knee X-ray (AP^standing) and (lateral^W hyperextension)
C1635007|Views (AP^standing) & (lateral^W hyperextension):Find:Pt:Knee:Doc:XR
C1635007|Views (AP^standing) & (lateral^W hyperextension):Finding:Point in time:Knee:Document:XR
C1714794|Multisection^WO & W contrast IV:Find:Pt:Spine.cervical+Spine.thoracic:Doc:MRI
C1714794|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.cervical+Spine.thoracic:Document:MRI
C1714794|Spine Cervical and Spine Thoracic MRI WO and W contrast IV
C1714794|C+T-spine MRI WO+W contr IV
C1714796|Orbit vessels MRI angiogram WO and W contrast IV
C1714796|Orbit ves MRI.Angio WO+W contr IV
C1714796|Multisection^WO & W contrast IV:Find:Pt:Orbit vessels:Doc:MRI.angio
C1714796|Multisection^WO & W contrast Intravenous:Finding:Point in time:Orbit vessels:Document:MRI.angio
C1714797|Views^during electroconvulsive shock treatment:Finding:Point in time:Heart:Narrative:Radnuc
C1714797|Deprecated Hrt RI During EST
C1714797|Views^during electroconvulsive shock treatment:Find:Pt:Heart:Nar:Radnuc
C1714797|Deprecated Heart Scan during electroconvulsive shock treatment
C1714787|Ankle-R MRI Dyn W contr IV
C1714787|Ankle - right MRI dynamic W contrast IV
C1714787|Multisection dynamic^W contrast IV:Find:Pt:Ankle.right:Doc:MRI
C1714787|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Ankle.right:Document:MRI
C1705865|Deprecated Finger.3rd-L XR GE 3V
C1705865|Deprecated Finger third Left X-ray GE 3 views
C1705865|Views GE 3:Find:Pt:Finger.third.left:Nar:XR
C1705865|Views GE 3:Finding:Point in time:Finger.third.left:Narrative:XR
C1715020|RI for ETr Mul Areas W I-131 mIBG IV
C1715020|Scan for endocrine tumor multiple areas W I-131 MIBG IV
C1715020|Views for endocrine tumor multiple areas^W I-131 MIBG IV:Find:Pt:^Patient:Doc:Radnuc
C1715020|Views for endocrine tumor multiple areas^W I-131 MIBG Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1715097|Multisection^WO & W contrast IV:Find:Pt:Brain+Internal auditory canal:Doc:MRI
C1715097|Brain and Internal auditory canal MRI WO and W contrast IV
C1715097|Brain+IAC MRI WO+W contr IV
C1715097|Multisection^WO & W contrast Intravenous:Finding:Point in time:Brain+Internal auditory canal:Document:MRI
C1631254|Liver Scan flow
C1631254|Liver RI Flow W RNC IV
C1631254|Views flow^W radionuclide IV:Find:Pt:Liver:Doc:Radnuc
C1631254|Views flow^W radionuclide Intravenous:Finding:Point in time:Liver:Document:Radnuc
C1644168|Multisection^WO & W contrast IV:Find:Pt:Extremity:Doc:CT
C1644168|Extremity CT WO and W contrast IV
C1644168|Multisection^WO & W contrast Intravenous:Finding:Point in time:Extremity:Document:Computerized Tomography
C1644168|Extr CT WO+W contr IV
C1642592|Knee-R XR port
C1642592|Knee - right X-ray portable
C1642592|Views portable:Find:Pt:Knee.right:Doc:XR
C1642592|Views portable:Finding:Point in time:Knee.right:Document:XR
C1977323|Hrt SPECT PF W ADE+Tc99mMIBI IV
C1977323|Heart SPECT perfusion W adenosine and W Tc-99m Sestamibi IV
C1977323|Multisection perfusion^W adenosine & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1977323|Multisection perfusion^W adenosine & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1953965|Clavicle - left MRI WO contrast
C1953965|Clavicle-L MRI WO contr
C1953965|Multisection^WO contrast:Find:Pt:Clavicle.left:Doc:MRI
C1953965|Multisection^WO contrast:Finding:Point in time:Clavicle.left:Document:MRI
C3169526|Head a+Neck a-L-R XRA W contr IA
C3169526|Head artery.right+Neck artery.right Fluoroscopic angiogram W contrast IA
C3169526|Views^W contrast IA:Find:Pt:Head artery.right+Neck artery.right:Doc:XR.fluor.angio
C3169526|Views^W contrast Intra-arterial:Finding:Point in time:Head artery.right+Neck artery.right:Document:XR.fluor.angio
C3533551|Guidance for repair of CVA catheter without port or pump:Finding:Point in time:Central vein:Document:XR.fluor
C3533551|Centl v Flr CVA cath WO pump repair guid
C3533551|Guidance for repair of CVA catheter without port or pump:Find:Pt:Central vein:Doc:XR.fluor
C3533551|Fluoroscopy Guidance for repair of CVA catheter without port or pump of Central vein
C3533550|L-spine Flr Kyphoplasty guid
C3533550|Guidance for kyphoplasty:Finding:Point in time:Spine.lumbar:Document:XR.fluor
C3533550|Guidance for kyphoplasty:Find:Pt:Spine.lumbar:Doc:XR.fluor
C3533550|Fluoroscopy Guidance for kyphoplasty of Lumbar spine
C3262949|Fluoroscopy Guidance for needle biopsy of Pancreas
C3262949|Pancreas Flr Bx needle guid
C3262949|Guidance for biopsy.needle:Finding:Point in time:Pancreas:Document:XR.fluor
C3262949|Guidance for biopsy.needle:Find:Pt:Pancreas:Doc:XR.fluor
C3263048|Scrotum+Test SPECT Flow W RNC IV
C3263048|Scrotum and Testicle SPECT flow
C3263048|Multisection flow^W radionuclide Intravenous:Finding:Point in time:Scrotum+Testicle:Document:Radnuc.SPECT
C3263048|Multisection flow^W radionuclide IV:Find:Pt:Scrotum+Testicle:Doc:Radnuc.SPECT
C3263062|Popliteal a XRA W contr IA
C3263062|Popliteal artery Fluoroscopic angiogram W contrast IA
C3263062|Views^W contrast Intra-arterial:Finding:Point in time:Popliteal artery:Document:XR.fluor.angio
C3263062|Views^W contrast IA:Find:Pt:Popliteal artery:Doc:XR.fluor.angio
C3263074|Shoulder - right X-ray AP and Grashey and axillary
C3263074|Should-R XR AP+Grashey+Ax
C3263074|Views AP & Grashey & axillary:Find:Pt:Shoulder.right:Doc:XR
C3263074|Views AP & Grashey & axillary:Finding:Point in time:Shoulder.right:Document:XR
C3263076|Sacrum X-ray standing
C3263076|Sacrum XR stand
C3263076|Views^standing:Find:Pt:Sacrum:Doc:XR
C3263076|Views^standing:Finding:Point in time:Sacrum:Document:XR
C3263081|Skull XR AP 1V
C3263081|Skull X-ray AP single view
C3263081|View AP:Find:Pt:Skull:Doc:XR
C3263081|View AP:Finding:Point in time:Skull:Document:XR
C3261717|Unspecified body region US.doppler limited
C3261717|XXX DOP Ltd
C3261717|Multisection limited:Find:Pt:XXX:Doc:US.doppler
C3261717|Multisection limited:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound.doppler
C3263104|Wrist XR Ulnar dev
C3263104|Wrist X-ray ulnar deviation
C3263104|Views ulnar deviation:Find:Pt:Wrist:Doc:XR
C3263104|Views ulnar deviation:Finding:Point in time:Wrist:Document:XR
C3263215|Extremity vessels Left US.doppler
C3263215|Extr ves-L DOP
C3263215|Multisection:Find:Pt:Extremity vessels.left:Doc:US.doppler
C3263215|Multisection:Finding:Point in time:Extremity vessels.left:Document:Ultrasound.doppler
C3262897|Fluoroscopy Guidance for biopsy of Pelvis
C3262897|Pelvis Flr Bx guid
C3262897|Guidance for biopsy:Finding:Point in time:Pelvis:Document:XR.fluor
C3262897|Guidance for biopsy:Find:Pt:Pelvis:Doc:XR.fluor
C0942160|Deprecated DEXA
C0942160|Views:Find:Pt:Radius+Ulna.right:Nar:XR.DEXA
C0942160|Views:Finding:Point in time:Radius+Ulna.right:Narrative:XR.DEXA
C0942160|Deprecated Radius & Ulna right DEXA Bone density views
C0942188|TO ves-Bl MRI.Angio W contr IV
C0942188|Thoracic outlet vessels - bilateral MRI angiogram W contrast IV
C0942188|Multisection^W contrast Intravenous:Finding:Point in time:Thoracic outlet vessels.bilateral:Document:MRI.angio
C0942188|Multisection^W contrast IV:Find:Pt:Thoracic outlet vessels.bilateral:Doc:MRI.angio
C0942192|Multisection^WO & W contrast IV:Find:Pt:Ankle.bilateral:Doc:MRI
C0942192|Ankle-Bl MRI WO+W contr IV
C0942192|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ankle.bilateral:Document:MRI
C0942192|Ankle - bilateral MRI WO and W contrast IV
C0942197|Elbow - bilateral MRI WO and W contrast IV
C0942197|Multisection^WO & W contrast Intravenous:Finding:Point in time:Elbow.bilateral:Document:MRI
C0942197|Multisection^WO & W contrast IV:Find:Pt:Elbow.bilateral:Doc:MRI
C0942197|Elbow-Bl MRI WO+W contr IV
C0942217|TO-R MRI
C0942217|Thoracic outlet - right MRI
C0942217|Multisection:Finding:Point in time:Thoracic outlet.right:Document:MRI
C0942217|Multisection:Find:Pt:Thoracic outlet.right:Doc:MRI
C0942233|UE-L MRI
C0942233|Upper extremity - left MRI
C0942233|Multisection:Finding:Point in time:Upper extremity.left:Document:MRI
C0942233|Multisection:Find:Pt:Upper extremity.left:Doc:MRI
C0942246|Hip-Bl US
C0942246|Hip - bilateral US
C0942246|Multisection:Finding:Point in time:Hip.bilateral:Document:Ultrasound
C0942246|Multisection:Find:Pt:Hip.bilateral:Doc:US
C0942251|Knee - bilateral MRI
C0942251|Knee-Bl MRI
C0942251|Multisection:Find:Pt:Knee.bilateral:Doc:MRI
C0942251|Multisection:Finding:Point in time:Knee.bilateral:Document:MRI
C0942253|Knee - right MRI
C0942253|Knee-R MRI
C0942253|Multisection:Find:Pt:Knee.right:Doc:MRI
C0942253|Multisection:Finding:Point in time:Knee.right:Document:MRI
C0945332|Brst-Bl Mam Bx Str Guid
C0945332|Guidance for stereotactic biopsy:Find:Pt:Breast.bilateral:Doc:Mam
C0945332|Guidance for stereotactic biopsy:Finding:Point in time:Breast.bilateral:Document:Mam
C0945332|Mammogram Guidance for stereotactic biopsy of Breast - bilateral
C0942290|Vein-R XRA Atherect guid W contr IV
C0942290|Fluoroscopic angiogram Guidance for atherectomy of Vein - right-- W contrast IV
C0942290|Guidance for atherectomy^W contrast IV:Find:Pt:Vein.right:Doc:XR.fluor.angio
C0942290|Guidance for atherectomy^W contrast Intravenous:Finding:Point in time:Vein.right:Document:XR.fluor.angio
C0942322|Mammogram Guidance for core needle percutaneous biopsy of Breast - right
C0942322|Brst-R Mam PC Bx CN guid
C0942322|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast.right:Document:Mam
C0942322|Guidance for percutaneous biopsy.core needle:Find:Pt:Breast.right:Doc:Mam
C0942327|US Guidance for biopsy of Kidney - right
C0942327|Kidney-R US Bx guid
C0942327|Guidance for biopsy:Find:Pt:Kidney.right:Doc:US
C0942327|Guidance for biopsy:Finding:Point in time:Kidney.right:Document:Ultrasound
C0942335|Wrist+Hand-Bl XR Bone Age
C0942335|Wrist - bilateral and Hand - bilateral X-ray bone age
C0942335|Views bone age:Finding:Point in time:Wrist.bilateral+Hand.bilateral:Document:XR
C0942335|Views bone age:Find:Pt:Wrist.bilateral+Hand.bilateral:Doc:XR
C0942353|Tibial artery - bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C0942353|Tibl a-Bl XRA Angpsty W contr IA
C0942353|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibial artery.bilateral:Document:XR.fluor.angio
C0942353|Angioplasty^W contrast IA:Find:Pt:Tibial artery.bilateral:Doc:XR.fluor.angio
C0942358|Hand-Bl XR 3V
C0942358|Hand - bilateral X-ray 3 views
C0942358|Views 3:Find:Pt:Hand.bilateral:Doc:XR
C0942358|Views 3:Finding:Point in time:Hand.bilateral:Document:XR
C0882066|Petrous part of temporal bone CT
C0882066|Petr part temp bone CT
C0882066|Multisection:Find:Pt:Petrous part of temporal bone:Doc:CT
C0882066|Multisection:Finding:Point in time:Petrous part of temporal bone:Document:Computerized Tomography
C0882085|Salivary gland Fluoroscopy W contrast intra salivary duct
C0882085|Salivary gland Flr W contr intra SD
C0882085|Views^W contrast intra salivary duct:Find:Pt:Salivary gland:Doc:XR.fluor
C0882085|Views^W contrast intra salivary duct:Finding:Point in time:Salivary gland:Document:XR.fluor
C0882088|Shoulder MRI
C0882088|Should MRI
C0882088|Multisection:Finding:Point in time:Shoulder:Narrative:MRI
C0882088|Multisection:Finding:Point in time:Shoulder:Document:MRI
C0882088|Multisection:Find:Pt:Shoulder:Doc:MRI
C0944155|Skull X-ray Single view
C0944155|Skull XR 1V
C0944155|View 1:Find:Pt:Skull:Doc:XR
C0944155|View 1:Finding:Point in time:Skull:Document:XR
C0882109|Spine Flr W contr ID
C0882109|Spine Fluoroscopy W contrast intradisc
C0882109|Views^W contrast intradisc:Find:Pt:Spine:Doc:XR.fluor
C0882109|Views^W contrast intradisc:Finding:Point in time:Spine:Document:XR.fluor
C0882110|T+L-spine XR Scoli W FE
C0882110|Views scoliosis^W flexion & W extension:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C0882110|Spine Thoracic and Lumbar X-ray scoliosis W flexion and W extension
C0882110|Views scoliosis^W flexion & W extension:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C0882113|C-spine CT W contr IV
C0882113|Multisection^W contrast Intravenous:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C0882113|Multisection^W contrast IV:Find:Pt:Spine.cervical:Doc:CT
C0882113|Cervical spine CT W contrast IV
C0882130|Multisection:Finding:Point in time:Spine.lumbar:Narrative:MRI
C0882130|L-spine MRI
C0882130|Multisection:Find:Pt:Spine.lumbar:Doc:MRI
C0882130|Multisection:Finding:Point in time:Spine.lumbar:Document:MRI
C0882130|Lumbar spine MRI
C2607991|L-spine XR
C2607991|Views:Find:Pt:Spine.lumbar:Doc:XR
C2607991|Views:Finding:Point in time:Spine.lumbar:Document:XR
C2607991|Lumbar spine X-ray
C0882140|T-spine CT W contr IV
C0882140|Multisection^W contrast IV:Find:Pt:Spine.thoracic:Doc:CT
C0882140|Multisection^W contrast Intravenous:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C0882140|Thoracic spine CT W contrast IV
C0882560|Views:Finding:Point in time:Toes:Narrative:XR
C0882560|Toes X-ray
C0882560|Toes XR
C0882560|Views:Finding:Point in time:Toes:Document:XR
C0882560|Views:Find:Pt:Toes:Doc:XR
C0882177|Deprecated Bladder+Urethra Flr W vdg
C0882177|Deprecated Urinary Bladder & Urethra Fluoroscopy W voiding
C0882177|Views^W voiding:Find:Pt:Urinary bladder+Urethra:Nar:XR.fluor
C0882177|Views^W voiding:Finding:Point in time:Urinary bladder+Urethra:Narrative:XR.fluor
C0882186|Abd aa XRA W contr IA
C0882186|Views^W contrast Intra-arterial:Finding:Point in time:Abdominal arteries:Document:XR.fluor.angio
C0882186|Views^W contrast IA:Find:Pt:Abdominal arteries:Doc:XR.fluor.angio
C0882186|Abdominal Arteries Fluoroscopic angiogram W contrast IA
C0882208|XXX CT Radiosurg guid W contr IV
C0882208|CT Guidance for radiosurgery of Unspecified body region-- W contrast IV
C0882208|Guidance for radiosurgery^W contrast IV:Find:Pt:XXX:Doc:CT
C0882208|Guidance for radiosurgery^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882563|Multisection:Finding:Point in time:To be specified in another part of the message:Narrative:MRI
C0882563|Unspecified body region MRI
C0882563|XXX MRI
C0882563|Multisection:Find:Pt:XXX:Doc:MRI
C0882563|Multisection:Finding:Point in time:To be specified in another part of the message:Document:MRI
C0942103|Spinal a-Bl XRA W contr IA
C0942103|Spinal artery - bilateral Fluoroscopic angiogram W contrast IA
C0942103|Views^W contrast IA:Find:Pt:Spinal artery.bilateral:Doc:XR.fluor.angio
C0942103|Views^W contrast Intra-arterial:Finding:Point in time:Spinal artery.bilateral:Document:XR.fluor.angio
C0881791|Stent Fluoroscopy W contrast intra stent
C0881791|Stent Flr W contr intra stnt
C0881791|Views^W contrast intra stent:Finding:Point in time:To be specified in another part of the message stent:Document:XR.fluor
C0881791|Views^W contrast intra stent:Find:Pt:XXX stent:Doc:XR.fluor
C0881807|AVF XRA Atherect W contr IV
C0881807|AV fistula Fluoroscopic angiogram Atherectomy W contrast IV
C0881807|Atherectomy^W contrast IV:Find:Pt:AV fistula:Doc:XR.fluor.angio
C0881807|Atherectomy^W contrast Intravenous:Finding:Point in time:AV fistula:Document:XR.fluor.angio
C0881815|Bone X-ray during surgery
C0881815|Bone XR in Surg
C0881815|Views^during surgery:Finding:Point in time:Bone.To be specified in another part of the message:Document:XR
C0881815|Views^during surgery:Find:Pt:Bone.XXX:Doc:XR
C0881824|Multisection^WO & W contrast Intravenous:Finding:Point in time:Brain:Document:MRI
C0881824|Brain MRI WO+W contr IV
C0881824|Brain MRI WO and W contrast IV
C0881824|Multisection^WO & W contrast IV:Find:Pt:Brain:Doc:MRI
C0881852|Cath Flr Patency Ck W contr via cath
C0881852|Catheter Fluoroscopy Patency check W contrast via catheter
C0881852|Patency check^W contrast via catheter:Find:Pt:Catheter.XXX:Doc:XR.fluor
C0881852|Patency check^W contrast via catheter:Finding:Point in time:Catheter.To be specified in another part of the message:Document:XR.fluor
C0881871|Chest XR PA+Lat+R-or L-Obl Upr
C0881871|Chest X-ray PA and lateral and right or-left oblique upright
C0881871|Views PA & lateral & R-or-L-oblique upright:Find:Pt:Chest:Doc:XR
C0881871|Views PA & lateral & R-or-L-oblique upright:Finding:Point in time:Chest:Document:XR
C0881889|Views:Finding:Point in time:Clavicle:Narrative:XR
C0881889|Clavicle XR
C0881889|Clavicle X-ray
C0881889|Views:Finding:Point in time:Clavicle:Document:XR
C0881889|Views:Find:Pt:Clavicle:Doc:XR
C0881934|Gastrointestine upper Fluoroscopy Single view W contrast PO
C0881934|UGI Flr 1V W contr PO
C0881934|View 1^W contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C0881934|View 1^W contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C0881948|Views^W radionuclide Intravenous:Finding:Point in time:Brain:Narrative:Radnuc
C0881948|Brain RI W RNC IV
C0881948|Brain Scan
C0881948|Views^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc
C0881948|Views^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc
C0881990|Kidney - bilateral X-ray tomograph W contrast IV
C0881990|Multisection^W contrast IV:Find:Pt:Kidney.bilateral:Doc:XR.tomo
C0881990|Multisection^W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:XR.tomo
C0881990|Kdny-Bl XRTomo W contr IV
C1114485|Sinuses MRI WO and W contrast IV
C1114485|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sinuses:Document:MRI
C1114485|Sinuses MRI WO+W contr IV
C1114485|Multisection^WO & W contrast IV:Find:Pt:Sinuses:Doc:MRI
C1114501|Ankle MRI WO contrast
C1114501|Ankle MRI WO contr
C1114501|Multisection^WO contrast:Finding:Point in time:Ankle:Document:MRI
C1114501|Multisection^WO contrast:Find:Pt:Ankle:Doc:MRI
C1114593|Knee X-ray 3 views
C1114593|Knee XR 3V
C1114593|Views 3:Find:Pt:Knee:Doc:XR
C1114593|Views 3:Finding:Point in time:Knee:Document:XR
C1114594|Knee X-ray 4 views
C1114594|Knee XR 4V
C1114594|Views 4:Finding:Point in time:Knee:Document:XR
C1114594|Views 4:Find:Pt:Knee:Doc:XR
C1114660|Aorta+Abd aa MRI.Angio
C1114660|Abdominal Aorta and Arteries MRI angiogram
C1114660|Multisection:Find:Pt:Aorta+Abdominal arteries:Doc:MRI.angio
C1114660|Multisection:Finding:Point in time:Aorta+Abdominal arteries:Document:MRI.angio
C1114662|Celiac ves+SM ves MRI.Angio
C1114662|Celiac vessels and Superior mesenteric Vessels MRI angiogram
C1114662|Multisection:Finding:Point in time:Celiac vessels+Superior mesenteric vessels:Document:MRI.angio
C1114662|Multisection:Find:Pt:Celiac vessels+Superior mesenteric vessels:Doc:MRI.angio
C1114670|UE joint MRI
C1114670|Multisection:Finding:Point in time:Upper extremity.joint:Document:MRI
C1114670|Multisection:Find:Pt:Upper extremity.joint:Doc:MRI
C1114670|Upper extremity.joint MRI
C1114412|CT Guidance for fine needle aspiration of Unspecified body region
C1114412|XXX CT FNA Asp
C1114412|Guidance for aspiration.fine needle:Find:Pt:XXX:Doc:CT
C1114412|Guidance for aspiration.fine needle:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1114425|T-spine CT W contr IT
C1114425|Multisection^W contrast Intrathecal:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C1114425|Multisection^W contrast IT:Find:Pt:Spine.thoracic:Doc:CT
C1114425|Thoracic spine CT W contrast IT
C1543420|Should-L XR AP(w IR+ER)+Ax
C1543420|Shoulder - left X-ray AP (W internal rotation and W external rotation) and axillary
C1543420|Views AP (W internal rotation & W external rotation) & axillary:Finding:Point in time:Shoulder.left:Document:XR
C1543420|Views AP (W internal rotation & W external rotation) & axillary:Find:Pt:Shoulder.left:Doc:XR
C1543431|Should-Bl XR AP(w IR)+West Point
C1543431|Shoulder - bilateral X-ray AP (W internal rotation) and West Point
C1543431|Views AP (W internal rotation) & West Point:Find:Pt:Shoulder.bilateral:Doc:XR
C1543431|Views AP (W internal rotation) & West Point:Finding:Point in time:Shoulder.bilateral:Document:XR
C1543769|Deprecated Views perfusion^at rest & W 99m Tc mibi IV:Find:Pt:Heart:Nar:Radnuc
C1543769|Views perfusion^at rest & W 99m Tc mibi IV:Find:Pt:Heart:Nar:Radnuc
C1543769|Deprecated Heart Scintigraphy perfusion at rest & W Tc-99m Sestamibi IV
C1543769|Deprecated Hrt RI PF
C1543769|Views perfusion^at rest & W 99m Tc mibi Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1543465|Knee-R XR 4V+Obl
C1543465|Knee - right X-ray 4 views and oblique
C1543465|Views 4 & oblique:Find:Pt:Knee.right:Doc:XR
C1543465|Views 4 & oblique:Finding:Point in time:Knee.right:Document:XR
C1543475|Should-R XR AP(w IR+ER)+West Point
C1543475|Shoulder - right X-ray AP (W internal rotation and W external rotation) and West Point
C1543475|Views AP (W internal rotation & W external rotation) & West Point:Finding:Point in time:Shoulder.right:Document:XR
C1543475|Views AP (W internal rotation & W external rotation) & West Point:Find:Pt:Shoulder.right:Doc:XR
C1543779|Hrt RI PF Rest+stress+W Tc99mMIBI IV
C1543779|Heart Scan perfusion at rest and W stress and W Tc-99m Sestamibi IV
C1543779|Views perfusion^at rest & W stress & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543779|Views perfusion^at rest & W stress & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543797|Kidney - bilateral Scan W Tc-99m DTPA IV
C1543797|Views^W Tc-99m DTPA Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1543797|Views^W Tc-99m DTPA IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1543797|Kdny-Bl RI W Tc99mDTPA IV
C1543799|Salivary gland Scan
C1543799|Salivary gland RI W RNC IV
C1543799|Views^W radionuclide IV:Find:Pt:Salivary gland:Doc:Radnuc
C1543799|Views^W radionuclide Intravenous:Finding:Point in time:Salivary gland:Document:Radnuc
C1543802|RI Tum local guid Ltd W RNC IV
C1543802|Scan Guidance for localization of tumor limited
C1543802|Guidance for localization of tumor limited^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C1543802|Guidance for localization of tumor limited^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543890|Hrt RI BP W Stress+W RNC IV
C1543890|Heart Scan blood pool W stress and W radionuclide IV
C1543890|Views blood pool^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543890|Views blood pool^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543918|RI Static for Tumor W Ga-67 IV
C1543918|Views static for tumor^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543918|Views static for tumor^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543918|Scan static for tumor W Ga-67 IV
C1543930|Hrt RI FP+WM+VV W Stress+W RNC IV
C1543930|Heart Scan first pass and wall motion and ventricular volume W stress and W radionuclide IV
C1543930|Views first pass & wall motion & ventricular volume^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543930|Views first pass & wall motion & ventricular volume^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543964|Views for tumor multiple areas^W Tc-99m Sestamibi IV:Find:Pt:^Patient:Doc:Radnuc
C1543964|Scan for tumor multiple areas W Tc-99m Sestamibi IV
C1543964|RI for Tumor Mul Areas W Tc99mMIBI IV
C1543964|Views for tumor multiple areas^W Tc-99m Sestamibi Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1526354|Radius+Ulna DXA T-score BDM
C1526354|Bone density:Tscore:Pt:Radius+Ulna:Qn:XR.DXA
C1526354|Radius and Ulna DXA [T-score] Bone density
C1526354|Bone density:T Score:Point in time:Radius+Ulna:Quantitative:XR.DXA
C1526356|Bone density:Tscore:Pt:Spine.lumbar:Qn:XR.DXA
C1526356|L-spine DXA T-score BDM
C1526356|Bone density:T Score:Point in time:Spine.lumbar:Quantitative:XR.DXA
C1526356|Lumbar spine DXA [T-score] Bone density
C1543173|Spine XR Lat
C1543173|Spine X-ray lateral
C1543173|View lateral:Find:Pt:Spine:Doc:XR
C1543173|View lateral:Finding:Point in time:Spine:Document:XR
C1543600|Vein DOP
C1543600|Vein US.doppler
C1543600|Multisection:Finding:Point in time:Vein:Document:Ultrasound.doppler
C1543600|Multisection:Find:Pt:Vein:Doc:US.doppler
C1543269|Brst.duct Mam W contr intra Dcts
C1543269|Breast duct Mammogram W contrast intra multiple ducts
C1543269|Views^W contrast intra multiple ducts:Finding:Point in time:Breast.duct:Document:Mam
C1543269|Views^W contrast intra multiple ducts:Find:Pt:Breast.duct:Doc:Mam
C1543682|Scan Guidance for abscess localization limited
C1543682|RI Abscess local guid Ltd W RNC IV
C1543682|Guidance for abscess localization limited^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C1543682|Guidance for abscess localization limited^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543693|Brain SPECT W Tc99mHMPAO IV
C1543693|Brain SPECT W Tc-99m HMPAO IV
C1543693|Multisection^W Tc-99m HMPAO IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1543693|Multisection^W Tc-99m HMPAO Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1524256|Should-R XR AP+Ax+Outlet
C1524256|Shoulder - right X-ray AP and axillary and outlet
C1524256|Views AP & axillary & outlet:Finding:Point in time:Shoulder.right:Document:XR
C1524256|Views AP & axillary & outlet:Find:Pt:Shoulder.right:Doc:XR
C1526757|Gastric a-R XRA W contr IA
C1526757|Gastric artery - right Fluoroscopic angiogram W contrast IA
C1526757|Views^W contrast Intra-arterial:Finding:Point in time:Gastric artery.right:Document:XR.fluor.angio
C1526757|Views^W contrast IA:Find:Pt:Gastric artery.right:Doc:XR.fluor.angio
C1543712|Hrt RI W RNC IV
C1543712|Heart Scan
C1543712|Views^W radionuclide Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1543712|Views^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543712|Views^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1526795|Wrist - left X-ray oblique
C1526795|Wrist-L XR Obl
C1526795|Views oblique:Finding:Point in time:Wrist.left:Document:XR
C1526795|Views oblique:Find:Pt:Wrist.left:Doc:XR
C1543417|Ft-L XR AP+Lat stand
C1543417|Foot - left X-ray AP and lateral standing
C1543417|Views AP & lateral^standing:Find:Pt:Foot.left:Doc:XR
C1543417|Views AP & lateral^standing:Finding:Point in time:Foot.left:Document:XR
C1524810|Ankle CT WO contrast
C1524810|Ankle CT WO contr
C1524810|Multisection^WO contrast:Find:Pt:Ankle:Doc:CT
C1524810|Multisection^WO contrast:Finding:Point in time:Ankle:Document:Computerized Tomography
C1524814|Ankle-R MRI WO contr
C1524814|Ankle - right MRI WO contrast
C1524814|Multisection^WO contrast:Find:Pt:Ankle.right:Doc:MRI
C1524814|Multisection^WO contrast:Finding:Point in time:Ankle.right:Document:MRI
C1524454|C-spine CT Ltd W contr IV
C1524454|Multisection limited^W contrast Intravenous:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C1524454|Multisection limited^W contrast IV:Find:Pt:Spine.cervical:Doc:CT
C1524454|Cervical spine CT limited W contrast IV
C1524461|Multisection^W contrast Intrasynovial:Finding:Point in time:Ankle.right:Document:MRI
C1524461|Multisection^W contrast IS:Find:Pt:Ankle.right:Doc:MRI
C1524461|Ankle-R MRI W contr IS
C1524461|Ankle - right MRI W contrast IS
C1524466|Multisection^W contrast Intrasynovial:Finding:Point in time:Hip.right:Document:MRI
C1524466|Multisection^W contrast IS:Find:Pt:Hip.right:Doc:MRI
C1524466|Hip-R MRI W contr IS
C1524466|Hip - right MRI W contrast IS
C1525213|Mastoid X-ray 3 views
C1525213|Mastoid XR 3V
C1525213|Views 3:Find:Pt:Mastoid:Doc:XR
C1525213|Views 3:Finding:Point in time:Mastoid:Document:XR
C1525214|Mastoid XR 4V
C1525214|Mastoid X-ray 4 views
C1525214|Views 4:Finding:Point in time:Mastoid:Document:XR
C1525214|Views 4:Find:Pt:Mastoid:Doc:XR
C1525254|Head ves MRI.Angio WO contr
C1525254|Head vessels MRI angiogram WO contrast
C1525254|Multisection^WO contrast:Finding:Point in time:Head vessels:Document:MRI.angio
C1525254|Multisection^WO contrast:Find:Pt:Head vessels:Doc:MRI.angio
C1525274|Chest and Abdomen MRI W contrast IV
C1525274|Chest+Abd MRI W contr IV
C1525274|Multisection^W contrast Intravenous:Finding:Point in time:Chest+Abdomen:Document:MRI
C1525274|Multisection^W contrast IV:Find:Pt:Chest+Abdomen:Doc:MRI
C1525327|Abdomen X-ray left lateral
C1525327|Abd XR L-Lat
C1525327|View L-lateral:Find:Pt:Abdomen:Doc:XR
C1525327|View L-lateral:Finding:Point in time:Abdomen:Document:XR
C1525336|Knee XR Laurin
C1525336|Knee X-ray Laurin
C1525336|View Laurin:Find:Pt:Knee:Doc:XR
C1525336|View Laurin:Finding:Point in time:Knee:Document:XR
C1525471|Deprecated Calcaneus - bilateral X-ray standing
C1525471|Deprecated Heel-Bl XR stand
C1525471|View^standing:Find:Pt:Calcaneus.bilateral:Doc:XR
C1525471|View^standing:Finding:Point in time:Calcaneus.bilateral:Document:XR
C1525471|Deprecated View^standing:Find:Pt:Calcaneus.bilateral:Doc:XR
C1525525|Should-L XR AP+Y
C1525525|Shoulder - left X-ray AP and Y
C1525525|Views AP & Y:Finding:Point in time:Shoulder.left:Document:XR
C1525525|Views AP & Y:Find:Pt:Shoulder.left:Doc:XR
C1525531|L-spine XR Lat W FE
C1525531|Views lateral^W flexion & W extension:Find:Pt:Spine.lumbar:Doc:XR
C1525531|Views lateral^W flexion & W extension:Finding:Point in time:Spine.lumbar:Document:XR
C1525531|Lumbar spine X-ray lateral W flexion and W extension
C1525553|Knee XR Obl+Sunrise
C1525553|Knee X-ray oblique and Sunrise
C1525553|Views oblique & Sunrise:Find:Pt:Knee:Doc:XR
C1525553|Views oblique & Sunrise:Finding:Point in time:Knee:Document:XR
C1525576|IM a XRA W contr IA
C1525576|Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C1525576|Views^W contrast IA:Find:Pt:Inferior mesenteric artery:Doc:XR.fluor.angio
C1525576|Views^W contrast Intra-arterial:Finding:Point in time:Inferior mesenteric artery:Document:XR.fluor.angio
C1525601|Views^standing:Find:Pt:Calcaneus:Doc:XR
C1525601|Deprecated Heel XR stand
C1525601|Deprecated Calcaneus X-ray standing
C1525601|Views^standing:Finding:Point in time:Calcaneus:Document:XR
C1525602|Views^standing:Finding:Point in time:Calcaneus.left:Document:XR
C1525602|Views^standing:Find:Pt:Calcaneus.left:Doc:XR
C1525602|Deprecated Heel-L XR stand
C1525602|Deprecated Calcaneus - left X-ray standing
C1525650|L-spine+Sacrum+SIJ+Coccyx XR 3V
C1525650|Spine Lumbar and Sacrum and Sacroiliac Joint and Coccyx X-ray 3 views
C1525650|Views 3:Find:Pt:Spine.lumbar+Sacrum+Sacroiliac joint+Coccyx:Doc:XR
C1525650|Views 3:Finding:Point in time:Spine.lumbar+Sacrum+Sacroiliac joint+Coccyx:Document:XR
C1525710|Ac arch+Vertebral a XRA W contr IA
C1525710|Aortic arch and Vertebral artery Fluoroscopic angiogram W contrast IA
C1525710|Views^W contrast IA:Find:Pt:Aortic arch+Vertebral artery:Doc:XR.fluor.angio
C1525710|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Vertebral artery:Document:XR.fluor.angio
C1525746|LE v XRA Angpsty W contr IV
C1525746|Lower extremity vein Fluoroscopic angiogram Angioplasty W contrast IV
C1525746|Angioplasty^W contrast Intravenous:Finding:Point in time:Lower extremity vein:Document:XR.fluor.angio
C1525746|Angioplasty^W contrast IV:Find:Pt:Lower extremity vein:Doc:XR.fluor.angio
C1525751|Wrist - left X-ray tomograph
C1525751|Wrist-L XRTomo
C1525751|Multisection:Find:Pt:Wrist.left:Doc:XR.tomo
C1525751|Multisection:Finding:Point in time:Wrist.left:Document:XR.tomo
C1525786|Wrist-Bl XR 2V
C1525786|Wrist - bilateral X-ray 2 views
C1525786|Views 2:Find:Pt:Wrist.bilateral:Doc:XR
C1525786|Views 2:Finding:Point in time:Wrist.bilateral:Document:XR
C1525849|Breast - left Mammogram spot compression
C1525849|Brst-L Mam Spot Compression
C1525849|Views spot^compression:Finding:Point in time:Breast.left:Document:Mam
C1525849|Views spot^compression:Find:Pt:Breast.left:Doc:Mam
C1525935|Pelvis X-ray 2 views
C1525935|Pelvis XR 2V
C1525935|Views 2:Find:Pt:Pelvis:Doc:XR
C1525935|Views 2:Finding:Point in time:Pelvis:Document:XR
C1525827|Finger third - left X-ray
C1525827|Finger.3rd-L XR
C1525827|Views:Find:Pt:Finger.third.left:Doc:XR
C1525827|Views:Finding:Point in time:Finger.third.left:Document:XR
C1525947|Pelvis X-ray lateral
C1525947|Pelvis XR Lat
C1525947|View lateral:Finding:Point in time:Pelvis:Document:XR
C1525947|View lateral:Find:Pt:Pelvis:Doc:XR
C1525968|Sacrum XR 2V
C1525968|Sacrum X-ray 2 views
C1525968|Views 2:Finding:Point in time:Sacrum:Document:XR
C1525968|Views 2:Find:Pt:Sacrum:Doc:XR
C1526024|Radius+Ulna-R XR AP+Lat
C1526024|Radius - right and Ulna - right X-ray AP and lateral
C1526024|Views AP & lateral:Find:Pt:Radius.right+Ulna.right:Doc:XR
C1526024|Views AP & lateral:Finding:Point in time:Radius.right+Ulna.right:Document:XR
C1526048|Hip-R XR Judet
C1526048|Hip - right X-ray Judet
C1526048|View Judet:Find:Pt:Hip.right:Doc:XR
C1526048|View Judet:Finding:Point in time:Hip.right:Document:XR
C1526058|Knee-R XR 3V
C1526058|Knee - right X-ray 3 views
C1526058|Views 3:Find:Pt:Knee.right:Doc:XR
C1526058|Views 3:Finding:Point in time:Knee.right:Document:XR
C1526071|Knee - right X-ray PA standing
C1526071|Knee-R XR PA V1 stand
C1526071|View PA^standing:Find:Pt:Knee.right:Doc:XR
C1526071|View PA^standing:Finding:Point in time:Knee.right:Document:XR
C1526102|Should-R XR AP+Stryker Notch
C1526102|Shoulder - right X-ray AP and Stryker Notch
C1526102|Views AP & Stryker Notch:Finding:Point in time:Shoulder.right:Document:XR
C1526102|Views AP & Stryker Notch:Find:Pt:Shoulder.right:Doc:XR
C1526191|T-spine XRTomo
C1526191|Multisection:Finding:Point in time:Spine.thoracic:Document:XR.tomo
C1526191|Multisection:Find:Pt:Spine.thoracic:Doc:XR.tomo
C1526191|Thoracic spine X-ray tomograph
C1526201|Chest US Needle local guid
C1526201|US Guidance for needle localization of Chest
C1526201|Guidance for needle localization:Find:Pt:Chest:Doc:US
C1526201|Guidance for needle localization:Finding:Point in time:Chest:Document:Ultrasound
C1526312|Spine.cavity Flr W contr
C1526312|Spine.cavity Fluoroscopy W contrast
C1526312|Views^W contrast:Find:Pt:Spine.cavity:Doc:XR.fluor
C1526312|Views^W contrast:Finding:Point in time:Spine.cavity:Document:XR.fluor
C1524486|Multisection^W contrast Intravenous:Finding:Point in time:Chest+Abdomen>Aorta:Document:Computerized Tomography
C1524486|Multisection^W contrast IV:Find:Pt:Chest+Abdomen>Aorta:Doc:CT
C1524486|Chest and Abdomen Aorta CT W contrast IV
C1524486|Chest+Abd Aorta CT W contr IV
C1524490|Carotid artery CT angiogram W contrast IV
C1524490|Multisection^W contrast IV:Find:Pt:Head+Neck>Carotid artery:Doc:CT.angio
C1524490|Multisection^W contrast Intravenous:Finding:Point in time:Head+Neck>Carotid artery:Document:Computerized Tomography.angio
C1524490|Carot art CT.Angio W contr IV
C1524502|Elbow MRI W contr IV
C1524502|Elbow MRI W contrast IV
C1524502|Multisection^W contrast Intravenous:Finding:Point in time:Elbow:Document:MRI
C1524502|Multisection^W contrast IV:Find:Pt:Elbow:Doc:MRI
C1524862|Hand CT WO contrast
C1524862|Hand CT WO contr
C1524862|Multisection^WO contrast:Find:Pt:Hand:Doc:CT
C1524862|Multisection^WO contrast:Finding:Point in time:Hand:Document:Computerized Tomography
C1524887|Sacroiliac Joint MRI WO contrast
C1524887|SIJ MRI WO contr
C1524887|Multisection^WO contrast:Find:Pt:Sacroiliac joint:Doc:MRI
C1524887|Multisection^WO contrast:Finding:Point in time:Sacroiliac joint:Document:MRI
C1524519|Thigh-L MRI W contr IV
C1524519|Thigh - left MRI W contrast IV
C1524519|Multisection^W contrast Intravenous:Finding:Point in time:Thigh.left:Document:MRI
C1524519|Multisection^W contrast IV:Find:Pt:Thigh.left:Doc:MRI
C1524523|Ft MRI W contr IV
C1524523|Foot MRI W contrast IV
C1524523|Multisection^W contrast IV:Find:Pt:Foot:Doc:MRI
C1524523|Multisection^W contrast Intravenous:Finding:Point in time:Foot:Document:MRI
C1524913|Lower leg CT WO contrast
C1524913|Lower leg CT WO contr
C1524913|Multisection^WO contrast:Find:Pt:Lower leg:Doc:CT
C1524913|Multisection^WO contrast:Finding:Point in time:Lower leg:Document:Computerized Tomography
C1524564|Larynx MRI W contr IV
C1524564|Larynx MRI W contrast IV
C1524564|Multisection^W contrast Intravenous:Finding:Point in time:Larynx:Document:MRI
C1524564|Multisection^W contrast IV:Find:Pt:Larynx:Doc:MRI
C1524567|Nasoph MRI W contr IV
C1524567|Nasopharynx MRI W contrast IV
C1524567|Multisection^W contrast IV:Find:Pt:Nasopharynx:Doc:MRI
C1524567|Multisection^W contrast Intravenous:Finding:Point in time:Nasopharynx:Document:MRI
C1524198|Should-Bl XR 1V
C1524198|Shoulder - bilateral X-ray Single view
C1524198|View 1:Find:Pt:Shoulder.bilateral:Doc:XR
C1524198|View 1:Finding:Point in time:Shoulder.bilateral:Document:XR
C1524213|Acromioclavicular joint - left X-ray AP single view
C1524213|AC joint-L XR AP 1V
C1524213|View AP:Finding:Point in time:Acromioclavicular joint.left:Document:XR
C1524213|View AP:Find:Pt:Acromioclavicular joint.left:Doc:XR
C1524598|Uterus CT W contr IV
C1524598|Uterus CT W contrast IV
C1524598|Multisection^W contrast Intravenous:Finding:Point in time:Uterus:Document:Computerized Tomography
C1524598|Multisection^W contrast IV:Find:Pt:Uterus:Doc:CT
C1524132|Chest+Abd MRI WO+W contr IV
C1524132|Chest and Abdomen MRI WO and W contrast IV
C1524132|Multisection^WO & W contrast IV:Find:Pt:Chest+Abdomen:Doc:MRI
C1524132|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest+Abdomen:Document:MRI
C1524650|Femur - left X-ray 4 views
C1524650|Femur-L XR 4V
C1524650|Views 4:Find:Pt:Femur.left:Doc:XR
C1524650|Views 4:Finding:Point in time:Femur.left:Document:XR
C1524663|Upper extremity - right MRI WO and W contrast IV
C1524663|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.right:Document:MRI
C1524663|UE-R MRI WO+W contr IV
C1524663|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.right:Doc:MRI
C1524664|Multisection^WO & W contrast IV:Find:Pt:Femur:Doc:CT
C1524664|Multisection^WO & W contrast Intravenous:Finding:Point in time:Femur:Document:Computerized Tomography
C1524664|Femur CT WO and W contrast IV
C1524664|Femur CT WO+W contr IV
C1524994|Clavicle-L XR 2V
C1524994|Clavicle - left X-ray 2 views
C1524994|Views 2:Finding:Point in time:Clavicle.left:Document:XR
C1524994|Views 2:Find:Pt:Clavicle.left:Doc:XR
C1524156|Radius+Ulna XR 2V
C1524156|Radius and Ulna X-ray 2 views
C1524156|Views 2:Find:Pt:Radius+Ulna:Doc:XR
C1524156|Views 2:Finding:Point in time:Radius+Ulna:Document:XR
C1525007|Shoulder - left X-ray 2 views
C1525007|Should-L XR 2V
C1525007|Views 2:Find:Pt:Shoulder.left:Doc:XR
C1525007|Views 2:Finding:Point in time:Shoulder.left:Document:XR
C1524382|Femur-L XRTomo
C1524382|Femur - left X-ray tomograph
C1524382|Multisection:Find:Pt:Femur.left:Doc:XR.tomo
C1524382|Multisection:Finding:Point in time:Femur.left:Document:XR.tomo
C1525039|Radius+Ulna-L XR AP+Lat
C1525039|Radius - left and Ulna.left X-ray AP and lateral
C1525039|Views AP & lateral:Finding:Point in time:Radius.left+Ulna.left:Document:XR
C1525039|Views AP & lateral:Find:Pt:Radius.left+Ulna.left:Doc:XR
C1524784|Spine CT WO and W contrast IV
C1524784|Multisection^WO & W contrast IV:Find:Pt:Spine:Doc:CT
C1524784|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine:Document:Computerized Tomography
C1524784|Spine CT WO+W contr IV
C1524675|Face XR Ltd
C1524675|Facial bones X-ray limited
C1524675|Views limited:Find:Pt:Facial bones:Doc:XR
C1524675|Views limited:Finding:Point in time:Facial bones:Document:XR
C1524676|Mandible XR Ltd
C1524676|Mandible X-ray limited
C1524676|Views limited:Find:Pt:Mandible:Doc:XR
C1524676|Views limited:Finding:Point in time:Mandible:Document:XR
C1525077|Tib+Fib-L XR Obl
C1525077|Tibia - left and Fibula - left X-ray oblique
C1525077|Views oblique:Find:Pt:Tibia.left+Fibula.left:Doc:XR
C1525077|Views oblique:Finding:Point in time:Tibia.left+Fibula.left:Document:XR
C1525094|Coronary aa XRA Atherect W contr IA
C1525094|Coronary arteries Fluoroscopic angiogram Atherectomy W contrast IA
C1525094|Atherectomy^W contrast IA:Find:Pt:Coronary arteries:Doc:XR.fluor.angio
C1525094|Atherectomy^W contrast Intra-arterial:Finding:Point in time:Coronary arteries:Document:XR.fluor.angio
C1830189|Prostate US Bx needle guid
C1830189|US Guidance for needle biopsy of Prostate
C1830189|Guidance for biopsy.needle:Find:Pt:Prostate:Doc:US
C1830189|Guidance for biopsy.needle:Finding:Point in time:Prostate:Document:Ultrasound
C1830263|Foot vessels US.doppler
C1830263|Ft ves DOP
C1830263|Multisection:Find:Pt:Foot vessels:Doc:US.doppler
C1830263|Multisection:Finding:Point in time:Foot vessels:Document:Ultrasound.doppler
C1830071|Chest XR GE 4 & PA+Lat
C1830071|Chest X-ray GE 4 and Pa and Lateral views
C1830071|Views GE 4 & PA & lateral:Find:Pt:Chest:Doc:XR
C1830071|Views GE 4 & PA & lateral:Finding:Point in time:Chest:Document:XR
C1715377|Muscle CT FNA Asp
C1715377|CT Guidance for fine needle aspiration of Muscle
C1715377|Guidance for aspiration.fine needle:Finding:Point in time:Muscle:Document:Computerized Tomography
C1715377|Guidance for aspiration.fine needle:Find:Pt:Muscle:Doc:CT
C1715387|Abd+Pelvis CT
C1715387|Abdomen and Pelvis CT
C1715387|Multisection:Finding:Point in time:Abdomen+Pelvis:Document:Computerized Tomography
C1715387|Multisection:Find:Pt:Abdomen+Pelvis:Doc:CT
C1715410|Abd+Pelvis RI for Tumor
C1715410|Abdomen and Pelvis Scan for tumor
C1715410|Views for tumor:Finding:Point in time:Abdomen+Pelvis:Document:Radnuc
C1715410|Views for tumor:Find:Pt:Abdomen+Pelvis:Doc:Radnuc
C1632265|Ribs - bilateral and Chest X-ray and PA chest
C1632265|Views & PA chest:Finding:Point in time:Ribs.bilateral+Chest:Document:XR
C1632265|Views & PA chest:Find:Pt:Ribs.bilateral+Chest:Doc:XR
C1632265|Ribs-Bl+Chest XR +PA Chst
C1634506|L-spine XR AP 1V W L-bending
C1634506|View AP^W L-bending:Find:Pt:Spine.lumbar:Doc:XR
C1634506|View AP^W L-bending:Finding:Point in time:Spine.lumbar:Document:XR
C1634506|Lumbar spine X-ray AP single view W left bending
C1714790|Knee-L MRI Dyn W contr IV
C1714790|Knee - left MRI dynamic W contrast IV
C1714790|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Knee.left:Document:MRI
C1714790|Multisection dynamic^W contrast IV:Find:Pt:Knee.left:Doc:MRI
C1714809|XXX Flr 90M
C1714809|Unspecified body region Fluoroscopy 90 minutes
C1714809|View:Find:90M:XXX:Doc:XR.fluor
C1714809|View:Finding:90 minutes:To be specified in another part of the message:Document:XR.fluor
C1714903|Guidance for drainage of abscess:Finding:Point in time:Subphrenic space:Document:Computerized Tomography
C1714903|Subphrenic Space CT Abscess drain guid
C1714903|CT Guidance for drainage of abscess of Subphrenic space
C1714903|Guidance for drainage of abscess:Find:Pt:Subphrenic space:Doc:CT
C1714928|Orbit+Face XR
C1714928|Views:Find:Pt:Orbit+Facial bones:Doc:XR
C1714928|Views:Finding:Point in time:Orbit+Facial bones:Document:XR
C1714928|Orbit and Facial bones X-ray
C1714957|Hand X-ray portable
C1714957|Hand XR port
C1714957|Views portable:Find:Pt:Hand:Doc:XR
C1714957|Views portable:Finding:Point in time:Hand:Document:XR
C1715026|Liver RI Flow W Tc99mRBC IV
C1715026|Liver Scan flow W Tc-99m tagged RBC IV
C1715026|Views flow^W Tc-99m tagged RBC IV:Find:Pt:Liver:Doc:Radnuc
C1715026|Views flow^W Tc-99m tagged RBC Intravenous:Finding:Point in time:Liver:Document:Radnuc
C1630190|T+L-spine XR Scoli AP 1V Stand+In Brace
C1630190|View scoliosis AP^standing & in brace:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1630190|Spine Thoracic and Lumbar X-ray scoliosis AP standing and in brace
C1630190|View scoliosis AP^standing & in brace:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1644662|Spleen Scan flow
C1644662|Spleen RI Flow W RNC IV
C1644662|Views flow^W radionuclide Intravenous:Finding:Point in time:Spleen:Document:Radnuc
C1644662|Views flow^W radionuclide IV:Find:Pt:Spleen:Doc:Radnuc
C1632388|Guidance for superficial biopsy:Finding:Point in time:Bone:Document:Computerized Tomography
C1632388|Bone CT Bx super guid
C1632388|Guidance for superficial biopsy:Find:Pt:Bone:Doc:CT
C1632388|CT Guidance for superficial biopsy of Bone
C1646329|Pelvis X-ray Single view portable
C1646329|Pelvis XR 1V port
C1646329|View 1 portable:Finding:Point in time:Pelvis:Document:XR
C1646329|View 1 portable:Find:Pt:Pelvis:Doc:XR
C1633446|Brst-R Mam Localization guid
C1633446|Mammogram Guidance for localization of Breast - right
C1633446|Guidance for localization:Find:Pt:Breast.right:Doc:Mam
C1633446|Guidance for localization:Finding:Point in time:Breast.right:Document:Mam
C1954364|Mammogram Guidance for sentinel lymph node injection of Breast - left
C1954364|Brst-L Mam Sentinel LN inj guid
C1954364|Guidance for sentinel lymph node injection:Finding:Point in time:Breast.left:Document:Mam
C1954364|Guidance for sentinel lymph node injection:Find:Pt:Breast.left:Doc:Mam
C1954368|Mammogram Guidance for sentinel lymph node injection of Breast - right
C1954368|Brst-R Mam Sentinel LN inj guid
C1954368|Guidance for sentinel lymph node injection:Finding:Point in time:Breast.right:Document:Mam
C1954368|Guidance for sentinel lymph node injection:Find:Pt:Breast.right:Doc:Mam
C1954371|Scrotum+Test DOP
C1954371|Scrotum and Testicle US.doppler
C1954371|Multisection:Find:Pt:Scrotum+Testicle:Doc:US.doppler
C1954371|Multisection:Finding:Point in time:Scrotum+Testicle:Document:Ultrasound.doppler
C1954372|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Retroperitoneum:Document:Computerized Tomography
C1954372|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Retroperitoneum:Doc:CT
C1954372|Retroperitoneum CT WO and W contrast IV
C1954372|Retroperitoneum CT WO+W contr IV
C1953326|Spine CT W contrast IT
C1953326|Spine CT W contr IT
C1953326|Multisection^W contrast IT:Find:Pt:Spine:Doc:CT
C1953326|Multisection^W contrast Intrathecal:Finding:Point in time:Spine:Document:Computerized Tomography
C1953943|Deprecated Temporal bones MRI W contr IV
C1953943|Deprecated Temporal bones MRI W contrast IV
C1953943|Multisection^W contrast Intravenous:Finding:Point in time:Temporal bones:Narrative:MRI
C1953943|Multisection^W contrast IV:Find:Pt:Temporal bone:Nar:MRI
C1953943|Multisection^W contrast Intravenous:Finding:Point in time:Temporal bone:Narrative:MRI
C1953952|Nasoph CT W contr IV
C1953952|Nasopharynx CT W contrast IV
C1953952|Multisection^W contrast IV:Find:Pt:Nasopharynx:Doc:CT
C1953952|Multisection^W contrast Intravenous:Finding:Point in time:Nasopharynx:Document:Computerized Tomography
C1953959|Brain.temporal MRI WO contrast
C1953959|Brain.temporal MRI WO contr
C1953959|Multisection^WO contrast:Finding:Point in time:Brain.temporal:Document:MRI
C1953959|Multisection^WO contrast:Find:Pt:Brain.temporal:Doc:MRI
C1953960|Multisection^WO & W contrast IV:Find:Pt:Clavicle.right:Doc:MRI
C1953960|Clavicle - right MRI WO and W contrast IV
C1953960|Clavicle-R MRI WO+W contr IV
C1953960|Multisection^WO & W contrast Intravenous:Finding:Point in time:Clavicle.right:Document:MRI
C3533571|Multisection^W contrast IV & W air contrast PR:Find:Pt:Abdomen+Pelvis>Colon+Rectum:Doc:CT
C3533571|Multisection^W contrast Intravenous & W air contrast Rectal:Finding:Point in time:Abdomen+Pelvis>Colon+Rectum:Document:Computerized Tomography
C3533571|Colon and Rectum CT W contrast IV and W air contrast PR
C3533571|Colon+Rectum CT W contr IV+Air contr PR
C3262939|Sacrum and Coccyx CT
C3262939|Sacrum+Coccyx CT
C3262939|Multisection:Find:Pt:Sacrum+Coccyx:Doc:CT
C3262939|Multisection:Finding:Point in time:Sacrum+Coccyx:Document:Computerized Tomography
C3262962|Knee-L XR 2V+Sunrise
C3262962|Knee - left X-ray 2 views and Sunrise
C3262962|Views 2 & Sunrise:Finding:Point in time:Knee.left:Document:XR
C3262962|Views 2 & Sunrise:Find:Pt:Knee.left:Doc:XR
C3263009|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast implant:Document:MRI
C3263009|Breast implant MRI WO and W contrast IV
C3263009|Brst implant MRI WO+W contr IV
C3263009|Multisection^WO & W contrast IV:Find:Pt:Breast implant:Doc:MRI
C3482440|T-spine Flr PC Vertebroplasty guid
C3482440|Guidance for percutaneous vertebroplasty:Finding:Point in time:Spine.thoracic:Document:XR.fluor
C3482440|Guidance for percutaneous vertebroplasty:Find:Pt:Spine.thoracic:Doc:XR.fluor
C3482440|Fluoroscopy Guidance for percutaneous vertebroplasty of Thoracic spine
C3482446|T-spine CT W contr ID
C3482446|Multisection^W contrast intradisc:Find:Pt:Spine.thoracic:Doc:CT
C3482446|Multisection^W contrast intradisc:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C3482446|Thoracic spine CT W contrast intradisc
C3262469|MRI Guidance for biopsy of Breast - left
C3262469|Brst-L MRI Bx guid
C3262469|Guidance for biopsy:Finding:Point in time:Breast.left:Document:MRI
C3262469|Guidance for biopsy:Find:Pt:Breast.left:Doc:MRI
C3263220|Spinal cord US Bx needle guid
C3263220|US Guidance for needle biopsy of Spinal cord
C3263220|Guidance for biopsy.needle:Finding:Point in time:Spinal cord:Document:Ultrasound
C3263220|Guidance for biopsy.needle:Find:Pt:Spinal cord:Doc:US
C3262923|Salivary gland CT Bx needle guid
C3262923|CT Guidance for needle biopsy of Salivary gland
C3262923|Guidance for biopsy.needle:Finding:Point in time:Salivary gland:Document:Computerized Tomography
C3262923|Guidance for biopsy.needle:Find:Pt:Salivary gland:Doc:CT
C0944171|Views:Finding:Point in time:Hand:Narrative:XR
C0944171|Hand XR
C0944171|Hand X-ray
C0944171|Views:Find:Pt:Hand:Doc:XR
C0944171|Views:Finding:Point in time:Hand:Document:XR
C0942178|Toes-R XR
C0942178|Toes - right X-ray
C0942178|Views:Find:Pt:Toes.right:Doc:XR
C0942178|Views:Finding:Point in time:Toes.right:Document:XR
C0942213|Ankle-L MRI
C0942213|Ankle - left MRI
C0942213|Multisection:Finding:Point in time:Ankle.left:Document:MRI
C0942213|Multisection:Find:Pt:Ankle.left:Doc:MRI
C0942254|Pelvis+Hip-Bl MRI
C0942254|Pelvis and Hip - bilateral MRI
C0942254|Multisection:Find:Pt:Pelvis+Hip.bilateral:Doc:MRI
C0942254|Multisection:Finding:Point in time:Pelvis+Hip.bilateral:Document:MRI
C0942271|Wrist - bilateral MRI
C0942271|Wrist-Bl MRI
C0942271|Multisection:Finding:Point in time:Wrist.bilateral:Document:MRI
C0942271|Multisection:Find:Pt:Wrist.bilateral:Doc:MRI
C0942344|Knee-Bl XR AP+Lat stand
C0942344|Knee - bilateral X-ray AP and lateral standing
C0942344|Views AP & lateral^standing:Finding:Point in time:Knee.bilateral:Document:XR
C0942344|Views AP & lateral^standing:Find:Pt:Knee.bilateral:Doc:XR
C0945349|Hip - left X-ray Single view
C0945349|Hip-L XR 1V
C0945349|View 1:Finding:Point in time:Hip.left:Document:XR
C0945349|View 1:Find:Pt:Hip.left:Doc:XR
C0884112|CT Guidance for biopsy of Lung
C0884112|Lung CT Bx guid
C0884112|Guidance for biopsy:Find:Pt:Chest>Lung:Doc:CT
C0884112|Guidance for biopsy:Finding:Point in time:Chest>Lung:Document:Computerized Tomography
C0882078|Views:Finding:Point in time:Radius+Ulna:Narrative:XR
C0882078|Radius+Ulna XR
C0882078|Radius and Ulna X-ray
C0882078|Views:Find:Pt:Radius+Ulna:Doc:XR
C0882078|Views:Finding:Point in time:Radius+Ulna:Document:XR
C0942117|Ankle-Bl XR
C0942117|Ankle - bilateral X-ray
C0942117|Views:Finding:Point in time:Ankle.bilateral:Document:XR
C0942117|Views:Find:Pt:Ankle.bilateral:Doc:XR
C0881783|Aorta XRA Angpsty W contr IA
C0881783|Aorta Fluoroscopic angiogram Angioplasty W contrast IA
C0881783|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Aorta:Document:XR.fluor.angio
C0881783|Angioplasty^W contrast IA:Find:Pt:Aorta:Doc:XR.fluor.angio
C0881800|Abdomen X-ray AP left lateral-decubitus
C0881800|Abd XR AP L-Lat Decub
C0881800|View AP L-lateral-decubitus:Find:Pt:Abdomen:Doc:XR
C0881800|View AP L-lateral-decubitus:Finding:Point in time:Abdomen:Document:XR
C0881839|Brst Mam Dx Ltd
C0881839|Breast Mammogram diagnostic limited
C0881839|Views diagnostic limited:Finding:Point in time:Breast:Document:Mam
C0881839|Views diagnostic limited:Find:Pt:Breast:Doc:Mam
C0881879|Chest XR AP+AP R-Lat Debub
C0881879|Chest X-ray AP and AP right lateral-decubitus
C0881879|Views AP & AP R-lateral-decubitus:Find:Pt:Chest:Doc:XR
C0881879|Views AP & AP R-lateral-decubitus:Finding:Point in time:Chest:Document:XR
C0881967|Views:Finding:Point in time:Hip:Narrative:XR
C0881967|Hip X-ray
C0881967|Hip XR
C0881967|Views:Find:Pt:Hip:Doc:XR
C0881967|Views:Finding:Point in time:Hip:Document:XR
C0881987|Kidney - bilateral X-ray tomograph WO contrast and 10M post contrast IV
C0881987|Multisection^WO contrast & 10M post contrast IV:Find:Pt:Kidney.bilateral:Doc:XR.tomo
C0881987|Multisection^WO contrast & 10 minutes post contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:XR.tomo
C0881987|Kdny-Bl XRTomo WO contr+10m p contr IV
C0881993|Abd XR AP+Lat port
C0881993|Abdomen X-ray AP and lateral portable
C0881993|Views AP & lateral portable:Finding:Point in time:Abdomen:Document:XR
C0881993|Views AP & lateral portable:Find:Pt:Abdomen:Doc:XR
C1114508|Upper arm MRI WO contr
C1114508|Upper arm MRI WO contrast
C1114508|Multisection^WO contrast:Finding:Point in time:Upper arm:Document:MRI
C1114508|Multisection^WO contrast:Find:Pt:Upper arm:Doc:MRI
C1114532|Deprecated Sinuses XR.Tomo PA+Lat
C1114532|Views PA & lateral:Find:Pt:Sinuses:Nar:XR.tomo
C1114532|Deprecated Views PA & lateral
C1114532|Views PA & lateral:Finding:Point in time:Sinuses:Narrative:XR.tomo
C2713289|View 1 portable:Finding:Point in time:Spine.cervical:Narrative:XR
C2713289|C-spine XR 1V port
C2713289|View 1 portable:Find:Pt:Spine.cervical:Doc:XR
C2713289|View 1 portable:Finding:Point in time:Spine.cervical:Document:XR
C2713289|Cervical spine X-ray Single view portable
C1114569|Multisection 3 views^W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:XR.tomo
C1114569|Multisection 3 views^W contrast IV:Find:Pt:Kidney.bilateral:Doc:XR.tomo
C1114569|Kidney - bilateral X-ray tomograph 3 views W contrast IV
C1114569|Kdny-Bl XRTomo 3V W contr IV
C1114576|Pelvis+Hip XR AP+Lat Frog
C1114576|Pelvis and Hip X-ray AP and lateral frog
C1114576|Views AP & lateral frog:Find:Pt:Pelvis+Hip:Doc:XR
C1114576|Views AP & lateral frog:Finding:Point in time:Pelvis+Hip:Document:XR
C1114581|L-spine XR 3V port
C1114581|Views 3 portable:Finding:Point in time:Spine.lumbar:Document:XR
C1114581|Views 3 portable:Find:Pt:Spine.lumbar:Doc:XR
C1114581|Lumbar spine X-ray 3 views portable
C1114611|UGI+SB Flr W contr PO
C1114611|Upper Gastrointestine and Small bowel Fluoroscopy W contrast PO
C1114611|View^W contrast Oral:Finding:Point in time:Gastrointestine.upper+Small bowel:Document:XR.fluor
C1114611|View^W contrast PO:Find:Pt:Gastrointestine.upper+Small bowel:Doc:XR.fluor
C1114682|Renal ves MRI.Angio W contr IV
C1114682|Renal vessels MRI angiogram W contrast IV
C1114682|Multisection^W contrast Intravenous:Finding:Point in time:Renal vessels:Document:MRI.angio
C1114682|Multisection^W contrast IV:Find:Pt:Renal vessels:Doc:MRI.angio
C1114416|Nasopharynx+Neck CT WO contr
C1114416|Nasopharynx and Neck CT WO contrast
C1114416|Multisection^WO contrast:Finding:Point in time:Nasopharynx+Neck:Document:Computerized Tomography
C1114416|Multisection^WO contrast:Find:Pt:Nasopharynx+Neck:Doc:CT
C1114428|Multisection^W contrast:Find:Pt:Abdomen:Doc:CT
C1114428|Deprecated Abd CT W contr
C1114428|Deprecated Abdomen CT W contrast
C1114428|Multisection^W contrast:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1114449|Spleen CT WO contrast
C1114449|Spleen CT WO contr
C1114449|Multisection^WO contrast:Finding:Point in time:Abdomen>Spleen:Document:Computerized Tomography
C1114449|Multisection^WO contrast:Find:Pt:Abdomen>Spleen:Doc:CT
C1114931|BDs+GB Flr W contr via T-tb
C1114931|Biliary ducts and Gallbladder Fluoroscopy W contrast via T-tube
C1114931|Views^W contrast via T-tube:Find:Pt:Biliary ducts+Gallbladder:Doc:XR.fluor
C1114931|Views^W contrast via T-tube:Finding:Point in time:Biliary ducts+Gallbladder:Document:XR.fluor
C1543447|Fistula Flr W contr retro
C1543447|Fistula Fluoroscopy W contrast retrograde
C1543447|Views^W contrast retrograde:Find:Pt:Fistula:Doc:XR.fluor
C1543447|Views^W contrast retrograde:Finding:Point in time:Fistula:Document:XR.fluor
C1543742|GI RI W Tc99mSC IV
C1543742|Gastrointestine Scan W Tc-99m SC IV
C1543742|Views^W Tc-99m SC IV:Find:Pt:Gastrointestine:Doc:Radnuc
C1543742|Views^W Tc-99m Subcutaneous Intravenous:Finding:Point in time:Gastrointestine:Document:Radnuc
C1543874|Liver Scan static
C1543874|Liver RI Static W RNC IV
C1543874|Views static^W radionuclide IV:Find:Pt:Liver:Doc:Radnuc
C1543874|Views static^W radionuclide Intravenous:Finding:Point in time:Liver:Document:Radnuc
C1542901|SPECT W I-131 mIBG IV
C1542901|Multisection^W I-131 MIBG IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1542901|Multisection^W I-131 MIBG Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543901|Bone SPECT
C1543901|Multisection^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1543901|Multisection^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1543901|Bone SPECT W RNC IV
C1543938|Heart SPECT gated
C1543938|Hrt SPECT Gated W RNC IV
C1543938|Multisection gated^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543938|Multisection gated^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543948|Deprecated View gated^W stress & W radionuclide IV:Find:Pt:Heart:Nar:Radnuc
C1543948|View gated^W stress & W radionuclide IV:Find:Pt:Heart:Nar:Radnuc
C1543948|Deprecated Hrt RI Gated V1 W Stress+W RN
C1543948|Deprecated Heart Scintigraphy gated W stress & W radionuclide IV
C1543948|View gated^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1542853|Hrt RI WM+EF W RNC IV
C1542853|Heart Scan wall motion and ejection fraction
C1542853|Views wall motion & ejection fraction^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1542853|Views wall motion & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543528|US Guidance for aspiration of Ovary
C1543528|Ovary US Asp guid
C1543528|Guidance for aspiration:Find:Pt:Ovary:Doc:US
C1543528|Guidance for aspiration:Finding:Point in time:Ovary:Document:Ultrasound
C1543153|Kidney transplant US
C1543153|Multisection:Finding:Point in time:Kidney transplant:Document:Ultrasound
C1543153|Multisection:Find:Pt:Kidney transplant:Doc:US
C1543577|Upper extremity vein - left US.doppler
C1543577|UE v-L DOP
C1543577|Multisection:Find:Pt:Upper extremity vein.left:Doc:US.doppler
C1543577|Multisection:Finding:Point in time:Upper extremity vein.left:Document:Ultrasound.doppler
C1543602|Unspecified body region US of foreign body
C1543602|XXX US of FB
C1543602|Multisection of foreign body:Find:Pt:XXX:Doc:US
C1543602|Multisection of foreign body:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1543217|Hep vs XRA W contr IV+Hemodynamics
C1543217|Hepatic veins Fluoroscopic angiogram W contrast IV and W hemodynamics
C1543217|Views^W contrast IV & W hemodynamics:Find:Pt:Hepatic veins:Doc:XR.fluor.angio
C1543217|Views^W contrast Intravenous & W hemodynamics:Finding:Point in time:Hepatic veins:Document:XR.fluor.angio
C1525168|Hip-R XR True Lat
C1525168|Hip - right X-ray true lateral
C1525168|View true lateral:Find:Pt:Hip.right:Doc:XR
C1525168|View true lateral:Finding:Point in time:Hip.right:Document:XR
C1525170|Orbit - right X-ray
C1525170|Orbit-R XR
C1525170|Views:Finding:Point in time:Orbit.right:Document:XR
C1525170|Views:Find:Pt:Orbit.right:Doc:XR
C1525932|Shoulder - right X-ray transthoracic
C1525932|Should-R XR Transthoracic
C1525932|View transthoracic:Finding:Point in time:Shoulder.right:Document:XR
C1525932|View transthoracic:Find:Pt:Shoulder.right:Doc:XR
C1526758|Multisection^WO & W contrast IV:Find:Pt:Wrist.right:Doc:CT
C1526758|Wrist - right CT WO and W contrast IV
C1526758|Multisection^WO & W contrast Intravenous:Finding:Point in time:Wrist.right:Document:Computerized Tomography
C1526758|Wrist-R CT WO+W contr IV
C1526768|Extremity lymphatics - right Fluoroscopy W contrast intra lymphatic
C1526768|Extr lymph-R Flr W contr IL
C1526768|Views^W contrast intra lymphatic:Find:Pt:Extremity lymphatics.right:Doc:XR.fluor
C1526768|Views^W contrast intra lymphatic:Finding:Point in time:Extremity lymphatics.right:Document:XR.fluor
C1542973|SPECT for Tumor W Ga-67 IV
C1542973|Multisection for tumor^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1542973|Multisection for tumor^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1526787|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.left:Doc:MRI
C1526787|Upper extremity - left MRI WO and W contrast IV
C1526787|UE-L MRI WO+W contr IV
C1526787|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.left:Document:MRI
C1526794|Wrist-L XR Ltd
C1526794|Wrist - left X-ray limited
C1526794|Views limited:Finding:Point in time:Wrist.left:Document:XR
C1526794|Views limited:Find:Pt:Wrist.left:Doc:XR
C1525186|Multisection^W contrast IS:Find:Pt:Upper joint:Doc:CT
C1525186|Deprecated Upper joint CT W contr IS
C1525186|Multisection^W contrast Intrasynovial:Finding:Point in time:Upper joint:Document:Computerized Tomography
C1525186|Deprecated Upper Joint CT W contrast IS
C1524238|C-spine CT Ltd WO contr
C1524238|Multisection limited^WO contrast:Find:Pt:Spine.cervical:Doc:CT
C1524238|Multisection limited^WO contrast:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C1524238|Cervical spine CT limited WO contrast
C1525307|View Harris:Find:Pt:Calcaneus.bilateral:Doc:XR
C1525307|View Harris:Finding:Point in time:Calcaneus.bilateral:Document:XR
C1525307|Deprecated Calcaneus - bilateral X-ray Harris
C1525307|Deprecated Heel-Bl XR Harris
C1525310|Knee XR Holmblad
C1525310|Knee X-ray Holmblad
C1525310|View Holmblad:Finding:Point in time:Knee:Document:XR
C1525310|View Holmblad:Find:Pt:Knee:Doc:XR
C1525325|Hip - bilateral X-ray lateral frog
C1525325|Hip-Bl XR Lat Frog
C1525325|View lateral frog:Finding:Point in time:Hip.bilateral:Document:XR
C1525325|View lateral frog:Find:Pt:Hip.bilateral:Doc:XR
C1525215|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.joint.left:Document:MRI
C1525215|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.joint.left:Doc:MRI
C1525215|Upper extremity joint - left MRI WO and W contrast IV
C1525215|UE joint-L MRI WO+W contr IV
C1525235|UE ves-R MRI.Angio WO+W contr IV
C1525235|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity vessels.right:Document:MRI.angio
C1525235|Multisection^WO & W contrast IV:Find:Pt:Upper extremity vessels.right:Doc:MRI.angio
C1525235|Upper extremity vessels - right MRI angiogram WO and W contrast IV
C1525242|Temporal bone-R CT WO contr
C1525242|Temporal bone - right CT WO contrast
C1525242|Multisection^WO contrast:Find:Pt:Temporal bone.right:Doc:CT
C1525242|Multisection^WO contrast:Finding:Point in time:Temporal bone.right:Document:Computerized Tomography
C1525262|Maxillofacial CT Bx guid
C1525262|CT Guidance for biopsy of Maxillofacial region
C1525262|Guidance for biopsy:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1525262|Guidance for biopsy:Find:Pt:Head>Maxillofacial region:Doc:CT
C1524687|Knee-L XR Rosenberg stand
C1524687|Knee - left X-ray Rosenberg standing
C1524687|View Rosenberg^standing:Finding:Point in time:Knee.left:Document:XR
C1524687|View Rosenberg^standing:Find:Pt:Knee.left:Doc:XR
C1525350|Breast Mammogram tangential
C1525350|Brst Mam Tangential
C1525350|View tangential:Finding:Point in time:Breast:Document:Mam
C1525350|View tangential:Find:Pt:Breast:Doc:Mam
C1525551|Should-Bl XR Outlet+Y
C1525551|Shoulder - bilateral X-ray outlet and Y
C1525551|Views outlet & Y:Find:Pt:Shoulder.bilateral:Doc:XR
C1525551|Views outlet & Y:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525565|Face XR Lat+Caldwell+Waters+SMV+Towne
C1525565|Facial bones X-ray lateral and Caldwell and Waters and submentovertex and Towne
C1525565|Views lateral & Caldwell & Waters & submentovertex & Towne:Find:Pt:Facial bones:Doc:XR
C1525565|Views lateral & Caldwell & Waters & submentovertex & Towne:Finding:Point in time:Facial bones:Document:XR
C1525588|Joint Fluoroscopy W contrast IS
C1525588|Views^W contrast Intrasynovial:Finding:Point in time:Joint:Document:XR.fluor
C1525588|Joint Flr W contr IS
C1525588|Views^W contrast IS:Find:Pt:Joint:Doc:XR.fluor
C1525598|Ankle - bilateral X-ray standing
C1525598|Ankle-Bl XR stand
C1525598|Views^standing:Finding:Point in time:Ankle.bilateral:Document:XR
C1525598|Views^standing:Find:Pt:Ankle.bilateral:Doc:XR
C1525620|Sternoclavicular Joint CT
C1525620|SC joint CT
C1525620|Multisection:Find:Pt:Sternoclavicular joint:Doc:CT
C1525620|Multisection:Finding:Point in time:Sternoclavicular joint:Document:Computerized Tomography
C1525638|TMJ MRI W contr IV
C1525638|Temporomandibular joint MRI W contrast IV
C1525638|Multisection^W contrast Intravenous:Finding:Point in time:Temporomandibular joint:Document:MRI
C1525638|Multisection^W contrast IV:Find:Pt:Temporomandibular joint:Doc:MRI
C1525641|TMJ-L MRI W contr IV
C1525641|Temporomandibular joint - left MRI W contrast IV
C1525641|Multisection^W contrast IV:Find:Pt:Temporomandibular joint.left:Doc:MRI
C1525641|Multisection^W contrast Intravenous:Finding:Point in time:Temporomandibular joint.left:Document:MRI
C1525701|Deprecated
C1525701|Views runoff^W contrast IA:Find:Pt:Aorta+Femoral artery:Nar:XR.fluor.angio
C1525701|Views runoff^W contrast Intra-arterial:Finding:Point in time:Aorta+Femoral artery:Narrative:XR.fluor.angio
C1525701|Deprecated Aorta and Femoral artery Narrative Fluoroscopic angiogram runoff W contrast IA
C1525709|Ac arch+Subclavian a-L XRA W contr IA
C1525709|Aortic arch and Subclavian artery - left Fluoroscopic angiogram W contrast IA
C1525709|Views^W contrast IA:Find:Pt:Aortic arch+Subclavian artery.left:Doc:XR.fluor.angio
C1525709|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Subclavian artery.left:Document:XR.fluor.angio
C1525714|Brachial artery - bilateral Fluoroscopic angiogram W contrast IA
C1525714|Brach a-Bl XRA W contr IA
C1525714|Views^W contrast IA:Find:Pt:Brachial artery.bilateral:Doc:XR.fluor.angio
C1525714|Views^W contrast Intra-arterial:Finding:Point in time:Brachial artery.bilateral:Document:XR.fluor.angio
C1524694|Wrist MRI W contr IV
C1524694|Wrist MRI W contrast IV
C1524694|Multisection^W contrast IV:Find:Pt:Wrist:Doc:MRI
C1524694|Multisection^W contrast Intravenous:Finding:Point in time:Wrist:Document:MRI
C1525779|Hand - left X-ray Bora
C1525779|Hand-L XR Bora
C1525779|View Bora:Find:Pt:Hand.left:Doc:XR
C1525779|View Bora:Finding:Point in time:Hand.left:Document:XR
C1525847|Breast Mammogram spot
C1525847|Brst Mam Spot
C1525847|Views spot:Finding:Point in time:Breast:Document:Mam
C1525847|Views spot:Find:Pt:Breast:Doc:Mam
C1525809|C-spine ves MRI.Angio WO+W contr IV
C1525809|Multisection^WO & W contrast IV:Find:Pt:Spine.cervical vessels:Doc:MRI.angio
C1525809|Cervical Spine vessels MRI angiogram WO and W contrast IV
C1525809|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.cervical vessels:Document:MRI.angio
C1525815|Thoracic Spine vessels MRI angiogram WO contrast
C1525815|T-spine ves MRI.Angio WO contr
C1525815|Multisection^WO contrast:Finding:Point in time:Spine.thoracic vessels:Document:MRI.angio
C1525815|Multisection^WO contrast:Find:Pt:Spine.thoracic vessels:Doc:MRI.angio
C1525970|Sacrum XRTomo
C1525970|Sacrum X-ray tomograph
C1525970|Multisection:Finding:Point in time:Sacrum:Document:XR.tomo
C1525970|Multisection:Find:Pt:Sacrum:Doc:XR.tomo
C1526010|Finger-R XR 2V
C1526010|Finger - right X-ray 2 views
C1526010|Views 2:Finding:Point in time:Finger.right:Document:XR
C1526010|Views 2:Find:Pt:Finger.right:Doc:XR
C1526029|Hand-R XR PA+Lat
C1526029|Hand - right X-ray PA and lateral
C1526029|Views PA & lateral:Find:Pt:Hand.right:Doc:XR
C1526029|Views PA & lateral:Finding:Point in time:Hand.right:Document:XR
C1526079|Knee-R XR 4V stand
C1526079|Knee - right X-ray 4 views standing
C1526079|Views 4^standing:Find:Pt:Knee.right:Doc:XR
C1526079|Views 4^standing:Finding:Point in time:Knee.right:Document:XR
C1526081|LE ves-R XRA W contr
C1526081|Lower extremity vessels - right Fluoroscopic angiogram W contrast
C1526081|Views^W contrast:Find:Pt:Lower extremity vessels.right:Doc:XR.fluor.angio
C1526081|Views^W contrast:Finding:Point in time:Lower extremity vessels.right:Document:XR.fluor.angio
C1524274|Sternum X-ray tomograph
C1524274|Sternum XRTomo
C1524274|Multisection:Find:Pt:Sternum:Doc:XR.tomo
C1524274|Multisection:Finding:Point in time:Sternum:Document:XR.tomo
C1526173|Tib+Fib XR Lat
C1526173|Tibia and Fibula X-ray lateral
C1526173|View lateral:Find:Pt:Tibia+Fibula:Doc:XR
C1526173|View lateral:Finding:Point in time:Tibia+Fibula:Document:XR
C1524707|Wrist XR Lat W FE
C1524707|Wrist X-ray lateral W flexion and W extension
C1524707|Views lateral^W flexion & W extension:Find:Pt:Wrist:Doc:XR
C1524707|Views lateral^W flexion & W extension:Finding:Point in time:Wrist:Document:XR
C1524708|Wrist X-ray lateral
C1524708|Wrist XR Lat
C1524708|View lateral:Finding:Point in time:Wrist:Document:XR
C1524708|View lateral:Find:Pt:Wrist:Doc:XR
C1524717|Upper extremity - left US
C1524717|UE-L US
C1524717|Multisection:Find:Pt:Upper extremity.left:Doc:US
C1524717|Multisection:Finding:Point in time:Upper extremity.left:Document:Ultrasound
C1526286|Sacrum US
C1526286|Multisection:Find:Pt:Sacrum:Doc:US
C1526286|Multisection:Finding:Point in time:Sacrum:Document:Ultrasound
C1526336|T+L-spine XR AP+Lat
C1526336|Spine Thoracic and Lumbar X-ray AP and lateral
C1526336|Views AP & lateral:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1526336|Views AP & lateral:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1525146|UE a DOP Ltd
C1525146|Upper extremity artery US.doppler limited
C1525146|Multisection limited:Finding:Point in time:Upper extremity artery:Document:Ultrasound.doppler
C1525146|Multisection limited:Find:Pt:Upper extremity artery:Doc:US.doppler
C1508084|Abd XR AP+L-Post Obl
C1508084|Abdomen X-ray AP and left posterior oblique
C1508084|Views AP & L-posterior oblique:Find:Pt:Abdomen:Doc:XR
C1508084|Views AP & L-posterior oblique:Finding:Point in time:Abdomen:Document:XR
C1526318|Bladder+Urethra Flr W contr Ante
C1526318|Urinary Bladder and Urethra Fluoroscopy W contrast antegrade
C1526318|Views^W contrast antegrade:Finding:Point in time:Urinary bladder+Urethra:Document:XR.fluor
C1526318|Views^W contrast antegrade:Find:Pt:Urinary bladder+Urethra:Doc:XR.fluor
C1524471|Multisection^W contrast IS:Find:Pt:Knee.right:Doc:MRI
C1524471|Knee-R MRI W contr IS
C1524471|Knee - right MRI W contrast IS
C1524471|Multisection^W contrast Intrasynovial:Finding:Point in time:Knee.right:Document:MRI
C1524494|Brst-Bl MRI W contr IV
C1524494|Breast - bilateral MRI W contrast IV
C1524494|Multisection^W contrast IV:Find:Pt:Breast.bilateral:Doc:MRI
C1524494|Multisection^W contrast Intravenous:Finding:Point in time:Breast.bilateral:Document:MRI
C1524512|UE-Bl CT W contr IV
C1524512|Upper extremity - bilateral CT W contrast IV
C1524512|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.bilateral:Document:Computerized Tomography
C1524512|Multisection^W contrast IV:Find:Pt:Upper extremity.bilateral:Doc:CT
C1524163|Hrt MRI W contr IV
C1524163|Heart MRI W contrast IV
C1524163|Multisection^W contrast Intravenous:Finding:Point in time:Heart:Document:MRI
C1524163|Multisection^W contrast IV:Find:Pt:Heart:Doc:MRI
C1524568|Neck ves CT.Angio W contr IV
C1524568|Neck vessels CT angiogram W contrast IV
C1524568|Multisection^W contrast Intravenous:Finding:Point in time:Neck>Vessels:Document:Computerized Tomography.angio
C1524568|Multisection^W contrast IV:Find:Pt:Neck>Vessels:Doc:CT.angio
C1524585|Should MRI W contr IV
C1524585|Shoulder MRI W contrast IV
C1524585|Multisection^W contrast IV:Find:Pt:Shoulder:Doc:MRI
C1524585|Multisection^W contrast Intravenous:Finding:Point in time:Shoulder:Document:MRI
C1524208|Finger third X-ray AP single view
C1524208|Finger.3rd XR AP 1V
C1524208|View AP:Find:Pt:Finger.third:Doc:XR
C1524208|View AP:Finding:Point in time:Finger.third:Document:XR
C1524214|Knee X-ray AP single view
C1524214|Knee XR AP 1V
C1524214|View AP:Find:Pt:Knee:Doc:XR
C1524214|View AP:Finding:Point in time:Knee:Document:XR
C1524289|Fluoroscopy Guidance for biopsy of Abdomen
C1524289|Abd Flr Bx guid
C1524289|Guidance for biopsy:Finding:Point in time:Abdomen:Document:XR.fluor
C1524289|Guidance for biopsy:Find:Pt:Abdomen:Doc:XR.fluor
C1524292|CT Guidance for biopsy of Breast
C1524292|Brst CT Bx guid
C1524292|Guidance for biopsy:Find:Pt:Breast:Doc:CT
C1524292|Guidance for biopsy:Finding:Point in time:Breast:Document:Computerized Tomography
C1524588|Should-R MRI W contr IV
C1524588|Shoulder - right MRI W contrast IV
C1524588|Multisection^W contrast Intravenous:Finding:Point in time:Shoulder.right:Document:MRI
C1524588|Multisection^W contrast IV:Find:Pt:Shoulder.right:Doc:MRI
C1524126|Breast - left MRI WO and W contrast IV
C1524126|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast.left:Document:MRI
C1524126|Multisection^WO & W contrast IV:Find:Pt:Breast.left:Doc:MRI
C1524126|Brst-L MRI WO+W contr IV
C1524313|CT Guidance for drainage of Anus
C1524313|Anus CT Drain guid
C1524313|Guidance for drainage:Find:Pt:Pelvis>Anus:Doc:CT
C1524313|Guidance for drainage:Finding:Point in time:Pelvis>Anus:Document:Computerized Tomography
C1524990|Brst-L Mam 2V
C1524990|Breast - left Mammogram 2 views
C1524990|Views 2:Finding:Point in time:Breast.left:Document:Mam
C1524990|Views 2:Find:Pt:Breast.left:Doc:Mam
C1524998|Elbow - left X-ray 2 views
C1524998|Elbow-L XR 2V
C1524998|Views 2:Find:Pt:Elbow.left:Doc:XR
C1524998|Views 2:Finding:Point in time:Elbow.left:Document:XR
C1524157|Radius+Ulna-Bl XR 2V
C1524157|Radius - bilateral and Ulna - bilateral X-ray 2 views
C1524157|Views 2:Find:Pt:Radius.bilateral+Ulna.bilateral:Doc:XR
C1524157|Views 2:Finding:Point in time:Radius.bilateral+Ulna.bilateral:Document:XR
C1525020|L-spine XR 7V
C1525020|Views 7:Find:Pt:Spine.lumbar:Doc:XR
C1525020|Views 7:Finding:Point in time:Spine.lumbar:Document:XR
C1525020|Lumbar spine X-ray 7 views
C1524354|Clavicle X-ray tomograph
C1524354|Clavicle XRTomo
C1524354|Multisection:Find:Pt:Clavicle:Doc:XR.tomo
C1524354|Multisection:Finding:Point in time:Clavicle:Document:XR.tomo
C1524385|Foot X-ray tomograph
C1524385|Ft XRTomo
C1524385|Multisection:Finding:Point in time:Foot:Document:XR.tomo
C1524385|Multisection:Find:Pt:Foot:Doc:XR.tomo
C1525041|Hip XR AP+Lat
C1525041|Hip X-ray AP and lateral
C1525041|Views AP & lateral:Finding:Point in time:Hip:Document:XR
C1525041|Views AP & lateral:Find:Pt:Hip:Doc:XR
C1524417|Upper arm - left MRI
C1524417|Upper arm-L MRI
C1524417|Multisection:Finding:Point in time:Upper arm.left:Document:MRI
C1524417|Multisection:Find:Pt:Upper arm.left:Doc:MRI
C1524775|Sacrum CT WO and W contrast IV
C1524775|Multisection^WO & W contrast IV:Find:Pt:Sacrum:Doc:CT
C1524775|Sacrum CT WO+W contr IV
C1524775|Multisection^WO & W contrast Intravenous:Finding:Point in time:Sacrum:Document:Computerized Tomography
C1524789|Spleen MRI WO+W contr IV
C1524789|Multisection^WO & W contrast IV:Find:Pt:Spleen:Doc:MRI
C1524789|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spleen:Document:MRI
C1524789|Spleen MRI WO and W contrast IV
C1524792|Thyroid MRI WO and W contrast IV
C1524792|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thyroid:Document:MRI
C1524792|Multisection^WO & W contrast IV:Find:Pt:Thyroid:Doc:MRI
C1524792|Thyroid MRI WO+W contr IV
C1524803|IVC MRI WO+W contr IV
C1524803|Multisection^WO & W contrast IV:Find:Pt:Vena cava.inferior:Doc:MRI
C1524803|Inferior vena cava MRI WO and W contrast IV
C1524803|Multisection^WO & W contrast Intravenous:Finding:Point in time:Vena cava.inferior:Document:MRI
C1524679|Elbow-L XR Obl
C1524679|Elbow - left X-ray oblique
C1524679|Views oblique:Finding:Point in time:Elbow.left:Document:XR
C1524679|Views oblique:Find:Pt:Elbow.left:Doc:XR
C1525086|Chest XR PA+Lat+Obl+Lordotic
C1525086|Chest X-ray PA and lateral and oblique and lordotic
C1525086|Views PA & lateral & oblique & lordotic:Find:Pt:Chest:Doc:XR
C1525086|Views PA & lateral & oblique & lordotic:Finding:Point in time:Chest:Document:XR
C1830205|Sinuses CT limited WO contrast
C1830205|Sinuses CT Ltd WO contr
C1830205|Multisection limited^WO contrast:Find:Pt:Head>Sinuses:Doc:CT
C1830205|Multisection limited^WO contrast:Finding:Point in time:Head>Sinuses:Document:Computerized Tomography
C1830235|Deprecated CBD XR Stone rem guid W contr
C1830235|Guidance for stone removal^W contrast intra biliary duct:Finding:Point in time:Biliary duct.common:Narrative:XR
C1830235|Guidance for stone removal^W contrast intra biliary duct:Find:Pt:Biliary duct.common:Nar:XR
C1830235|Deprecated X-ray Guidance for stone removal of Biliary duct common-- W contrast intra biliary duct
C1830248|Ankle-R XR GE 3V
C1830248|Ankle - right X-ray GE 3 views
C1830248|Views GE 3:Find:Pt:Ankle.right:Doc:XR
C1830248|Views GE 3:Finding:Point in time:Ankle.right:Document:XR
C1830250|Should-Bl XR AP+Transthoracic
C1830250|Shoulder - bilateral X-ray AP and transthoracic
C1830250|Views AP & transthoracic:Find:Pt:Shoulder.bilateral:Doc:XR
C1830250|Views AP & transthoracic:Finding:Point in time:Shoulder.bilateral:Document:XR
C1831075|Knee-R XR LE 4V
C1831075|Knee - right X-ray LE 4 views
C1831075|Views LE 4:Finding:Point in time:Knee.right:Document:XR
C1831075|Views LE 4:Find:Pt:Knee.right:Doc:XR
C1830073|Mandible X-ray GE 4 views
C1830073|Mandible XR GE 4V
C1830073|Views GE 4:Finding:Point in time:Mandible:Document:XR
C1830073|Views GE 4:Find:Pt:Mandible:Doc:XR
C1830076|L-spine XR GE 4V
C1830076|Views GE 4:Find:Pt:Spine.lumbar:Doc:XR
C1830076|Views GE 4:Finding:Point in time:Spine.lumbar:Document:XR
C1830076|Lumbar spine X-ray GE 4 views
C1715379|Retroperitoneum CT FNA Asp
C1715379|Guidance for aspiration.fine needle:Find:Pt:Abdomen>Retroperitoneum:Doc:CT
C1715379|CT Guidance for fine needle aspiration of Retroperitoneum
C1715379|Guidance for aspiration.fine needle:Finding:Point in time:Abdomen>Retroperitoneum:Document:Computerized Tomography
C1715385|T-spine CT WO+W contr IT
C1715385|Multisection^WO & W contrast IT:Find:Pt:Spine.thoracic:Doc:CT
C1715385|Multisection^WO & W contrast Intrathecal:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C1715385|Thoracic spine CT WO and W contrast IT
C1715386|L-spine CT WO+W contr IT
C1715386|Multisection^WO & W contrast Intrathecal:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1715386|Multisection^WO & W contrast IT:Find:Pt:Spine.lumbar:Doc:CT
C1715386|Lumbar spine CT WO and W contrast IT
C1715392|Mammogram Guidance for percutaneous needle biopsy of Breast
C1715392|Brst Mam PC Bx needle guid
C1715392|Guidance for percutaneous biopsy.needle:Find:Pt:Breast:Doc:Mam
C1715392|Guidance for percutaneous biopsy.needle:Finding:Point in time:Breast:Document:Mam
C1715413|Parathyroid RI W Tc99mMIBI IV
C1715413|Parathyroid Scan W Tc-99m Sestamibi IV
C1715413|Views^W Tc-99m Sestamibi Intravenous:Finding:Point in time:Parathyroid:Document:Radnuc
C1715413|Views^W Tc-99m Sestamibi IV:Find:Pt:Parathyroid:Doc:Radnuc
C1717315|US Guidance for biopsy of Abdomen retroperitoneum
C1717315|Abd.reper US Bx guid
C1717315|Guidance for biopsy:Finding:Point in time:Abdomen.retroperitoneum:Document:Ultrasound
C1717315|Guidance for biopsy:Find:Pt:Abdomen.retroperitoneum:Doc:US
C1715446|SIJ XR 2V or 3V
C1715446|Sacroiliac Joint X-ray 2 or 3 views
C1715446|Views 2 or 3:Find:Pt:Sacroiliac joint:Doc:XR
C1715446|Views 2 or 3:Finding:Point in time:Sacroiliac joint:Document:XR
C1635069|GB XR W 2x dose contr PO
C1635069|Gallbladder X-ray W double dose contrast PO
C1635069|Views^W double dose contrast PO:Find:Pt:Gallbladder:Doc:XR
C1635069|Views^W double dose contrast Oral:Finding:Point in time:Gallbladder:Document:XR
C1645329|Multisection transvaginal:Find:Pt:XXX:Doc:MRI
C1645329|MRI Transvag
C1645329|Transvaginal MRI
C1645329|Multisection transvaginal:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1632802|Foot sesamoid bones - bilateral X-ray axial
C1632802|View axial:Finding:Point in time:Foot.sesamoid bones.bilateral:Document:XR
C1632802|View axial:Find:Pt:Foot.sesamoid bones.bilateral:Doc:XR
C1632802|Ft.Sesamoids-Bl XR Axial
C1714907|Ovary - bilateral MRI
C1714907|Multisection:Find:Pt:Ovary.bilateral:Doc:MRI
C1714907|Multisection:Finding:Point in time:Ovary.bilateral:Document:MRI
C1714907|Ovary-Bl MRI
C1714926|Deprecated Unspecified body region CT dynamic W contrast IV
C1714926|Deprecated XXX CT Dyn W contr IV
C1714926|Multisection dynamic^W contrast IV:Find:Pt:XXX:Doc:CT
C1714926|Multisection dynamic^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1706619|Deprecated Finger.5th-L XR GE 3V
C1706619|Views GE 3:Find:Pt:Finger.fifth.left:Nar:XR
C1706619|Deprecated Finger fifth Left X-ray GE 3 views
C1706619|Views GE 3:Finding:Point in time:Finger.fifth.left:Narrative:XR
C1705863|Deprecated Finger.2nd-R XR GE 3V
C1705863|Views GE 3:Find:Pt:Finger.second.right:Nar:XR
C1705863|Deprecated Finger second Right X-ray GE 3 views
C1705863|Views GE 3:Finding:Point in time:Finger.second.right:Narrative:XR
C1715018|Hrt RI for Infarct Ql W RNC IV
C1715018|Heart Scan for infarct qualitative
C1715018|Views for infarct qualitative^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1715018|Views for infarct qualitative^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1715090|Vein-L XRA Thrombect guid W contr IV
C1715090|Fluoroscopic angiogram Guidance for thrombectomy of Vein - left-- W contrast IV
C1715090|Guidance for thrombectomy^W contrast IV:Find:Pt:Vein.left:Doc:XR.fluor.angio
C1715090|Guidance for thrombectomy^W contrast Intravenous:Finding:Point in time:Vein.left:Document:XR.fluor.angio
C1637278|Ankle-Bl XR AP+Lat+Obl W Stress
C1637278|Ankle - bilateral X-ray AP and lateral and oblique W manual stress
C1637278|Views AP & lateral & oblique^W manual stress:Find:Pt:Ankle.bilateral:Doc:XR
C1637278|Views AP & lateral & oblique^W manual stress:Finding:Point in time:Ankle.bilateral:Document:XR
C1626322|Upper extremity vessel graft - left US.doppler
C1626322|UE ves graft-L DOP
C1626322|Multisection:Find:Pt:Upper extremity vessel graft.left:Doc:US.doppler
C1626322|Multisection:Finding:Point in time:Upper extremity vessel graft.left:Document:Ultrasound.doppler
C1626174|US Guidance for aspiration of Thyroid
C1626174|Thyroid US Asp guid
C1626174|Guidance for aspiration:Finding:Point in time:Thyroid:Document:Ultrasound
C1626174|Guidance for aspiration:Find:Pt:Thyroid:Doc:US
C1641530|Shoulder - right X-ray portable
C1641530|Should-R XR port
C1641530|Views portable:Find:Pt:Shoulder.right:Doc:XR
C1641530|Views portable:Finding:Point in time:Shoulder.right:Document:XR
C1643596|Chest XR R-Obl+L-Obl
C1643596|Chest X-ray right oblique and left oblique
C1643596|Views R-oblique & L-oblique:Finding:Point in time:Chest:Document:XR
C1643596|Views R-oblique & L-oblique:Find:Pt:Chest:Doc:XR
C1631261|CT Guidance for needle biopsy of Pancreas
C1631261|Pancreas CT Bx needle guid
C1631261|Guidance for biopsy.needle:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C1631261|Guidance for biopsy.needle:Find:Pt:Abdomen>Pancreas:Doc:CT
C1632226|RI for Tumor W Tl-201 IV
C1632226|Scan for tumor W Tl-201 IV
C1632226|Views for tumor^W Tl-201 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1632226|Views for tumor^W Tl-201 IV:Find:Pt:^Patient:Doc:Radnuc
C1624132|Unspecified body region Fluoroscopy Greater than 1 hour
C1624132|XXX Flr >1h
C1624132|View:Find:Gt 1H:XXX:Doc:XR.fluor
C1624132|View:Finding:Greater than 1 hour:To be specified in another part of the message:Document:XR.fluor
C1977258|XXX MRI W contr IV
C1977258|Unspecified body region MRI W contrast IV
C1977258|Multisection^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1977258|Multisection^W contrast IV:Find:Pt:XXX:Doc:MRI
C1954303|Upper extremity vein - left US
C1954303|UE v-L US
C1954303|Multisection:Finding:Point in time:Upper extremity vein.left:Document:Ultrasound
C1954303|Multisection:Find:Pt:Upper extremity vein.left:Doc:US
C1954311|Views:Finding:Point in time:Skull.base:Narrative:XR
C1954311|Skull.base XR
C1954311|Skull.base X-ray
C1954311|Views:Finding:Point in time:Skull.base:Document:XR
C1954311|Views:Find:Pt:Skull.base:Doc:XR
C1953328|LE aa-R XRA W contr IA
C1953328|Lower extremity arteries - right Fluoroscopic angiogram W contrast IA
C1953328|Views^W contrast IA:Find:Pt:Lower extremity arteries.right:Doc:XR.fluor.angio
C1953328|Views^W contrast Intra-arterial:Finding:Point in time:Lower extremity arteries.right:Document:XR.fluor.angio
C1953945|T-spine MRI W contr IT
C1953945|Multisection^W contrast IT:Find:Pt:Spine.thoracic:Doc:MRI
C1953945|Multisection^W contrast Intrathecal:Finding:Point in time:Spine.thoracic:Document:MRI
C1953945|Thoracic spine MRI W contrast IT
C1953955|Orbit CT W contr IV
C1953955|Orbit CT W contrast IV
C1953955|Multisection^W contrast IV:Find:Pt:Head>Orbit:Doc:CT
C1953955|Multisection^W contrast Intravenous:Finding:Point in time:Head>Orbit:Document:Computerized Tomography
C3533805|Multisection^W contrast IV:Find:Pt:Toes.right:Doc:MRI
C3533805|Toes - right MRI W contrast IV
C3533805|Multisection^W contrast Intravenous:Finding:Point in time:Toes.right:Document:MRI
C3533805|Toes-R MRI W contr IV
C3533803|Multisection^WO contrast:Find:Pt:Toes.left:Doc:MRI
C3533803|Toes-L MRI WO contr
C3533803|Toes - left MRI WO contrast
C3533803|Multisection^WO contrast:Finding:Point in time:Toes.left:Document:MRI
C3655083|Multisection & physiologic artery study:Find:Pt:Extremity arteries.bilateral:Doc:US.doppler
C3655083|Extremity arteries - bilateral US.doppler Multisection and physiologic artery study
C3655083|Multisection & physiologic artery study:Finding:Point in time:Extremity arteries.bilateral:Document:Ultrasound.doppler
C3655083|Extr aa-Bl DOP +Phys stdy
C3655081|Multisection & physiologic artery study^at rest & W exercise:Finding:Point in time:Extremity arteries.bilateral:Document:Ultrasound.doppler
C3655081|Multisection & physiologic artery study^at rest & W exercise:Find:Pt:Extremity arteries.bilateral:Doc:US.doppler
C3655081|Extr aa-Bl DOP +Phys stdy Rest+excz
C3655081|Extremity arteries - bilateral US.doppler Multisection and physiologic artery study at rest and with exercise
C3262948|Liver Flr Bx needle guid
C3262948|Fluoroscopy Guidance for needle biopsy of Liver
C3262948|Guidance for biopsy.needle:Finding:Point in time:Liver:Document:XR.fluor
C3262948|Guidance for biopsy.needle:Find:Pt:Liver:Doc:XR.fluor
C3262955|Hip Flr Drain guid
C3262955|Fluoroscopy Guidance for drainage of Hip
C3262955|Guidance for drainage:Find:Pt:Hip:Doc:XR.fluor
C3262955|Guidance for drainage:Finding:Point in time:Hip:Document:XR.fluor
C3262956|Iliac a XRA Stent plac guid
C3262956|Fluoroscopic angiogram Guidance for placement of stent in Iliac artery
C3262956|Guidance for placement of stent:Find:Pt:Iliac artery:Doc:XR.fluor.angio
C3262956|Guidance for placement of stent:Finding:Point in time:Iliac artery:Document:XR.fluor.angio
C3262995|Forearm - bilateral MRI W contrast IV
C3262995|Forearm-Bl MRI W contr IV
C3262995|Multisection^W contrast IV:Find:Pt:Forearm.bilateral:Doc:MRI
C3262995|Multisection^W contrast Intravenous:Finding:Point in time:Forearm.bilateral:Document:MRI
C3263078|Shoulder X-ray AP and Y
C3263078|Should XR AP+Y
C3263078|Views AP & Y:Find:Pt:Shoulder:Doc:XR
C3263078|Views AP & Y:Finding:Point in time:Shoulder:Document:XR
C3263086|T-spine XR 2V stand
C3263086|Views 2^standing:Find:Pt:Spine.thoracic:Doc:XR
C3263086|Views 2^standing:Finding:Point in time:Spine.thoracic:Document:XR
C3263086|Thoracic spine X-ray 2 views standing
C3263098|Salivary gland US
C3263098|Multisection:Find:Pt:Salivary gland:Doc:US
C3263098|Multisection:Finding:Point in time:Salivary gland:Document:Ultrasound
C3263106|Fluoroscopy Guidance for aspiration of cyst of Bone
C3263106|Bone Flr Cyst Asp guid
C3263106|Guidance for aspiration of cyst:Find:Pt:Bone:Doc:XR.fluor
C3263106|Guidance for aspiration of cyst:Finding:Point in time:Bone:Document:XR.fluor
C3263206|Ovary US
C3263206|Multisection:Find:Pt:Ovary:Doc:US
C3263206|Multisection:Finding:Point in time:Ovary:Document:Ultrasound
C3262896|XXX Flr Bx CN guid
C3262896|Fluoroscopy Guidance for core needle biopsy of Unspecified body region
C3262896|Guidance for biopsy.core needle:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C3262896|Guidance for biopsy.core needle:Find:Pt:XXX:Doc:XR.fluor
C0487981|Chest XR Diam AP
C0487981|Diameter.anterior-posterior:Len:Pt:Chest:Qn:XR
C0487981|Chest X-ray Diameter.anterior-posterior
C0487981|Diameter.anterior-posterior:Length:Point in time:Chest:Quantitative:XR
C0944167|Joint MRI
C0944167|Multisection:Finding:Point in time:Joint:Document:MRI
C0944167|Multisection:Find:Pt:Joint:Doc:MRI
C0942198|Multisection^WO & W contrast Intravenous:Finding:Point in time:Elbow.left:Document:MRI
C0942198|Multisection^WO & W contrast IV:Find:Pt:Elbow.left:Doc:MRI
C0942198|Elbow-L MRI WO+W contr IV
C0942198|Elbow - left MRI WO and W contrast IV
C0942244|Forearm - right MRI
C0942244|Forearm-R MRI
C0942244|Multisection:Find:Pt:Forearm.right:Doc:MRI
C0942244|Multisection:Finding:Point in time:Forearm.right:Document:MRI
C0942260|Should-Bl US
C0942260|Shoulder - bilateral US
C0942260|Multisection:Finding:Point in time:Shoulder.bilateral:Document:Ultrasound
C0942260|Multisection:Find:Pt:Shoulder.bilateral:Doc:US
C0942294|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - right
C0942294|Cent v-R XRA LT per cath plac guid
C0942294|Guidance for placement of longterm peripheral catheter:Find:Pt:Central vein.right:Doc:XR.fluor.angio
C0942294|Guidance for placement of longterm peripheral catheter:Finding:Point in time:Central vein.right:Document:XR.fluor.angio
C0942372|Knee - left X-ray 2 views
C0942372|Knee-L XR 2V
C0942372|Views 2:Finding:Point in time:Knee.left:Document:XR
C0942372|Views 2:Find:Pt:Knee.left:Doc:XR
C0882065|Peripheral vessel US.doppler Peripheral plane
C0882065|Periph ves DOP Periph plane
C0882065|Peripheral plane:Find:Pt:Peripheral vessel:Doc:US.doppler
C0882065|Peripheral plane:Finding:Point in time:Peripheral vessel:Document:Ultrasound.doppler
C0882089|Shoulder MRI WO and W contrast IV
C0882089|Multisection^WO & W contrast IV:Find:Pt:Shoulder:Doc:MRI
C0882089|Should MRI WO+W contr IV
C0882089|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder:Document:MRI
C0882098|Sinuses MRI W contr IV
C0882098|Sinuses MRI W contrast IV
C0882098|Multisection^W contrast Intravenous:Finding:Point in time:Sinuses:Document:MRI
C0882098|Multisection^W contrast IV:Find:Pt:Sinuses:Doc:MRI
C0882552|C-spine CT
C0882552|Multisection:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C0882552|Multisection:Find:Pt:Spine.cervical:Doc:CT
C0882552|Cervical spine CT
C0882138|L-spine MRI W anesthesia
C0882138|Multisection^W anesthesia:Find:Pt:Spine.lumbar:Doc:MRI
C0882138|Multisection^W anesthesia:Finding:Point in time:Spine.lumbar:Document:MRI
C0882138|Lumbar spine MRI W anesthesia
C0882173|Urethra Fluoroscopy W contrast intra urethra
C0882173|Urth Flr W contr intra ureth
C0882173|Views^W contrast intra urethra:Find:Pt:Urethra:Doc:XR.fluor
C0882173|Views^W contrast intra urethra:Finding:Point in time:Urethra:Document:XR.fluor
C0882183|Guidance for placement of large bore catheter into vessel in Central vein
C0882183|Centl v LB Cath plac guid into ves
C0882183|Guidance for placement of large bore catheter into vessel:Find:Pt:Central vein:Doc
C0882183|Guidance for placement of large bore catheter into vessel:Finding:Point in time:Central vein:Document
C0942100|Carotid artery - bilateral Fluoroscopic angiogram W contrast IA
C0942100|Carot a-Bl XRA W contr IA
C0942100|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.bilateral:Document:XR.fluor.angio
C0942100|Views^W contrast IA:Find:Pt:Carotid artery.bilateral:Doc:XR.fluor.angio
C0942132|Lower extremity - right X-ray
C0942132|LE-R XR
C0942132|Views:Find:Pt:Lower extremity.right:Doc:XR
C0942132|Views:Finding:Point in time:Lower extremity.right:Document:XR
C0881779|Ankle MRI
C0881779|Multisection:Finding:Point in time:Ankle:Narrative:MRI
C0881779|Multisection:Find:Pt:Ankle:Doc:MRI
C0881779|Multisection:Finding:Point in time:Ankle:Document:MRI
C0881866|View AP L-lateral-decubitus:Finding:Point in time:Chest:Narrative:XR
C0881866|Chest XR AP L-Lat Decub
C0881866|Chest X-ray AP left lateral-decubitus
C0881866|View AP L-lateral-decubitus:Find:Pt:Chest:Doc:XR
C0881866|View AP L-lateral-decubitus:Finding:Point in time:Chest:Document:XR
C0881959|Views^at rest & W Tl-201 Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C0881959|Hrt RI Rest+W Tl201 IV
C0881959|Heart Scan at rest and W Tl-201 IV
C0881959|Views^at rest & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C0881959|Views^at rest & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1114486|XXX MRI RT guid W contr IV
C1114486|MRI Guidance for radiation treatment of Unspecified body region-- W contrast IV
C1114486|Guidance for radiation treatment^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1114486|Guidance for radiation treatment^W contrast IV:Find:Pt:XXX:Doc:MRI
C1114540|C-spine XR AP+Lat port
C1114540|Views AP & lateral portable:Finding:Point in time:Spine.cervical:Document:XR
C1114540|Views AP & lateral portable:Find:Pt:Spine.cervical:Doc:XR
C1114540|Cervical spine X-ray AP and lateral portable
C1114565|T-spine XR AP V1 port
C1114565|View AP portable:Find:Pt:Spine.thoracic:Doc:XR
C1114565|View AP portable:Finding:Point in time:Spine.thoracic:Document:XR
C1114565|Thoracic spine X-ray AP portable single view
C1114572|Acetabulum - bilateral X-ray portable
C1114572|Acetabulum-Bl XR port
C1114572|Views portable:Find:Pt:Acetabulum.bilateral:Doc:XR
C1114572|Views portable:Finding:Point in time:Acetabulum.bilateral:Document:XR
C1114583|L-spine XR Obl 1V
C1114583|View oblique:Find:Pt:Spine.lumbar:Doc:XR
C1114583|View oblique:Finding:Point in time:Spine.lumbar:Document:XR
C1114583|Lumbar spine X-ray oblique single view
C1114422|C-spine CT WO contr
C1114422|Multisection^WO contrast:Find:Pt:Spine.cervical:Doc:CT
C1114422|Multisection^WO contrast:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C1114422|Cervical spine CT WO contrast
C1114433|Pancreas CT FNA Asp
C1114433|CT Guidance for fine needle aspiration of Pancreas
C1114433|Guidance for aspiration.fine needle:Find:Pt:Abdomen>Pancreas:Doc:CT
C1114433|Guidance for aspiration.fine needle:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C1114451|Pelvic vessels CT angiogram WO and W contrast IV
C1114451|Multisection^WO & W contrast IV:Find:Pt:Pelvis>Vessels:Doc:CT.angio
C1114451|Pelv ves CT.Angio WO+W contr IV
C1114451|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pelvis>Vessels:Document:Computerized Tomography.angio
C1543437|Ribs posterior - bilateral X-ray
C1543437|Ribs post-Bl XR
C1543437|Views:Finding:Point in time:Ribs.posterior.bilateral:Document:XR
C1543437|Views:Find:Pt:Ribs.posterior.bilateral:Doc:XR
C1543448|Wrist-R XR 3V+Radial Deviation
C1543448|Wrist - right X-ray 3 views and radial deviation
C1543448|Views 3 & radial deviation:Find:Pt:Wrist.right:Doc:XR
C1543448|Views 3 & radial deviation:Finding:Point in time:Wrist.right:Document:XR
C2718315|Views & oblique:Finding:Point in time:Elbow.right:Narrative:XR
C2718315|Elbow-R XR +Obl
C2718315|Elbow - right X-ray and oblique
C2718315|Views & oblique:Finding:Point in time:Elbow.right:Document:XR
C2718315|Views & oblique:Find:Pt:Elbow.right:Doc:XR
C1543747|Lung RI Ltd W RNC IV
C1543747|Lung Scan limited
C1543747|Views limited^W radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1543747|Views limited^W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1543461|Knee-R XR 2V+Tunnel
C1543461|Knee - right X-ray 2 views and tunnel
C1543461|Views 2 & tunnel:Finding:Point in time:Knee.right:Document:XR
C1543461|Views 2 & tunnel:Find:Pt:Knee.right:Doc:XR
C1543489|T-spine XR +Swimmers
C1543489|Views & Swimmers:Find:Pt:Spine.thoracic:Doc:XR
C1543489|Views & Swimmers:Finding:Point in time:Spine.thoracic:Document:XR
C1543489|Thoracic spine X-ray and Swimmers
C1543491|Gastrointestine US
C1543491|GI US
C1543491|Multisection:Find:Pt:Gastrointestine:Doc:US
C1543491|Multisection:Finding:Point in time:Gastrointestine:Document:Ultrasound
C1543873|RI for Tumor Ltd W Ga-67 IV
C1543873|Views for tumor limited^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543873|Views for tumor limited^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543873|Scan for tumor limited W Ga-67 IV
C1543520|UE ves-R DOP
C1543520|Upper extremity vessels - right US.doppler
C1543520|Multisection:Finding:Point in time:Upper extremity vessels.right:Document:Ultrasound.doppler
C1543520|Multisection:Find:Pt:Upper extremity vessels.right:Doc:US.doppler
C1543159|Orbit+Face MRI W contr IV
C1543159|Orbit and Face MRI W contrast IV
C1543159|Multisection^W contrast IV:Find:Pt:Orbit+Face:Doc:MRI
C1543159|Multisection^W contrast Intravenous:Finding:Point in time:Orbit+Face:Document:MRI
C1543568|Ribs upper post-R XR
C1543568|Ribs upper posterior - right X-ray
C1543568|Views:Find:Pt:Ribs.upper.posterior.right:Doc:XR
C1543568|Views:Finding:Point in time:Ribs.upper.posterior.right:Document:XR
C1543190|Ft XR AP+Lat
C1543190|Foot X-ray AP and lateral
C1543190|Views AP & lateral:Find:Pt:Foot:Doc:XR
C1543190|Views AP & lateral:Finding:Point in time:Foot:Document:XR
C1543688|Vein - bilateral Scan
C1543688|Vein-Bl RI W RNC IV
C1543688|Views^W radionuclide IV:Find:Pt:Vein.bilateral:Doc:Radnuc
C1543688|Views^W radionuclide Intravenous:Finding:Point in time:Vein.bilateral:Document:Radnuc
C1524261|Patella-R XR AP+Lat+Sunrise
C1524261|Patella - right X-ray AP and lateral and Sunrise
C1524261|Views AP & lateral & Sunrise:Find:Pt:Patella.right:Doc:XR
C1524261|Views AP & lateral & Sunrise:Finding:Point in time:Patella.right:Document:XR
C1526750|Should-R XR Grashey+Outlet+Serendipity
C1526750|Shoulder - right X-ray Grashey and outlet and Serendipity
C1526750|Views Grashey & outlet & Serendipity:Find:Pt:Shoulder.right:Doc:XR
C1526750|Views Grashey & outlet & Serendipity:Finding:Point in time:Shoulder.right:Document:XR
C1543709|Hrt SPECT W Tc99mTF IV
C1543709|Heart SPECT W Tc-99m Tetrofosmin IV
C1543709|Multisection^W Tc-99m Tetrofosmin IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543709|Multisection^W Tc-99m Tetrofosmin Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543734|SPECT Ltd W Ga-67 IV
C1543734|Multisection limited^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543734|Multisection limited^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543734|SPECT limited W Ga-67 IV
C1526808|Knee - left X-ray 4 views standing
C1526808|Knee-L XR 4V stand
C1526808|Views 4^standing:Find:Pt:Knee.left:Doc:XR
C1526808|Views 4^standing:Finding:Point in time:Knee.left:Document:XR
C1526817|Ankle aa-L XRA W contr IA
C1526817|Ankle arteries - left Fluoroscopic angiogram W contrast IA
C1526817|Views^W contrast IA:Find:Pt:Ankle arteries.left:Doc:XR.fluor.angio
C1526817|Views^W contrast Intra-arterial:Finding:Point in time:Ankle arteries.left:Document:XR.fluor.angio
C1524433|Mandible XRTomo
C1524433|Mandible X-ray tomograph
C1524433|Multisection:Find:Pt:Mandible:Doc:XR.tomo
C1524433|Multisection:Finding:Point in time:Mandible:Document:XR.tomo
C1524173|Sacrum CT
C1524173|Multisection:Finding:Point in time:Sacrum:Document:Computerized Tomography
C1524173|Multisection:Find:Pt:Sacrum:Doc:CT
C1524181|C-spine XRTomo
C1524181|Multisection:Find:Pt:Spine.cervical:Doc:XR.tomo
C1524181|Multisection:Finding:Point in time:Spine.cervical:Document:XR.tomo
C1524181|Cervical spine X-ray tomograph
C1524184|Sternum MRI
C1524184|Multisection:Find:Pt:Sternum:Doc:MRI
C1524184|Multisection:Finding:Point in time:Sternum:Document:MRI
C1524188|Lower leg - right MRI
C1524188|Lower leg-R MRI
C1524188|Multisection:Finding:Point in time:Lower leg.right:Document:MRI
C1524188|Multisection:Find:Pt:Lower leg.right:Doc:MRI
C1524818|TA MRI.Angio WO contr
C1524818|Aorta thoracic MRI angiogram WO contrast
C1524818|Multisection^WO contrast:Finding:Point in time:Aorta.thoracic:Document:MRI.angio
C1524818|Multisection^WO contrast:Find:Pt:Aorta.thoracic:Doc:MRI.angio
C1524820|Face MRI WO contr
C1524820|Face MRI WO contrast
C1524820|Multisection^WO contrast:Finding:Point in time:Face:Document:MRI
C1524820|Multisection^WO contrast:Find:Pt:Face:Doc:MRI
C1524838|LE-L MRI WO contr
C1524838|Lower extremity - left MRI WO contrast
C1524838|Multisection^WO contrast:Finding:Point in time:Lower extremity.left:Document:MRI
C1524838|Multisection^WO contrast:Find:Pt:Lower extremity.left:Doc:MRI
C1524850|Thigh-R MRI WO contr
C1524850|Thigh - right MRI WO contrast
C1524850|Multisection^WO contrast:Find:Pt:Thigh.right:Doc:MRI
C1524850|Multisection^WO contrast:Finding:Point in time:Thigh.right:Document:MRI
C1525106|Toe MRI
C1525106|Multisection:Find:Pt:Toe:Doc:MRI
C1525106|Multisection:Finding:Point in time:Toe:Document:MRI
C1524459|Multisection^W contrast IS:Find:Pt:Ankle:Doc:MRI
C1524459|Multisection^W contrast Intrasynovial:Finding:Point in time:Ankle:Document:MRI
C1524459|Ankle MRI W contrast IS
C1524459|Ankle MRI W contr IS
C1525290|Ribs-Bl XR AP 1V
C1525290|Ribs - bilateral X-ray AP single view
C1525290|View AP:Finding:Point in time:Ribs.bilateral:Document:XR
C1525290|View AP:Find:Pt:Ribs.bilateral:Doc:XR
C1525293|Should-L XR AP+West Point+Outlet
C1525293|Shoulder - left X-ray AP and West Point and outlet
C1525293|Views AP & West Point & outlet:Finding:Point in time:Shoulder.left:Document:XR
C1525293|Views AP & West Point & outlet:Find:Pt:Shoulder.left:Doc:XR
C1525301|Deprecated View decubitus:Finding:Point in time:Abdomen:Narrative:XR
C1525301|Deprecated View decubitus
C1525301|View decubitus:Find:Pt:Abdomen:Nar:XR
C1525301|Deprecated Abd XR decubitus
C1525301|View decubitus:Finding:Point in time:Abdomen:Narrative:XR
C1525198|Ovary MRI W contr IV
C1525198|Ovary MRI W contrast IV
C1525198|Multisection^W contrast IV:Find:Pt:Ovary:Doc:MRI
C1525198|Multisection^W contrast Intravenous:Finding:Point in time:Ovary:Document:MRI
C1525216|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.joint.right:Doc:MRI
C1525216|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.joint.right:Document:MRI
C1525216|UE joint-R MRI WO+W contr IV
C1525216|Upper extremity joint - right MRI WO and W contrast IV
C1525260|Tib+Fib XR Obl
C1525260|Tibia and Fibula X-ray oblique
C1525260|Views oblique:Find:Pt:Tibia+Fibula:Doc:XR
C1525260|Views oblique:Finding:Point in time:Tibia+Fibula:Document:XR
C1524682|Knee - left X-ray PA standing
C1524682|Knee-L XR PA V1 stand
C1524682|View PA^standing:Find:Pt:Knee.left:Doc:XR
C1524682|View PA^standing:Finding:Point in time:Knee.left:Document:XR
C1524689|Deprecated Calcaneus - bilateral X-ray ski jump
C1524689|Deprecated Heel-Bl XR Ski Jump
C1524689|Views ski jump:Finding:Point in time:Calcaneus.bilateral:Document:XR
C1524689|Views ski jump:Find:Pt:Calcaneus.bilateral:Doc:XR
C1525475|XXX Flr of FB
C1525475|Unspecified body region Fluoroscopy of foreign body
C1525475|Views of foreign body:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1525475|Views of foreign body:Find:Pt:XXX:Doc:XR.fluor
C1525493|Should-L XR AP+Ax+Outlet
C1525493|Shoulder - left X-ray AP and axillary and outlet
C1525493|Views AP & axillary & outlet:Finding:Point in time:Shoulder.left:Document:XR
C1525493|Views AP & axillary & outlet:Find:Pt:Shoulder.left:Doc:XR
C1525507|Knee-Bl XR AP+Lat+Sunrise
C1525507|Knee - bilateral X-ray AP and lateral and Sunrise
C1525507|Views AP & lateral & Sunrise:Finding:Point in time:Knee.bilateral:Document:XR
C1525507|Views AP & lateral & Sunrise:Find:Pt:Knee.bilateral:Doc:XR
C1525537|Abd XR R-Obl+L-Obl
C1525537|Abdomen X-ray right oblique and left oblique
C1525537|Views R-oblique & L-oblique:Find:Pt:Abdomen:Doc:XR
C1525537|Views R-oblique & L-oblique:Finding:Point in time:Abdomen:Document:XR
C1525538|C-spine XR Obl+Lat W FE
C1525538|Views oblique & lateral^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C1525538|Views oblique & lateral^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C1525538|Cervical spine X-ray oblique and lateral W flexion and W extension
C1525569|Humerus X-ray portable
C1525569|Humerus XR port
C1525569|Views portable:Finding:Point in time:Humerus:Document:XR
C1525569|Views portable:Find:Pt:Humerus:Doc:XR
C1525573|Fem a+Popliteal a XRA W contr IA
C1525573|Femoral artery and Popliteal artery Fluoroscopic angiogram W contrast IA
C1525573|Views^W contrast IA:Find:Pt:Femoral artery+Popliteal artery:Doc:XR.fluor.angio
C1525573|Views^W contrast Intra-arterial:Finding:Point in time:Femoral artery+Popliteal artery:Document:XR.fluor.angio
C1525593|Jugular v XRA W contr IV
C1525593|Jugular vein Fluoroscopic angiogram W contrast IV
C1525593|Views^W contrast IV:Find:Pt:Jugular vein:Doc:XR.fluor.angio
C1525593|Views^W contrast Intravenous:Finding:Point in time:Jugular vein:Document:XR.fluor.angio
C1525646|Pelvis+L-spine XR 3V
C1525646|Pelvis and Spine Lumbar X-ray 3 views
C1525646|Views 3:Find:Pt:Pelvis+Spine.lumbar:Doc:XR
C1525646|Views 3:Finding:Point in time:Pelvis+Spine.lumbar:Document:XR
C1525649|L-spine+Sacrum+Coccyx XR 3V
C1525649|Spine Lumbar and Sacrum and Coccyx X-ray 3 views
C1525649|Views 3:Find:Pt:Spine.lumbar+Sacrum+Coccyx:Doc:XR
C1525649|Views 3:Finding:Point in time:Spine.lumbar+Sacrum+Coccyx:Document:XR
C1525679|Face+Zygomatic Arch XR
C1525679|Facial bones and Zygomatic arch X-ray
C1525679|Views:Find:Pt:Facial bones+Zygomatic arch:Doc:XR
C1525679|Views:Finding:Point in time:Facial bones+Zygomatic arch:Document:XR
C1525692|Toes - bilateral X-ray 2 views
C1525692|Toes-Bl XR 2V
C1525692|Views 2:Finding:Point in time:Toes.bilateral:Document:XR
C1525692|Views 2:Find:Pt:Toes.bilateral:Doc:XR
C1525712|Ac arch+VA-R XRA W contr IA
C1525712|Aortic arch and Vertebral artery - right Fluoroscopic angiogram W contrast IA
C1525712|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Vertebral artery.right:Document:XR.fluor.angio
C1525712|Views^W contrast IA:Find:Pt:Aortic arch+Vertebral artery.right:Doc:XR.fluor.angio
C1525715|Bronchial artery Fluoroscopic angiogram W contrast IA
C1525715|Bronchial a XRA W contr IA
C1525715|Views^W contrast IA:Find:Pt:Bronchial artery:Doc:XR.fluor.angio
C1525715|Views^W contrast Intra-arterial:Finding:Point in time:Bronchial artery:Document:XR.fluor.angio
C1525728|Celiac a+Gastric a-L+SMA XRA W contr IA
C1525728|Celiac artery and Gastric artery - left and Superior mesenteric artery Fluoroscopic angiogram W contrast IA
C1525728|Views^W contrast Intra-arterial:Finding:Point in time:Celiac artery+Gastric artery.left+Superior mesenteric artery:Document:XR.fluor.angio
C1525728|Views^W contrast IA:Find:Pt:Celiac artery+Gastric artery.left+Superior mesenteric artery:Doc:XR.fluor.angio
C1525794|VA-L XRA W contr IA
C1525794|Vertebral artery - left Fluoroscopic angiogram W contrast IA
C1525794|Views^W contrast Intra-arterial:Finding:Point in time:Vertebral artery.left:Document:XR.fluor.angio
C1525794|Views^W contrast IA:Find:Pt:Vertebral artery.left:Doc:XR.fluor.angio
C1525933|Pelvis ves XRA W contr
C1525933|Pelvis vessels Fluoroscopic angiogram W contrast
C1525933|Views^W contrast:Finding:Point in time:Pelvis vessels:Document:XR.fluor.angio
C1525933|Views^W contrast:Find:Pt:Pelvis vessels:Doc:XR.fluor.angio
C1525941|Pelvis XR AP+Inlet+Outlet
C1525941|Pelvis X-ray AP and inlet and outlet
C1525941|Views AP & inlet & outlet:Finding:Point in time:Pelvis:Document:XR
C1525941|Views AP & inlet & outlet:Find:Pt:Pelvis:Doc:XR
C1525803|Multisection^W contrast Intravenous:Finding:Point in time:Aortic stent:Document:Computerized Tomography.angio
C1525803|Deprecated Ac stent CT.Angio W contr IV
C1525803|Multisection^W contrast IV:Find:Pt:Aortic stent:Doc:CT.angio
C1525803|Deprecated Aortic stent CT angiogram W contrast IV
C1525817|Tib-L XR 10 Deg Cau Angle
C1525817|Tibia - left X-ray 10 degree caudal angle
C1525817|View 10 degree caudal angle:Find:Pt:Tibia.left:Doc:XR
C1525817|View 10 degree caudal angle:Finding:Point in time:Tibia.left:Document:XR
C1525957|Views^W contrast:Find:Pt:Abdomen>Renal vessels:Doc:XR.fluor.angio
C1525957|Views^W contrast:Finding:Point in time:Abdomen>Renal vessels:Document:XR.fluor.angio
C1525957|Abd>Renal vls XRA W contr
C1525957|Abdominal Renal vessels Fluoroscopic angiogram W contrast
C1525976|T+L-spine XR Scoli Lat stand
C1525976|Spine Thoracic and Lumbar X-ray scoliosis lateral standing
C1525976|View scoliosis lateral^standing:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1525976|View scoliosis lateral^standing:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1526030|Hand - right X-ray PA
C1526030|Hand-R XR PA V1
C1526030|View PA:Find:Pt:Hand.right:Doc:XR
C1526030|View PA:Finding:Point in time:Hand.right:Document:XR
C1526040|Hip-R XR AP+Lat Frog
C1526040|Hip - right X-ray AP and lateral frog
C1526040|Views AP & lateral frog:Finding:Point in time:Hip.right:Document:XR
C1526040|Views AP & lateral frog:Find:Pt:Hip.right:Doc:XR
C1526042|Hip-R XR AP 1V
C1526042|Hip - right X-ray AP single view
C1526042|View AP:Finding:Point in time:Hip.right:Document:XR
C1526042|View AP:Find:Pt:Hip.right:Doc:XR
C1526088|Ribs-R XR AP 1V
C1526088|Ribs - right X-ray AP single view
C1526088|View AP:Find:Pt:Ribs.right:Doc:XR
C1526088|View AP:Finding:Point in time:Ribs.right:Document:XR
C1526094|Scapula-R XR AP+Y
C1526094|Scapula - right X-ray AP and Y
C1526094|Views AP & Y:Finding:Point in time:Scapula.right:Document:XR
C1526094|Views AP & Y:Find:Pt:Scapula.right:Doc:XR
C1526136|Should XR Grashey
C1526136|Shoulder X-ray Grashey
C1526136|View Grashey:Finding:Point in time:Shoulder:Document:XR
C1526136|View Grashey:Find:Pt:Shoulder:Doc:XR
C1526176|Tib+Fib XR AP+Lat
C1526176|Tibia and Fibula X-ray AP and lateral
C1526176|Views AP & lateral:Finding:Point in time:Tibia+Fibula:Document:XR
C1526176|Views AP & lateral:Find:Pt:Tibia+Fibula:Doc:XR
C1526205|Pelvis aa+LE aa-Bl XRA W contr IA
C1526205|Pelvis arteries and Lower extremity arteries - bilateral Fluoroscopic angiogram W contrast IA
C1526205|Views^W contrast IA:Find:Pt:Pelvis arteries+Lower extremity arteries.bilateral:Doc:XR.fluor.angio
C1526205|Views^W contrast Intra-arterial:Finding:Point in time:Pelvis arteries+Lower extremity arteries.bilateral:Document:XR.fluor.angio
C1526254|Chest XR W Insp
C1526254|Chest X-ray W inspiration
C1526254|View^W inspiration:Find:Pt:Chest:Doc:XR
C1526254|View^W inspiration:Finding:Point in time:Chest:Document:XR
C1525141|Carot a US Ltd
C1525141|Carotid artery US limited
C1525141|Multisection limited:Finding:Point in time:Carotid artery:Document:Ultrasound
C1525141|Multisection limited:Find:Pt:Carotid artery:Doc:US
C1526274|US Guidance for fine needle aspiration of Breast - right
C1526274|Brst-R US FNA Asp
C1526274|Guidance for aspiration.fine needle:Find:Pt:Breast.right:Doc:US
C1526274|Guidance for aspiration.fine needle:Finding:Point in time:Breast.right:Document:Ultrasound
C1526281|Femur-R US
C1526281|Femur - right US
C1526281|Multisection:Finding:Point in time:Femur.right:Document:Ultrasound
C1526281|Multisection:Find:Pt:Femur.right:Doc:US
C1508081|Multisection sagittal:Find:Pt:Spine.lumbosacral+Cervical+Thoracic:Doc:MRI
C1508081|Multisection sagittal:Finding:Point in time:Spine.lumbosacral+Cervical+Thoracic:Document:MRI
C1508081|Deprecated Spine.lumbosacral+Cervical+Thoracic MRI sagittal
C1508081|Deprecated Lumbrosac+C+T-spine MRI Sagit
C1525912|Spine US CSF asp guid
C1525912|US Guidance for CSF aspiration of Spine
C1525912|Guidance for CSF aspiration:Find:Pt:Spine:Doc:US
C1525912|Guidance for CSF aspiration:Finding:Point in time:Spine:Document:Ultrasound
C1508085|Knee-L XR Sunrise 20+40+60 Deg
C1508085|Knee - left X-ray Sunrise 20 and 40 and 60 degrees
C1508085|Views Sunrise 20 & 40 & 60 degrees:Finding:Point in time:Knee.left:Document:XR
C1508085|Views Sunrise 20 & 40 & 60 degrees:Find:Pt:Knee.left:Doc:XR
C1524477|Deprecated Head.cistern CT W contr IT
C1524477|Multisection^W contrast IT:Find:Pt:Head.cistern:Nar:CT
C1524477|Deprecated Head Cistern CT Multisection W contrast IT
C1524477|Multisection^W contrast Intrathecal:Finding:Point in time:Head.cistern:Narrative:Computerized Tomography
C1524495|Brst-L MRI W contr IV
C1524495|Breast - left MRI W contrast IV
C1524495|Multisection^W contrast Intravenous:Finding:Point in time:Breast.left:Document:MRI
C1524495|Multisection^W contrast IV:Find:Pt:Breast.left:Doc:MRI
C1524507|LE-Bl MRI W contr IV
C1524507|Lower extremity - bilateral MRI W contrast IV
C1524507|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.bilateral:Document:MRI
C1524507|Multisection^W contrast IV:Find:Pt:Lower extremity.bilateral:Doc:MRI
C1524509|LE-L MRI W contr IV
C1524509|Lower extremity - left MRI W contrast IV
C1524509|Multisection^W contrast IV:Find:Pt:Lower extremity.left:Doc:MRI
C1524509|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.left:Document:MRI
C1524882|LE.joint MRI WO contr
C1524882|Lower Extremity Joint MRI WO contrast
C1524882|Multisection^WO contrast:Find:Pt:Lower extremity.joint:Doc:MRI
C1524882|Multisection^WO contrast:Finding:Point in time:Lower extremity.joint:Document:MRI
C1524901|Thoracic outlet - right MRI WO contrast
C1524901|TO-R MRI WO contr
C1524901|Multisection^WO contrast:Find:Pt:Thoracic outlet.right:Doc:MRI
C1524901|Multisection^WO contrast:Finding:Point in time:Thoracic outlet.right:Document:MRI
C1524923|Chest ves MRI.Angio WO contr
C1524923|Chest vessels MRI angiogram WO contrast
C1524923|Multisection^WO contrast:Finding:Point in time:Chest vessels:Document:MRI.angio
C1524923|Multisection^WO contrast:Find:Pt:Chest vessels:Doc:MRI.angio
C1524556|Knee CT W contr IV
C1524556|Knee CT W contrast IV
C1524556|Multisection^W contrast IV:Find:Pt:Knee:Doc:CT
C1524556|Multisection^W contrast Intravenous:Finding:Point in time:Knee:Document:Computerized Tomography
C1524557|Knee MRI W contr IV
C1524557|Knee MRI W contrast IV
C1524557|Multisection^W contrast Intravenous:Finding:Point in time:Knee:Document:MRI
C1524557|Multisection^W contrast IV:Find:Pt:Knee:Doc:MRI
C1524202|Chest XR AP 1V
C1524202|Chest X-ray AP single view
C1524202|View AP:Find:Pt:Chest:Doc:XR
C1524202|View AP:Finding:Point in time:Chest:Document:XR
C1524210|Ft-Bl XR AP 1V
C1524210|Foot - bilateral X-ray AP single view
C1524210|View AP:Find:Pt:Foot.bilateral:Doc:XR
C1524210|View AP:Finding:Point in time:Foot.bilateral:Document:XR
C1524607|Aorta abdominal MRI WO and W contrast IV
C1524607|Ab Ao MRI WO+W contr IV
C1524607|Multisection^WO & W contrast Intravenous:Finding:Point in time:Aorta.abdominal:Document:MRI
C1524607|Multisection^WO & W contrast IV:Find:Pt:Aorta.abdominal:Doc:MRI
C1524956|Elbow X-ray oblique
C1524956|Elbow XR Obl
C1524956|Views oblique:Finding:Point in time:Elbow:Document:XR
C1524956|Views oblique:Find:Pt:Elbow:Doc:XR
C1524965|Hip XR Obl 1V
C1524965|Hip X-ray oblique single view
C1524965|View oblique:Finding:Point in time:Hip:Document:XR
C1524965|View oblique:Find:Pt:Hip:Doc:XR
C1524982|Sacroiliac joint - left X-ray
C1524982|SIJ-L XR
C1524982|Views:Finding:Point in time:Sacroiliac joint.left:Document:XR
C1524982|Views:Find:Pt:Sacroiliac joint.left:Doc:XR
C1524983|Knee - bilateral X-ray
C1524983|Knee-Bl XR
C1524983|Views:Finding:Point in time:Knee.bilateral:Document:XR
C1524983|Views:Find:Pt:Knee.bilateral:Doc:XR
C1524986|Patella-Bl XR
C1524986|Patella - bilateral X-ray
C1524986|Views:Finding:Point in time:Patella.bilateral:Document:XR
C1524986|Views:Find:Pt:Patella.bilateral:Doc:XR
C1524656|Shoulder - left X-ray 4 views
C1524656|Should-L XR 4V
C1524656|Views 4:Find:Pt:Shoulder.left:Doc:XR
C1524656|Views 4:Finding:Point in time:Shoulder.left:Document:XR
C1525002|Femur-L XR 2V
C1525002|Femur - left X-ray 2 views
C1525002|Views 2:Find:Pt:Femur.left:Doc:XR
C1525002|Views 2:Finding:Point in time:Femur.left:Document:XR
C1525014|Face XR 5V
C1525014|Facial bones X-ray 5 views
C1525014|Views 5:Find:Pt:Facial bones:Doc:XR
C1525014|Views 5:Finding:Point in time:Facial bones:Document:XR
C1525022|Wrist - left X-ray 8 views
C1525022|Wrist-L XR 8V
C1525022|Views 8:Finding:Point in time:Wrist.left:Document:XR
C1525022|Views 8:Find:Pt:Wrist.left:Doc:XR
C1524383|Femur - right CT
C1524383|Femur-R CT
C1524383|Multisection:Find:Pt:Femur.right:Doc:CT
C1524383|Multisection:Finding:Point in time:Femur.right:Document:Computerized Tomography
C1525028|Elbow XR AP+Lat
C1525028|Elbow X-ray AP and lateral
C1525028|Views AP & lateral:Find:Pt:Elbow:Doc:XR
C1525028|Views AP & lateral:Finding:Point in time:Elbow:Document:XR
C1527041|Kidney MRI
C1527041|Multisection:Finding:Point in time:Kidney:Narrative:MRI
C1527041|Multisection:Find:Pt:Kidney:Doc:MRI
C1527041|Multisection:Finding:Point in time:Kidney:Document:MRI
C1524669|Deprecated Heel XR AP+Lat+Obl
C1524669|Views AP & lateral & oblique:Find:Pt:Calcaneus:Doc:XR
C1524669|Views AP & lateral & oblique:Finding:Point in time:Calcaneus:Document:XR
C1524669|Deprecated Calcaneus X-ray AP and lateral and oblique
C1830201|Multisection coronal:Find:Pt:Sinuses:Doc:CT
C1830201|Multisection coronal:Finding:Point in time:Sinuses:Document:Computerized Tomography
C1830201|Deprecated Sinuses CT coronal
C1830224|Brst-UL MRI W contr IV
C1830224|Breast - unilateral MRI W contrast IV
C1830224|Multisection^W contrast IV:Find:Pt:Breast.unilateral:Doc:MRI
C1830224|Multisection^W contrast Intravenous:Finding:Point in time:Breast.unilateral:Document:MRI
C1830270|Elbow+Radius+Ulna XR
C1830270|Elbow+Radius+Ulna X-ray
C1830270|Views:Find:Pt:Elbow+Radius+Ulna:Doc:XR
C1830270|Views:Finding:Point in time:Elbow+Radius+Ulna:Document:XR
C1715440|Neck vessels US.doppler
C1715440|Neck ves DOP
C1715440|Multisection:Finding:Point in time:Neck vessels:Document:Ultrasound.doppler
C1715440|Multisection:Find:Pt:Neck vessels:Doc:US.doppler
C1715447|Hand XR 2V port
C1715447|Hand X-ray 2 views portable
C1715447|Views 2 portable:Find:Pt:Hand:Doc:XR
C1715447|Views 2 portable:Finding:Point in time:Hand:Document:XR
C1715448|Radius+Ulna XR 2V port
C1715448|Radius and Ulna X-ray 2 views portable
C1715448|Views 2 portable:Find:Pt:Radius+Ulna:Doc:XR
C1715448|Views 2 portable:Finding:Point in time:Radius+Ulna:Document:XR
C1717321|Fluoroscopy Guidance for fine needle aspiration of Thyroid
C1717321|Thyroid Flr FNA Asp
C1717321|Guidance for aspiration.fine needle:Find:Pt:Thyroid:Doc:XR.fluor
C1717321|Guidance for aspiration.fine needle:Finding:Point in time:Thyroid:Document:XR.fluor
C1715480|Liver Flr FNA Asp
C1715480|Fluoroscopy Guidance for fine needle aspiration of Liver
C1715480|Guidance for aspiration.fine needle:Find:Pt:Liver:Doc:XR.fluor
C1715480|Guidance for aspiration.fine needle:Finding:Point in time:Liver:Document:XR.fluor
C1649481|Shoulder - left X-ray portable
C1649481|Should-L XR port
C1649481|Views portable:Find:Pt:Shoulder.left:Doc:XR
C1649481|Views portable:Finding:Point in time:Shoulder.left:Document:XR
C1649484|Hand - left X-ray portable
C1649484|Hand-L XR port
C1649484|Views portable:Finding:Point in time:Hand.left:Document:XR
C1649484|Views portable:Find:Pt:Hand.left:Doc:XR
C1632789|IMAl-L Flr Inj guid
C1632789|Fluoroscopy Guidance for injection of Mammary artery.internal - left
C1632789|Guidance for injection:Find:Pt:Mammary artery.internal.left:Doc:XR.fluor
C1632789|Guidance for injection:Finding:Point in time:Mammary artery.internal.left:Document:XR.fluor
C1717258|Views survey:Finding:Point in time:To be specified in another part of the message bones:Narrative:XR
C1717258|Bones X-ray survey
C1717258|Bones XR Survey
C1717258|Views survey:Find:Pt:Bones:Doc:XR
C1717258|Views survey:Finding:Point in time:Bones:Document:XR
C1714924|Unspecified body region CT WO contrast
C1714924|XXX CT WO contr
C1714924|Multisection^WO contrast:Find:Pt:XXX:Doc:CT
C1714924|Multisection^WO contrast:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1714929|Orbit+Face+Neck MRI
C1714929|Orbit and Face and Neck MRI
C1714929|Multisection:Find:Pt:Orbit+Face+Neck:Doc:MRI
C1714929|Multisection:Finding:Point in time:Orbit+Face+Neck:Document:MRI
C1714939|Brain RI Static+Flow W RNC IV
C1714939|Brain Scan static and flow
C1714939|Views static & flow^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc
C1714939|Views static & flow^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1714499|Renal ves RI Flow W Tc99mMAG3 IV
C1714499|Renal vessels Scan flow W Tc-99m Mertiatide IV
C1714499|Views flow^W Tc-99m Mertiatide Intravenous:Finding:Point in time:Renal vessels:Document:Radnuc
C1714499|Views flow^W Tc-99m Mertiatide IV:Find:Pt:Renal vessels:Doc:Radnuc
C1714501|KD-Bl+Renal ves RI W Tc99mDTPA IV
C1714501|Views^W Tc-99m DTPA IV:Find:Pt:Kidney.bilateral+Renal vessels:Doc:Radnuc
C1714501|Views^W Tc-99m DTPA Intravenous:Finding:Point in time:Kidney.bilateral+Renal vessels:Document:Radnuc
C1714501|Kidney - bilateral and Renal vessels Scan W Tc-99m DTPA IV
C1715091|Vein XRA Thrombect guid W contr IV
C1715091|Fluoroscopic angiogram Guidance for thrombectomy of Vein-- W contrast IV
C1715091|Guidance for thrombectomy^W contrast Intravenous:Finding:Point in time:Vein:Document:XR.fluor.angio
C1715091|Guidance for thrombectomy^W contrast IV:Find:Pt:Vein:Doc:XR.fluor.angio
C1715105|Knee - left X-ray Sunrise
C1715105|Knee-L XR Sunrise
C1715105|View Sunrise:Find:Pt:Knee.left:Doc:XR
C1715105|View Sunrise:Finding:Point in time:Knee.left:Document:XR
C1715121|Tibioperoneal arteries - left Fluoroscopic angiogram Angioplasty W contrast IA
C1715121|Tibioperon aa-L XRA Angpsty W contr IA
C1715121|Angioplasty^W contrast IA:Find:Pt:Tibioperoneal arteries.left:Doc:XR.fluor.angio
C1715121|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibioperoneal arteries.left:Document:XR.fluor.angio
C1636075|Lower extremity vessel graft - left US.doppler
C1636075|LE ves graft-L DOP
C1636075|Multisection:Finding:Point in time:Lower extremity vessel graft.left:Document:Ultrasound.doppler
C1636075|Multisection:Find:Pt:Lower extremity vessel graft.left:Doc:US.doppler
C1626177|Breast - bilateral FFD mammogram screening
C1626177|Views screening:Finding:Point in time:Breast.bilateral:Document:Mam.FFD
C1626177|Views screening:Find:Pt:Breast.bilateral:Doc:Mam.FFD
C1626177|Brst-Bl FFDM Screening
C1642593|Deprecated Views:Finding:Point in time:Tibia.right:Narrative:XR
C1642593|Views:Find:Pt:Tibia.right:Nar:XR
C1642593|Deprecated Tib-R XR
C1642593|Views:Finding:Point in time:Tibia.right:Narrative:XR
C1642593|Deprecated Tibia Right X-ray
C1632224|Retroperitoneum CT WO contr
C1632224|Retroperitoneum CT WO contrast
C1632224|Multisection^WO contrast:Find:Pt:Abdomen>Retroperitoneum:Doc:CT
C1632224|Multisection^WO contrast:Finding:Point in time:Abdomen>Retroperitoneum:Document:Computerized Tomography
C1632956|Hrt RI Rest+stress+W Tl201 IV
C1632956|Heart Scan at rest and W stress and W Tl-201 IV
C1632956|Views^at rest & W stress & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1632956|Views^at rest & W stress & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1632231|Ribs-L XR 1V
C1632231|Ribs - left X-ray Single view
C1632231|View 1:Finding:Point in time:Ribs.left:Document:XR
C1632231|View 1:Find:Pt:Ribs.left:Doc:XR
C1641064|C-spine XR 6V
C1641064|Views 6:Find:Pt:Spine.cervical:Doc:XR
C1641064|Views 6:Finding:Point in time:Spine.cervical:Document:XR
C1641064|Cervical spine X-ray 6 views
C1954374|Deprecated Mandible - left X-ray
C1954374|Views:Finding:Point in time:Mandible.left:Document:XR
C1954374|Views:Find:Pt:Mandible.left:Doc:XR
C1954374|Deprecated Mandible-L XR
C1954376|Orbit - bilateral X-ray GE 4 views
C1954376|Orbit-Bl XR GE 4V
C1954376|Views GE 4:Find:Pt:Orbit.bilateral:Doc:XR
C1954376|Views GE 4:Finding:Point in time:Orbit.bilateral:Document:XR
C1953324|Mastoid - bilateral X-ray 1 or 2 views
C1953324|Mastoid-Bl XR 1V or 2V
C1953324|Views 1 or 2:Finding:Point in time:Mastoid.bilateral:Document:XR
C1953324|Views 1 or 2:Find:Pt:Mastoid.bilateral:Doc:XR
C1953950|Brain.temporal MRI W contr IV
C1953950|Brain.temporal MRI W contrast IV
C1953950|Multisection^W contrast IV:Find:Pt:Brain.temporal:Doc:MRI
C1953950|Multisection^W contrast Intravenous:Finding:Point in time:Brain.temporal:Document:MRI
C1953979|T-spine XR 3V+Swimmers
C1953979|Views 3 & Swimmers:Finding:Point in time:Spine.thoracic:Document:XR
C1953979|Views 3 & Swimmers:Find:Pt:Spine.thoracic:Doc:XR
C1953979|Thoracic spine X-ray 3 views and Swimmers
C1952655|Mastoid - left X-ray 1 or 2 views
C1952655|Mastoid-L XR 1V or 2V
C1952655|Views 1 or 2:Find:Pt:Mastoid.left:Doc:XR
C1952655|Views 1 or 2:Finding:Point in time:Mastoid.left:Document:XR
C2925710|CT Guidance for ablation of tissue of Unspecified body region
C2925710|XXX CT Ablation guid
C2925710|Guidance for ablation of tissue:Find:Pt:XXX:Doc:CT
C2925710|Guidance for ablation of tissue:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C3533556|Fluoroscopy Guidance for removal of CVA lumen obstruction from Central vein
C3533556|Guidance for removal of CVA lumen obstruction:Find:Pt:Central vein:Doc:XR.fluor
C3533556|Centl v Flr CVA lumen obs rem guid
C3533556|Guidance for removal of CVA lumen obstruction:Finding:Point in time:Central vein:Document:XR.fluor
C3533478|US Guidance for injection of sclerosing agent of Extremity vein - left
C3533478|Guidance for injection of sclerosing agent:Find:Pt:Extremity vein.left:Doc:US
C3533478|Guidance for injection of sclerosing agent:Finding:Point in time:Extremity vein.left:Document:Ultrasound
C3533478|Extr v-L US Sclerosing agent inj guid
C3262932|Ankle-R CT W contr IS
C3262932|Multisection^W contrast IS:Find:Pt:Ankle.right:Doc:CT
C3262932|Ankle - right CT W contrast IS
C3262932|Multisection^W contrast Intrasynovial:Finding:Point in time:Ankle.right:Document:Computerized Tomography
C3262975|Should-L XR Grashey & Y
C3262975|Shoulder - left X-ray Grashey and Y
C3262975|Views Grashey & Y:Find:Pt:Shoulder.left:Doc:XR
C3262975|Views Grashey & Y:Finding:Point in time:Shoulder.left:Document:XR
C3483134|L-spine US CSF asp guid
C3483134|Guidance for CSF aspiration:Find:Pt:Spine.lumbar:Doc:US
C3483134|Guidance for CSF aspiration:Finding:Point in time:Spine.lumbar:Document:Ultrasound
C3483134|US Guidance for CSF aspiration of Lumbar spine
C3263057|Fluoroscopy Guidance for percutaneous drainage of abscess of Pelvis
C3263057|Pelvis Flr PC Abscess Drain guid
C3263057|Guidance for percutaneous drainage of abscess:Finding:Point in time:Pelvis:Document:XR.fluor
C3263057|Guidance for percutaneous drainage of abscess:Find:Pt:Pelvis:Doc:XR.fluor
C3261714|LN US Bx CN guid
C3261714|US Guidance for core needle biopsy of Lymph node
C3261714|Guidance for biopsy.core needle:Find:Pt:Lymph node:Doc:US
C3261714|Guidance for biopsy.core needle:Finding:Point in time:Lymph node:Document:Ultrasound
C3263205|Femoral artery and Popliteal artery US
C3263205|Fem a+Popliteal a US
C3263205|Multisection:Find:Pt:Femoral artery+Popliteal artery:Doc:US
C3263205|Multisection:Finding:Point in time:Femoral artery+Popliteal artery:Document:Ultrasound
C3262895|Wrist-Bl XR Ulnar+Radial Deviation
C3262895|Wrist - bilateral X-ray ulnar deviation and radial deviation
C3262895|Views ulnar deviation & radial deviation:Find:Pt:Wrist.bilateral:Doc:XR
C3262895|Views ulnar deviation & radial deviation:Finding:Point in time:Wrist.bilateral:Document:XR
C3262917|CT Guidance for biopsy of Pelvis-- WO contrast
C3262917|Pelvis CT Bx guid WO contr
C3262917|Guidance for biopsy^WO contrast:Finding:Point in time:Pelvis:Document:Computerized Tomography
C3262917|Guidance for biopsy^WO contrast:Find:Pt:Pelvis:Doc:CT
C0944156|Views:Finding:Point in time:Knee:Narrative:XR
C0944156|Knee X-ray
C0944156|Knee XR
C0944156|Views:Finding:Point in time:Knee:Document:XR
C0944156|Views:Find:Pt:Knee:Doc:XR
C0942154|Optic foramen - bilateral X-ray
C0942154|Optic foramen-Bl XR
C0942154|Views:Find:Pt:Optic foramen.bilateral:Doc:XR
C0942154|Views:Finding:Point in time:Optic foramen.bilateral:Document:XR
C0945316|Ribs - bilateral X-ray
C0945316|Ribs-Bl XR
C0945316|Views:Find:Pt:Ribs.bilateral:Doc:XR
C0945316|Views:Finding:Point in time:Ribs.bilateral:Document:XR
C0942312|US Guidance for drainage of Extremity - bilateral
C0942312|Extr-Bl US Drain guid
C0942312|Guidance for drainage:Find:Pt:Extremity.bilateral:Doc:US
C0942312|Guidance for drainage:Finding:Point in time:Extremity.bilateral:Document:Ultrasound
C0942333|Brst-L Mam Dx Ltd
C0942333|Breast - left Mammogram diagnostic limited
C0942333|Views diagnostic limited:Find:Pt:Breast.left:Doc:Mam
C0942333|Views diagnostic limited:Finding:Point in time:Breast.left:Document:Mam
C0942341|Knee-Bl XR AP+PA stand
C0942341|Knee - bilateral X-ray AP and PA standing
C0942341|Views AP & PA^standing:Find:Pt:Knee.bilateral:Doc:XR
C0942341|Views AP & PA^standing:Finding:Point in time:Knee.bilateral:Document:XR
C0942371|Knee-Bl XR 2V
C0942371|Knee - bilateral X-ray 2 views
C0942371|Views 2:Find:Pt:Knee.bilateral:Doc:XR
C0942371|Views 2:Finding:Point in time:Knee.bilateral:Document:XR
C0882017|Lower leg ves MRI.Angio W contr IV
C0882017|Lower leg vessels MRI angiogram W contrast IV
C0882017|Multisection^W contrast IV:Find:Pt:Lower leg vessels:Doc:MRI.angio
C0882017|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg vessels:Document:MRI.angio
C0882024|Views:Finding:Point in time:Mandible:Narrative:XR
C0882024|Mandible XR
C0882024|Mandible X-ray
C0882024|Views:Finding:Point in time:Mandible:Document:XR
C0882024|Views:Find:Pt:Mandible:Doc:XR
C0882080|Rect+Bladder Flr W contr PR+IB def+void
C0882080|Rectum and Urinary bladder Fluoroscopy W contrast PR and intra bladder during defecation and voiding
C0882080|Views^W contrast PR & intra bladder during defecation & voiding:Find:Pt:Rectum+Urinary bladder:Doc:XR.fluor
C0882080|Views^W contrast Rectal & intra bladder during defecation & voiding:Finding:Point in time:Rectum+Urinary bladder:Document:XR.fluor
C0882155|Fluoroscopy Guidance for placement of tube in Stomach
C0882155|Stom Flr Tube plac guid
C0882155|Guidance for placement of tube:Find:Pt:Stomach:Doc:XR.fluor
C0882155|Guidance for placement of tube:Finding:Point in time:Stomach:Document:XR.fluor
C0882188|Bone RI W In-111 WBC IV
C0882188|Bone Scan W In-111 tagged WBC IV
C0882188|Views^W In-111 tagged WBC IV:Find:Pt:Bone:Doc:Radnuc
C0882188|Views^W In-111 tagged WBC Intravenous:Finding:Point in time:Bone:Document:Radnuc
C0882195|XXX CT Ltd
C0882195|Unspecified body region CT limited
C0882195|Multisection limited:Find:Pt:XXX:Doc:CT
C0882195|Multisection limited:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0942091|Salivary gland - left Fluoroscopy W contrast intra salivary duct
C0942091|Salivary gland-L Flr W contr intra SD
C0942091|Views^W contrast intra salivary duct:Finding:Point in time:Salivary gland.left:Document:XR.fluor
C0942091|Views^W contrast intra salivary duct:Find:Pt:Salivary gland.left:Doc:XR.fluor
C0882517|TA CT W contr IV
C0882517|Multisection^W contrast Intravenous:Finding:Point in time:Chest>Aorta.thoracic:Document:Computerized Tomography
C0882517|Multisection^W contrast IV:Find:Pt:Chest>Aorta.thoracic:Doc:CT
C0882517|Thoracic Aorta CT W contrast IV
C0881799|Abd XR AP L-Lat Decub Port
C0881799|Abdomen X-ray AP left lateral-decubitus portable
C0881799|View AP L-lateral-decubitus portable:Finding:Point in time:Abdomen:Document:XR
C0881799|View AP L-lateral-decubitus portable:Find:Pt:Abdomen:Doc:XR
C0882518|BDs+GB RI for Bil Pat+EF W Sinc+RNC IV
C0882518|Biliary ducts and Gallbladder Scan for patency of biliary structures and ejection fraction W sincalide and W radionuclide IV
C0882518|Views for patency of biliary structures & ejection fraction^W sincalide & W radionuclide Intravenous:Finding:Point in time:Biliary ducts+Gallbladder:Document:Radnuc
C0882518|Views for patency of biliary structures & ejection fraction^W sincalide & W radionuclide IV:Find:Pt:Biliary ducts+Gallbladder:Doc:Radnuc
C0881855|Centl v XRA CC change guid W contr IV
C0881855|Fluoroscopic angiogram Guidance for change of central catheter in Central vein-- W contrast IV
C0881855|Guidance for change of central catheter^W contrast Intravenous:Finding:Point in time:Central vein:Document:XR.fluor.angio
C0881855|Guidance for change of central catheter^W contrast IV:Find:Pt:Central vein:Doc:XR.fluor.angio
C0881868|Chest XR L-Lat Upr
C0881868|Chest X-ray left lateral upright
C0881868|View L-lateral upright:Finding:Point in time:Chest:Document:XR
C0881868|View L-lateral upright:Find:Pt:Chest:Doc:XR
C0881904|Esophagus Fluoroscopy W gastrografin PO
C0881904|Esoph Flr W Gastrografin PO
C0881904|Views^W gastrografin Oral:Finding:Point in time:Esophagus:Document:XR.fluor
C0881904|Views^W gastrografin PO:Find:Pt:Esophagus:Doc:XR.fluor
C0884111|Views:Finding:Point in time:Facial bones:Narrative:XR
C0884111|Facial bones X-ray
C0884111|Face XR
C0884111|Views:Find:Pt:Facial bones:Doc:XR
C0884111|Views:Finding:Point in time:Facial bones:Document:XR
C0881918|Facial bones CT
C0881918|Multisection:Finding:Point in time:Facial bones:Document:Computerized Tomography
C0881918|Multisection:Find:Pt:Facial bones:Doc:CT
C0881918|Face CT
C0881944|Multisection^WO & W contrast IV:Find:Pt:Head:Doc:CT
C0881944|Head CT WO+W contr IV
C0881944|Head CT WO and W contrast IV
C0881944|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head:Document:Computerized Tomography
C0881965|Hip US
C0881965|Multisection:Find:Pt:Hip:Doc:US
C0881965|Multisection:Finding:Point in time:Hip:Document:Ultrasound
C1114936|US Guidance for aspiration of cyst of Unspecified body region
C1114936|XXX US Cyst Asp guid
C1114936|Guidance for aspiration of cyst:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1114936|Guidance for aspiration of cyst:Find:Pt:XXX:Doc:US
C1114937|Liver US during surgery
C1114937|Liver US in Surg
C1114937|Multisection^during surgery:Find:Pt:Liver:Doc:US
C1114937|Multisection^during surgery:Finding:Point in time:Liver:Document:Ultrasound
C1114523|LE US
C1114523|Lower extremity US
C1114523|Multisection:Finding:Point in time:Lower extremity:Document:Ultrasound
C1114523|Multisection:Find:Pt:Lower extremity:Doc:US
C1114563|T-spine XR AP 1V
C1114563|View AP:Find:Pt:Spine.thoracic:Doc:XR
C1114563|View AP:Finding:Point in time:Spine.thoracic:Document:XR
C1114563|Thoracic spine X-ray AP single view
C1114571|Abd XR AP+Lat Xtable port
C1114571|Abdomen X-ray AP and lateral crosstable portable
C1114571|Views AP & lateral crosstable portable:Find:Pt:Abdomen:Doc:XR
C1114571|Views AP & lateral crosstable portable:Finding:Point in time:Abdomen:Document:XR
C1114668|Forearm vessels MRI angiogram
C1114668|Forearm ves MRI.Angio
C1114668|Multisection:Find:Pt:Forearm vessels:Doc:MRI.angio
C1114668|Multisection:Finding:Point in time:Forearm vessels:Document:MRI.angio
C1114415|IAC CT WO contr
C1114415|Internal auditory canal CT WO contrast
C1114415|Multisection^WO contrast:Finding:Point in time:Internal auditory canal:Document:Computerized Tomography
C1114415|Multisection^WO contrast:Find:Pt:Internal auditory canal:Doc:CT
C1114424|CT Guidance for fine needle aspiration of Lung
C1114424|Lung CT FNA Asp
C1114424|Guidance for aspiration.fine needle:Find:Pt:Chest>Lung:Doc:CT
C1114424|Guidance for aspiration.fine needle:Finding:Point in time:Chest>Lung:Document:Computerized Tomography
C1114430|CT Guidance for fine needle aspiration of Abdomen
C1114430|Abd CT FNA Asp
C1114430|Guidance for aspiration.fine needle:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1114430|Guidance for aspiration.fine needle:Find:Pt:Abdomen:Doc:CT
C1114446|Multisection^W & WO contrast Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:Computerized Tomography
C1114446|Deprecated Kidney - bilateral and Collecting system CT W and WO contrast IV
C1114446|Multisection^W & WO contrast IV:Find:Pt:Kidney.bilateral+Collecting system:Nar:CT
C1114446|Deprecated KD-Bl+CS CT W+WO contr IV
C1114926|Fluoroscopy Guidance for removal of foreign body from Unspecified body region
C1114926|XXX Flr FB rem guid
C1114926|Guidance for removal of foreign body:Find:Pt:XXX:Doc:XR.fluor
C1114926|Guidance for removal of foreign body:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1543451|T+L-spine XR Scoli AP+Lat stand
C1543451|Spine Thoracic and Lumbar X-ray scoliosis AP and lateral standing
C1543451|Views scoliosis AP & lateral^standing:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1543451|Views scoliosis AP & lateral^standing:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1543739|RI for Lymphoma W Ga-67 IV
C1543739|Views for lymphoma^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543739|Views for lymphoma^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543739|Scan for lymphoma W Ga-67 IV
C1543759|Hrt RI PF W DPY+Tl-201 IV
C1543759|Heart Scan perfusion W dipyridamole and W Tl-201 IV
C1543759|Views perfusion^W dipyridamole & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1543759|Views perfusion^W dipyridamole & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543473|Should-R XR AP(w IR+ER)
C1543473|Shoulder - right X-ray AP (W internal rotation and W external rotation)
C1543473|Views AP (W internal rotation & W external rotation):Find:Pt:Shoulder.right:Doc:XR
C1543473|Views AP (W internal rotation & W external rotation):Finding:Point in time:Shoulder.right:Document:XR
C1543795|Prostate SPECT W Tc99mPMSA IV
C1543795|Prostate SPECT W Tc-99m capromab pendatide IV
C1543795|Multisection^W Tc-99m capromab pendatide Intravenous:Finding:Point in time:Prostate:Document:Radnuc.SPECT
C1543795|Multisection^W Tc-99m capromab pendatide IV:Find:Pt:Prostate:Doc:Radnuc.SPECT
C1543859|Bone Scan static whole body
C1543859|Bone RI Static WB W RNC IV
C1543859|Views static whole body ^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543859|Views static whole body^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543888|Bone RI Flow W RNC IV
C1543888|Bone Scan flow
C1543888|Views flow^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543888|Views flow^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543925|Bone RI Static Mul Areas W RNC IV
C1543925|Bone Scan static multiple areas
C1543925|Views static multiple areas^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543925|Views static multiple areas^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543939|Hrt RI Gated+EF W RNC IV
C1543939|Heart Scan gated and ejection fraction
C1543939|Views gated & ejection fraction^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543939|Views gated & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543515|Extr a-R DOP
C1543515|Extremity artery - right US.doppler
C1543515|Multisection:Find:Pt:Extremity artery.right:Doc:US.doppler
C1543515|Multisection:Finding:Point in time:Extremity artery.right:Document:Ultrasound.doppler
C1543516|Extremity vein - right US.doppler
C1543516|Extr v-R DOP
C1543516|Multisection:Finding:Point in time:Extremity vein.right:Document:Ultrasound.doppler
C1543516|Multisection:Find:Pt:Extremity vein.right:Doc:US.doppler
C1543157|Vein US
C1543157|Multisection:Find:Pt:Vein:Doc:US
C1543157|Multisection:Finding:Point in time:Vein:Document:Ultrasound
C1543574|Fem ves-L DOP
C1543574|Femoral vessels - left US.doppler
C1543574|Multisection:Find:Pt:Femoral vessels.left:Doc:US.doppler
C1543574|Multisection:Finding:Point in time:Femoral vessels.left:Document:Ultrasound.doppler
C1543167|Pelvis CT Ltd Pelvimetry WO contr
C1543167|Multisection limited for pelvimetry^WO contrast:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1543167|Multisection limited for pelvimetry^WO contrast:Find:Pt:Pelvis:Doc:CT
C1543167|Pelvis CT limited for pelvimetry WO contrast
C1543172|Chest XR Lat
C1543172|Chest X-ray lateral
C1543172|View lateral:Finding:Point in time:Chest:Document:XR
C1543172|View lateral:Find:Pt:Chest:Doc:XR
C1543188|C+T+L-spine XR AP+Lat
C1543188|Spine Cervical and Thoracic and Lumbar X-ray AP and lateral
C1543188|Views AP & lateral:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:XR
C1543188|Views AP & lateral:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:XR
C1543197|Ft XR AP+Obl
C1543197|Foot X-ray AP and oblique
C1543197|Views AP & oblique:Finding:Point in time:Foot:Document:XR
C1543197|Views AP & oblique:Find:Pt:Foot:Doc:XR
C1526763|Brst-R Mam Spot
C1526763|Breast - right Mammogram spot
C1526763|Views spot:Finding:Point in time:Breast.right:Document:Mam
C1526763|Views spot:Find:Pt:Breast.right:Doc:Mam
C1543704|Brain RI W Tc99mGHA IV
C1543704|Brain Scan W Tc-99m glucoheptonate IV
C1543704|Views^W Tc-99m glucoheptonate IV:Find:Pt:Brain:Doc:Radnuc
C1543704|Views^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1543733|SPECT WB W Ga-67 IV
C1543733|Multisection whole body^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543733|Multisection whole body^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1543733|SPECT whole body W Ga-67 IV
C1543414|Should-Bl XR AP(w IR+ER)
C1543414|Shoulder - bilateral X-ray AP (W internal rotation and W external rotation)
C1543414|Views AP (W internal rotation & W external rotation):Find:Pt:Shoulder.bilateral:Doc:XR
C1543414|Views AP (W internal rotation & W external rotation):Finding:Point in time:Shoulder.bilateral:Document:XR
C1525114|Neck veins MRI angiogram
C1525114|Neck vv MRI.Angio
C1525114|Multisection:Find:Pt:Neck veins:Doc:MRI.angio
C1525114|Multisection:Finding:Point in time:Neck veins:Document:MRI.angio
C1525174|Upper extremity vessels - right MRI angiogram
C1525174|UE ves-R MRI.Angio
C1525174|Multisection:Finding:Point in time:Upper extremity vessels.right:Document:MRI.angio
C1525174|Multisection:Find:Pt:Upper extremity vessels.right:Doc:MRI.angio
C1524447|Hip CT Ltd
C1524447|Hip CT limited
C1524447|Multisection limited:Find:Pt:Hip:Doc:CT
C1524447|Multisection limited:Finding:Point in time:Hip:Document:Computerized Tomography
C1524463|Multisection^W contrast IS:Find:Pt:Elbow.right:Doc:MRI
C1524463|Multisection^W contrast Intrasynovial:Finding:Point in time:Elbow.right:Document:MRI
C1524463|Elbow - right MRI W contrast IS
C1524463|Elbow-R MRI W contr IS
C1525284|Abd+Pelvis CT WO contr
C1525284|Abdomen and Pelvis CT WO contrast
C1525284|Multisection^WO contrast:Find:Pt:Abdomen+Pelvis:Doc:CT
C1525284|Multisection^WO contrast:Finding:Point in time:Abdomen+Pelvis:Document:Computerized Tomography
C1525294|Brst Mam Ax
C1525294|Breast Mammogram axillary
C1525294|View axillary:Find:Pt:Breast:Doc:Mam
C1525294|View axillary:Finding:Point in time:Breast:Document:Mam
C1525317|Hip XR Lat Xtable
C1525317|Hip X-ray lateral crosstable
C1525317|View lateral crosstable:Finding:Point in time:Hip:Document:XR
C1525317|View lateral crosstable:Find:Pt:Hip:Doc:XR
C1525202|Neck vv MRI.Angio W contr IV
C1525202|Neck veins MRI angiogram W contrast IV
C1525202|Multisection^W contrast Intravenous:Finding:Point in time:Neck veins:Document:MRI.angio
C1525202|Multisection^W contrast IV:Find:Pt:Neck veins:Doc:MRI.angio
C1524224|Hip X-ray Von rossen
C1524224|Hip XR Von Rossen
C1524224|View Von rossen:Find:Pt:Hip:Doc:XR
C1524224|View Von rossen:Finding:Point in time:Hip:Document:XR
C1525472|Hip - bilateral X-ray standing
C1525472|Hip-Bl XR stand
C1525472|View^standing:Find:Pt:Hip.bilateral:Doc:XR
C1525472|View^standing:Finding:Point in time:Hip.bilateral:Document:XR
C1525503|Hip-Bl XR AP+Lat Frog
C1525503|Hip - bilateral X-ray AP and lateral frog
C1525503|Views AP & lateral frog:Find:Pt:Hip.bilateral:Doc:XR
C1525503|Views AP & lateral frog:Finding:Point in time:Hip.bilateral:Document:XR
C1525506|Ankle XR AP+Lat+Mortise
C1525506|Ankle X-ray AP and lateral and Mortise
C1525506|Views AP & lateral & Mortise:Finding:Point in time:Ankle:Document:XR
C1525506|Views AP & lateral & Mortise:Find:Pt:Ankle:Doc:XR
C1524248|C-spine XR AP+Obl+Odont+Lat W FE
C1524248|Views AP & oblique & odontoid & lateral^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C1524248|Views AP & oblique & odontoid & lateral^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C1524248|Cervical spine X-ray AP and oblique and odontoid and lateral W flexion and W extension
C1525534|Ankle-L XR Lat+Mortise
C1525534|Ankle - left X-ray lateral and Mortise
C1525534|Views lateral & Mortise:Find:Pt:Ankle.left:Doc:XR
C1525534|Views lateral & Mortise:Finding:Point in time:Ankle.left:Document:XR
C1525570|Cerebral artery Fluoroscopic angiogram W contrast IA
C1525570|Cerebral a XRA W contr IA
C1525570|Views^W contrast Intra-arterial:Finding:Point in time:Cerebral artery:Document:XR.fluor.angio
C1525570|Views^W contrast IA:Find:Pt:Cerebral artery:Doc:XR.fluor.angio
C1525658|Multisection^WO & W contrast IV:Find:Pt:Mediastinum:Doc:MRI
C1525658|Mediastinum MRI WO+W contr IV
C1525658|Mediastinum MRI WO and W contrast IV
C1525658|Multisection^WO & W contrast Intravenous:Finding:Point in time:Mediastinum:Document:MRI
C1525703|Bones X-ray survey for metastasis
C1525703|Bones XR Survey for Metastasis
C1525703|Views survey for metastasis:Find:Pt:Bones:Doc:XR
C1525703|Views survey for metastasis:Finding:Point in time:Bones:Document:XR
C1525713|Adrenal a-L XRA W contr IA
C1525713|Adrenal artery - left Fluoroscopic angiogram W contrast IA
C1525713|Views^W contrast IA:Find:Pt:Adrenal artery.left:Doc:XR.fluor.angio
C1525713|Views^W contrast Intra-arterial:Finding:Point in time:Adrenal artery.left:Document:XR.fluor.angio
C1525799|Skull.base CT
C1525799|Multisection:Find:Pt:Skull.base:Doc:CT
C1525799|Multisection:Finding:Point in time:Skull.base:Document:Computerized Tomography
C1525855|Ft-L XR W Stress
C1525855|Foot - left X-ray W manual stress
C1525855|Views^W manual stress:Find:Pt:Foot.left:Doc:XR
C1525855|Views^W manual stress:Finding:Point in time:Foot.left:Document:XR
C1524133|Ac arch+Carot a.com-R XRA W contr IA
C1524133|Aortic arch and Carotid artery.common - right Fluoroscopic angiogram W contrast IA
C1524133|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery.common.right:Doc:XR.fluor.angio
C1524133|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery.common.right:Document:XR.fluor.angio
C1525808|Multisection^WO & W contrast IV:Find:Pt:Spine vessels:Doc:MRI.angio
C1525808|Spine vessels MRI angiogram WO and W contrast IV
C1525808|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine vessels:Document:MRI.angio
C1525808|Spine ves MRI.Angio WO+W contr IV
C1525822|Finger fourth - bilateral X-ray
C1525822|Finger.4th-Bl XR
C1525822|Views:Finding:Point in time:Finger.fourth.bilateral:Document:XR
C1525822|Views:Find:Pt:Finger.fourth.bilateral:Doc:XR
C1525948|Pelvis XR Obl
C1525948|Pelvis XR +Obl
C1525948|Pelvis X-ray oblique
C1525948|Pelvis X-ray and oblique
C1525948|Views & oblique:Finding:Point in time:Pelvis:Document:XR
C1525948|Views oblique:Finding:Point in time:Pelvis:Document:XR
C1525948|Views oblique:Find:Pt:Pelvis:Doc:XR
C1525948|Views & oblique:Find:Pt:Pelvis:Doc:XR
C1525961|Wrist-R XRTomo
C1525961|Wrist - right X-ray tomograph
C1525961|Multisection:Find:Pt:Wrist.right:Doc:XR.tomo
C1525961|Multisection:Finding:Point in time:Wrist.right:Document:XR.tomo
C1525966|SIJ XR AP+Obl
C1525966|Sacroiliac Joint X-ray AP and oblique
C1525966|Views AP & oblique:Finding:Point in time:Sacroiliac joint:Document:XR
C1525966|Views AP & oblique:Find:Pt:Sacroiliac joint:Doc:XR
C1525997|Elbow - right X-ray 2 views
C1525997|Elbow-R XR 2V
C1525997|Views 2:Finding:Point in time:Elbow.right:Document:XR
C1525997|Views 2:Find:Pt:Elbow.right:Doc:XR
C1525998|Elbow-R XR 3V
C1525998|Elbow - right X-ray 3 views
C1525998|Views 3:Finding:Point in time:Elbow.right:Document:XR
C1525998|Views 3:Find:Pt:Elbow.right:Doc:XR
C1525999|Elbow - right X-ray 4 views
C1525999|Elbow-R XR 4V
C1525999|Views 4:Find:Pt:Elbow.right:Doc:XR
C1525999|Views 4:Finding:Point in time:Elbow.right:Document:XR
C1526014|Ft-R XR 2V stand
C1526014|Foot - right X-ray 2 views standing
C1526014|Views 2^standing:Find:Pt:Foot.right:Doc:XR
C1526014|Views 2^standing:Finding:Point in time:Foot.right:Document:XR
C1526035|Views AP & lateral:Finding:Point in time:Calcaneus.right:Document:XR
C1526035|Views AP & lateral:Find:Pt:Calcaneus.right:Doc:XR
C1526035|Deprecated Calcaneus - right X-ray AP and lateral
C1526035|Deprecated Heel-R XR AP+Lat
C1525127|Patella - right X-ray
C1525127|Patella-R XR
C1525127|Views:Find:Pt:Patella.right:Doc:XR
C1525127|Views:Finding:Point in time:Patella.right:Document:XR
C1526089|Ribs - right X-ray lateral
C1526089|Ribs-R XR Lat
C1526089|View lateral:Finding:Point in time:Ribs.right:Document:XR
C1526089|View lateral:Find:Pt:Ribs.right:Doc:XR
C1526160|Skull X-ray 4 views
C1526160|Skull XR 4V
C1526160|Views 4:Finding:Point in time:Skull:Document:XR
C1526160|Views 4:Find:Pt:Skull:Doc:XR
C1526181|Views^W contrast Intrasynovial:Finding:Point in time:Temporomandibular joint:Document:XR.fluor
C1526181|TMJ Flr W contr IS
C1526181|Views^W contrast IS:Find:Pt:Temporomandibular joint:Doc:XR.fluor
C1526181|Temporomandibular joint Fluoroscopy W contrast IS
C1526253|Chest X-ray W expiration
C1526253|Chest XR W Exp
C1526253|View^W expiration:Finding:Point in time:Chest:Document:XR
C1526253|View^W expiration:Find:Pt:Chest:Doc:XR
C1526272|US Guidance for needle biopsy of Thyroid
C1526272|Thyroid US Bx needle guid
C1526272|Guidance for biopsy.needle:Finding:Point in time:Thyroid:Document:Ultrasound
C1526272|Guidance for biopsy.needle:Find:Pt:Thyroid:Doc:US
C1526278|Parathyroid US
C1526278|Multisection:Finding:Point in time:Parathyroid:Document:Ultrasound
C1526278|Multisection:Find:Pt:Parathyroid:Doc:US
C1526305|Should-L XR AP+Transthoracic
C1526305|Shoulder - left X-ray AP and transthoracic
C1526305|Views AP & transthoracic:Finding:Point in time:Shoulder.left:Document:XR
C1526305|Views AP & transthoracic:Find:Pt:Shoulder.left:Doc:XR
C1526313|Breast duct - bilateral Mammogram W contrast intra duct
C1526313|Brst.duct-Bl Mam W contr intra Dct
C1526313|Views^W contrast intra duct:Find:Pt:Breast.duct.bilateral:Doc:Mam
C1526313|Views^W contrast intra duct:Finding:Point in time:Breast.duct.bilateral:Document:Mam
C1524492|Face MRI W contr IV
C1524492|Face MRI W contrast IV
C1524492|Multisection^W contrast IV:Find:Pt:Face:Doc:MRI
C1524492|Multisection^W contrast Intravenous:Finding:Point in time:Face:Document:MRI
C1524867|Hrt MRI WO contr
C1524867|Heart MRI WO contrast
C1524867|Multisection^WO contrast:Find:Pt:Heart:Doc:MRI
C1524867|Multisection^WO contrast:Finding:Point in time:Heart:Document:MRI
C1524873|Hip - left MRI WO contrast
C1524873|Hip-L MRI WO contr
C1524873|Multisection^WO contrast:Finding:Point in time:Hip.left:Document:MRI
C1524873|Multisection^WO contrast:Find:Pt:Hip.left:Doc:MRI
C1524905|Sacrum CT WO contr
C1524905|Sacrum CT WO contrast
C1524905|Multisection^WO contrast:Finding:Point in time:Sacrum:Document:Computerized Tomography
C1524905|Multisection^WO contrast:Find:Pt:Sacrum:Doc:CT
C1524546|Upper arm-R MRI W contr IV
C1524546|Upper arm - right MRI W contrast IV
C1524546|Multisection^W contrast Intravenous:Finding:Point in time:Upper arm.right:Document:MRI
C1524546|Multisection^W contrast IV:Find:Pt:Upper arm.right:Doc:MRI
C1524547|LE.joint MRI W contr IV
C1524547|Lower Extremity Joint MRI W contrast IV
C1524547|Multisection^W contrast IV:Find:Pt:Lower extremity.joint:Doc:MRI
C1524547|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.joint:Document:MRI
C1524217|Shoulder - left X-ray AP single view
C1524217|Should-L XR AP 1V
C1524217|View AP:Find:Pt:Shoulder.left:Doc:XR
C1524217|View AP:Finding:Point in time:Shoulder.left:Document:XR
C1524297|Salivary gland CT Bx guid
C1524297|CT Guidance for biopsy of Salivary gland
C1524297|Guidance for biopsy:Find:Pt:Salivary gland:Doc:CT
C1524297|Guidance for biopsy:Finding:Point in time:Salivary gland:Document:Computerized Tomography
C1524597|Lower leg-R MRI W contr IV
C1524597|Lower leg - right MRI W contrast IV
C1524597|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg.right:Document:MRI
C1524597|Multisection^W contrast IV:Find:Pt:Lower leg.right:Doc:MRI
C1524599|Uterus MRI W contr IV
C1524599|Uterus MRI W contrast IV
C1524599|Multisection^W contrast Intravenous:Finding:Point in time:Uterus:Document:MRI
C1524599|Multisection^W contrast IV:Find:Pt:Uterus:Doc:MRI
C1524651|Knee - bilateral X-ray 4 views
C1524651|Knee-Bl XR 4V
C1524651|Views 4:Find:Pt:Knee.bilateral:Doc:XR
C1524651|Views 4:Finding:Point in time:Knee.bilateral:Document:XR
C1524751|Multisection^WO & W contrast IV:Find:Pt:Hip.right:Doc:MRI
C1524751|Hip-R MRI WO+W contr IV
C1524751|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip.right:Document:MRI
C1524751|Hip - right MRI WO and W contrast IV
C1525033|Femur-Bl XR AP+Lat
C1525033|Femur - bilateral X-ray AP and lateral
C1525033|Views AP & lateral:Finding:Point in time:Femur.bilateral:Document:XR
C1525033|Views AP & lateral:Find:Pt:Femur.bilateral:Doc:XR
C1525042|Hip-Bl XR AP+Lat
C1525042|Hip - bilateral X-ray AP and lateral
C1525042|Views AP & lateral:Find:Pt:Hip.bilateral:Doc:XR
C1525042|Views AP & lateral:Finding:Point in time:Hip.bilateral:Document:XR
C1525058|Toes-L XR AP+Lat
C1525058|Toes - left X-ray AP and lateral
C1525058|Views AP & lateral:Finding:Point in time:Toes.left:Document:XR
C1525058|Views AP & lateral:Find:Pt:Toes.left:Doc:XR
C1524799|Multisection^WO & W contrast IV:Find:Pt:Portal vein:Doc:MRI.angio
C1524799|Portal v MRI.Angio WO+W contr IV
C1524799|Portal vein MRI angiogram WO and W contrast IV
C1524799|Multisection^WO & W contrast Intravenous:Finding:Point in time:Portal vein:Document:MRI.angio
C1525080|Hand-Bl XR PA+Lat
C1525080|Hand - bilateral X-ray PA and lateral
C1525080|Views PA & lateral:Finding:Point in time:Hand.bilateral:Document:XR
C1525080|Views PA & lateral:Find:Pt:Hand.bilateral:Doc:XR
C1830195|Stom Flr Replac of PC drain tube guid
C1830195|Fluoroscopy Guidance for replacement of percutaneous drainage tube in Stomach
C1830195|Guidance for replacement of percutaneous drainage tube:Finding:Point in time:Stomach:Document:XR.fluor
C1830195|Guidance for replacement of percutaneous drainage tube:Find:Pt:Stomach:Doc:XR.fluor
C1830210|Upper extremity - right Vessels CT angiogram WO and W contrast IV
C1830210|EU ves-R CT.Angio WO+W contr IV
C1830210|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.right>Vessels:Doc:CT.angio
C1830210|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.right>Vessels:Document:Computerized Tomography.angio
C1830214|Multisection^WO & W reduced contrast volume IV:Find:Pt:Pelvis:Doc:CT
C1830214|Multisection^WO & W reduced contrast volume Intravenous:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1830214|Pelvis CT WO+W red contr vol IV
C1830214|Pelvis CT WO and W reduced contrast volume IV
C1830242|Abd Flr
C1830242|Abdomen Fluoroscopy
C1830242|Views:Find:Pt:Abdomen:Doc:XR.fluor
C1830242|Views:Finding:Point in time:Abdomen:Document:XR.fluor
C1830255|Breast - right FFD mammogram screening
C1830255|Views screening:Finding:Point in time:Breast.right:Document:Mam.FFD
C1830255|Brst-R FFDM Screening
C1830255|Views screening:Find:Pt:Breast.right:Doc:Mam.FFD
C1830279|Ankle-L XR GE 3V
C1830279|Ankle - left X-ray GE 3 views
C1830279|Views GE 3:Find:Pt:Ankle.left:Doc:XR
C1830279|Views GE 3:Finding:Point in time:Ankle.left:Document:XR
C1715373|Liver CT Ablation guid
C1715373|CT Guidance for ablation of tissue of Liver
C1715373|Guidance for ablation of tissue:Find:Pt:Abdomen>Liver:Doc:CT
C1715373|Guidance for ablation of tissue:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1715388|Mandible CT limited
C1715388|Mandible CT Ltd
C1715388|Multisection limited:Find:Pt:Mandible:Doc:CT
C1715388|Multisection limited:Finding:Point in time:Mandible:Document:Computerized Tomography
C1715390|Brst-Bl CT WO contr
C1715390|Breast - bilateral CT WO contrast
C1715390|Multisection^WO contrast:Find:Pt:Breast.bilateral:Doc:CT
C1715390|Multisection^WO contrast:Finding:Point in time:Breast.bilateral:Document:Computerized Tomography
C1715426|US Guidance for fine needle aspiration of Liver
C1715426|Liver US FNA Asp
C1715426|Guidance for aspiration.fine needle:Finding:Point in time:Liver:Document:Ultrasound
C1715426|Guidance for aspiration.fine needle:Find:Pt:Liver:Doc:US
C1715478|Fluoroscopy Guidance for fine needle aspiration of Pancreas
C1715478|Pancreas Flr FNA Asp
C1715478|Guidance for aspiration.fine needle:Finding:Point in time:Pancreas:Document:XR.fluor
C1715478|Guidance for aspiration.fine needle:Find:Pt:Pancreas:Doc:XR.fluor
C1644152|Ribs - left X-ray portable
C1644152|Ribs-L XR port
C1644152|Views portable:Find:Pt:Ribs.left:Doc:XR
C1644152|Views portable:Finding:Point in time:Ribs.left:Document:XR
C1646773|Guidance for biopsy:Find:Pt:Chest>Pleura:Doc:US
C1646773|Guidance for biopsy:Finding:Point in time:Chest>Pleura:Document:Ultrasound
C1646773|US Guidance for biopsy of Chest Pleura
C1646773|Chest Pleura US Bx guid
C1714528|Sinuses X-ray GE 3 views
C1714528|Sinuses XR GE 3V
C1714528|Views GE 3:Finding:Point in time:Sinuses:Document:XR
C1714528|Views GE 3:Find:Pt:Sinuses:Doc:XR
C1714913|Lower leg vessels - bilateral MRI angiogram W contrast IV
C1714913|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg vessels.bilateral:Document:MRI.angio
C1714913|Multisection^W contrast IV:Find:Pt:Lower leg vessels.bilateral:Doc:MRI.angio
C1714913|Lower leg ves-Bl MRI.Angio W contr IV
C1714788|Elbow-L MRI Dyn W contr IV
C1714788|Elbow - left MRI dynamic W contrast IV
C1714788|Multisection dynamic^W contrast IV:Find:Pt:Elbow.left:Doc:MRI
C1714788|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Elbow.left:Document:MRI
C1714956|T+L-spine XR Scoli AP upr+sup
C1714956|Views scoliosis AP^upright & supine:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1714956|Spine Thoracic and Lumbar X-ray scoliosis AP upright and supine
C1714956|Views scoliosis AP^upright & supine:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1715034|Spleen SPECT flow
C1715034|Spleen SPECT Flow W RNC IV
C1715034|Multisection flow^W radionuclide IV:Find:Pt:Spleen:Doc:Radnuc.SPECT
C1715034|Multisection flow^W radionuclide Intravenous:Finding:Point in time:Spleen:Document:Radnuc.SPECT
C1715110|C+T+L-spine XR 2V
C1715110|Spine Cervical and Thoracic and Lumbar X-ray 2 views
C1715110|Views 2:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:XR
C1715110|Views 2:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:XR
C1715111|CTJ XR AP+Lat
C1715111|Spine Cervicothoracic Junction X-ray AP and lateral
C1715111|Views AP & lateral:Find:Pt:Spine.cervicothoracic junction:Doc:XR
C1715111|Views AP & lateral:Finding:Point in time:Spine.cervicothoracic junction:Document:XR
C1715117|L-spine XR Obl
C1715117|Views oblique:Finding:Point in time:Spine.lumbar:Document:XR
C1715117|Views oblique:Find:Pt:Spine.lumbar:Doc:XR
C1715117|Lumbar spine X-ray oblique
C1626319|T+L-spine XR Scoli AP 1V Stand+R-bending
C1626319|View scoliosis AP^standing & W R-bending:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1626319|View scoliosis AP^standing & W R-bending:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1626319|Spine Thoracic and Lumbar X-ray scoliosis AP standing and W right bending
C1639905|Extremity vein - right US
C1639905|Extr v-R US
C1639905|Multisection:Finding:Point in time:Extremity vein.right:Document:Ultrasound
C1639905|Multisection:Find:Pt:Extremity vein.right:Doc:US
C1627298|C-spine XR +Obl
C1627298|Views & oblique:Finding:Point in time:Spine.cervical:Document:XR
C1627298|Views & oblique:Find:Pt:Spine.cervical:Doc:XR
C1627298|Cervical spine X-ray and oblique
C1643242|Face XR port
C1643242|Facial bones X-ray portable
C1643242|Views portable:Find:Pt:Facial bones:Doc:XR
C1643242|Views portable:Finding:Point in time:Facial bones:Document:XR
C1642595|Hand-R XR Ltd
C1642595|Hand - right X-ray limited
C1642595|Views limited:Finding:Point in time:Hand.right:Document:XR
C1642595|Views limited:Find:Pt:Hand.right:Doc:XR
C1653523|Views PA & lateral:Finding:Point in time:Chest:Narrative:XR
C1653523|Chest XR PA+Lat
C1653523|Chest X-ray PA and lateral
C1653523|Views PA & lateral:Finding:Point in time:Chest:Document:XR
C1653523|Views PA & lateral:Find:Pt:Chest:Doc:XR
C1630749|Multisection^WO & W contrast IV:Find:Pt:Abdomen+Pelvis:Doc:CT
C1630749|Abdomen and Pelvis CT WO and W contrast IV
C1630749|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis:Document:Computerized Tomography
C1630749|Abd+Pelvis CT WO+W contr IV
C1631257|Chest and Abdomen CT WO contrast
C1631257|Chest+Abd CT WO contr
C1631257|Multisection^WO contrast:Find:Pt:Chest+Abdomen:Doc:CT
C1631257|Multisection^WO contrast:Finding:Point in time:Chest+Abdomen:Document:Computerized Tomography
C1632954|SPECT for tumor W Tl-201 IV
C1632954|Multisection for tumor^W Tl-201 IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1632954|Multisection for tumor^W Tl-201 Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1632337|Pelv ves CT.Angio W contr IV
C1632337|Multisection^W contrast IV:Find:Pt:Pelvis>Vessels:Doc:CT.angio
C1632337|Pelvic vessels CT angiogram W contrast IV
C1632337|Multisection^W contrast Intravenous:Finding:Point in time:Pelvis>Vessels:Document:Computerized Tomography.angio
C1978446|Ankle+Foot-R XR
C1978446|Ankle - right and Foot - right X-ray
C1978446|Views:Find:Pt:Ankle.right+Foot.right:Doc:XR
C1978446|Views:Finding:Point in time:Ankle.right+Foot.right:Document:XR
C1954306|Lower extremity vein - left US
C1954306|LE v-L US
C1954306|Multisection:Find:Pt:Lower extremity vein.left:Doc:US
C1954306|Multisection:Finding:Point in time:Lower extremity vein.left:Document:Ultrasound
C1954369|Mammogram Guidance for sentinel lymph node injection of Breast
C1954369|Brst Mam Sentinel LN inj guid
C1954369|Guidance for sentinel lymph node injection:Finding:Point in time:Breast:Document:Mam
C1954369|Guidance for sentinel lymph node injection:Find:Pt:Breast:Doc:Mam
C1952652|Ribs-L+Chest XR GE 3V+PA Chst
C1952652|Ribs - left and Chest X-ray GE 3 and PA Chest views
C1952652|Views GE 3 & PA chest:Finding:Point in time:Ribs.left+Chest:Document:XR
C1952652|Views GE 3 & PA chest:Find:Pt:Ribs.left+Chest:Doc:XR
C1952654|Mastoid - right X-ray 1 or 2 views
C1952654|Mastoid-R XR 1V or 2V
C1952654|Views 1 or 2:Find:Pt:Mastoid.right:Doc:XR
C1952654|Views 1 or 2:Finding:Point in time:Mastoid.right:Document:XR
C3655047|Surg Spec XR
C3655047|Views:Find:Pt:Surgical specimen:Doc:XR
C3655047|Views:Finding:Point in time:Surgical specimen:Document:XR
C3655047|Surgical specimen X-ray
C3533570|Guidance for ambulatory phlebectomy:Find:Pt:Extremity vein.right:Doc:US
C3533570|Extr v-R US Amb phleb guid
C3533570|Guidance for ambulatory phlebectomy:Finding:Point in time:Extremity vein.right:Document:Ultrasound
C3533570|US Guidance for ambulatory phlebectomy of Extremity vein - right
C3533566|US Guidance for injection of sclerosing agent of Extremity veins - bilateral
C3533566|Extr vv-Bl US Sclerosing agent inj guid
C3533566|Guidance for injection of sclerosing agent:Find:Pt:Extremity veins.bilateral:Doc:US
C3533566|Guidance for injection of sclerosing agent:Finding:Point in time:Extremity veins.bilateral:Document:Ultrasound
C3533563|XXX Flr PN DN guid
C3533563|Fluoroscopy Guidance for peripheral nerve denervation of Unspecified body region
C3533563|Guidance for peripheral nerve denervation:Find:Pt:XXX:Doc:XR.fluor
C3533563|Guidance for peripheral nerve denervation:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C3262997|Hand - bilateral MRI WO and W contrast IV
C3262997|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hand.bilateral:Document:MRI
C3262997|Hand-Bl MRI WO+W contr IV
C3262997|Multisection^WO & W contrast IV:Find:Pt:Hand.bilateral:Doc:MRI
C3263030|Multisection^WO & W contrast Intrasynovial:Finding:Point in time:Hip.right:Document:MRI
C3263030|Hip - right MRI WO and W contrast IS
C3263030|Multisection^WO & W contrast IS:Find:Pt:Hip.right:Doc:MRI
C3263030|Hip-R MRI WO+W contr IS
C3263036|XXX MRI WO contr
C3263036|Unspecified body region MRI WO contrast
C3263036|Multisection^WO contrast:Find:Pt:XXX:Doc:MRI
C3263036|Multisection^WO contrast:Finding:Point in time:To be specified in another part of the message:Document:MRI
C3203435|Ft-R XR 1V
C3203435|Foot - right X-ray Single view
C3203435|View 1:Find:Pt:Foot.right:Doc:XR
C3203435|View 1:Finding:Point in time:Foot.right:Document:XR
C3262911|Knee - bilateral CT W contrast IV
C3262911|Knee-Bl CT W contr IV
C3262911|Multisection^W contrast Intravenous:Finding:Point in time:Knee.bilateral:Document:Computerized Tomography
C3262911|Multisection^W contrast IV:Find:Pt:Knee.bilateral:Doc:CT
C3262927|Extremity - left CT WO contrast
C3262927|Extr-L CT WO contr
C3262927|Multisection^WO contrast:Find:Pt:Extremity.left:Doc:CT
C3262927|Multisection^WO contrast:Finding:Point in time:Extremity.left:Document:Computerized Tomography
C0942174|Tib+Fib-L XR
C0942174|Tibia - left and Fibula - left X-ray
C0942174|Views:Finding:Point in time:Tibia.left+Fibula.left:Document:XR
C0942174|Views:Find:Pt:Tibia.left+Fibula.left:Doc:XR
C0942195|TO-L MRI WO+W contr IV
C0942195|Multisection^WO & W contrast IV:Find:Pt:Thoracic outlet.left:Doc:MRI
C0942195|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thoracic outlet.left:Document:MRI
C0942195|Thoracic outlet - left MRI WO and W contrast IV
C0942212|Ankle - bilateral MRI
C0942212|Ankle-Bl MRI
C0942212|Multisection:Finding:Point in time:Ankle.bilateral:Document:MRI
C0942212|Multisection:Find:Pt:Ankle.bilateral:Doc:MRI
C0942234|Upper extremity - right MRI
C0942234|UE-R MRI
C0942234|Multisection:Find:Pt:Upper extremity.right:Doc:MRI
C0942234|Multisection:Finding:Point in time:Upper extremity.right:Document:MRI
C0942298|Cent v-L XRA Cath plac guid W contr IV
C0942298|Fluoroscopic angiogram Guidance for placement of catheter in Central vein - left-- W contrast IV
C0942298|Guidance for placement of catheter^W contrast Intravenous:Finding:Point in time:Central vein.left:Document:XR.fluor.angio
C0942298|Guidance for placement of catheter^W contrast IV:Find:Pt:Central vein.left:Doc:XR.fluor.angio
C0945339|Brst-L Mam Bx guid
C0945339|Mammogram Guidance for biopsy of Breast - left
C0945339|Guidance for biopsy:Find:Pt:Breast.left:Doc:Mam
C0945339|Guidance for biopsy:Finding:Point in time:Breast.left:Document:Mam
C0945345|Vein-Bl VD admin into cath
C0945345|Administration of vasodilator into catheter of Vein - bilateral
C0945345|Administration of vasodilator into catheter:Finding:Point in time:Vein.bilateral:Document
C0945345|Administration of vasodilator into catheter:Find:Pt:Vein.bilateral:Doc
C0882545|Pelvis X-ray pelvimetry
C0882545|Pelvis XR Pelvimetry
C0882545|View pelvimetry:Find:Pt:Pelvis:Doc:XR
C0882545|View pelvimetry:Finding:Point in time:Pelvis:Document:XR
C0882077|Bone density:Mass Aeric:Point in time:Radius+Ulna:Quantitative:XR.DXA
C0882077|Radius and Ulna DXA Bone density
C0882077|Bone density:MAric:Pt:Radius+Ulna:Qn:XR.DXA
C0882077|Radius+Ulna DXA BDM
C0882081|Kidney US Drain guid
C0882081|US Guidance for drainage of Kidney
C0882081|Guidance for drainage:Find:Pt:Kidney:Doc:US
C0882081|Guidance for drainage:Finding:Point in time:Kidney:Document:Ultrasound
C2608010|Views:Finding:Point in time:Shoulder:Narrative:XR
C2608010|Should XR
C2608010|Shoulder X-ray
C2608010|Views:Find:Pt:Shoulder:Doc:XR
C2608010|Views:Finding:Point in time:Shoulder:Document:XR
C0882153|Views:Finding:Point in time:Sternoclavicular joints:Narrative:XR
C0882153|SC joints XR
C0882153|Sternoclavicular Joints X-ray
C0882153|Views:Finding:Point in time:Sternoclavicular joints:Document:XR
C0882153|Views:Find:Pt:Sternoclavicular joints:Doc:XR
C0882157|Stomach Scan for gastric emptying solid phase W Tc-99m SC PO
C0882157|Stom RI SPGE W Tc99mSC PO
C0882157|Views for gastric emptying solid phase^W Tc-99m SC PO:Find:Pt:Stomach:Doc:Radnuc
C0882157|Views for gastric emptying solid phase^W Tc-99m Subcutaneous Oral:Finding:Point in time:Stomach:Document:Radnuc
C0882164|Three vessels Fluoroscopic angiogram W contrast
C0882164|Views^W contrast:Finding:Point in time:Three vessels:Document:XR.fluor.angio
C0882164|Views^W contrast:Find:Pt:Three vessels:Doc:XR.fluor.angio
C0882164|3 vess XRA W contr
C0882220|Unspecified body region Fluoroscopy during surgery
C0882220|XXX Flr in Surg
C0882220|Views^during surgery:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C0882220|Views^during surgery:Find:Pt:XXX:Doc:XR.fluor
C0942130|LE-Bl XR
C0942130|Lower extremity - bilateral X-ray
C0942130|Views:Find:Pt:Lower extremity.bilateral:Doc:XR
C0942130|Views:Finding:Point in time:Lower extremity.bilateral:Document:XR
C0942133|Upper extremity - right X-ray
C0942133|UE-R XR
C0942133|Views:Finding:Point in time:Upper extremity.right:Document:XR
C0942133|Views:Find:Pt:Upper extremity.right:Doc:XR
C0947254|Finger-L XR
C0947254|Finger - left X-ray
C0947254|Views:Finding:Point in time:Finger.left:Document:XR
C0947254|Views:Find:Pt:Finger.left:Doc:XR
C0881817|Bones long X-ray survey
C0881817|Bones.long XR Survey
C0881817|Views survey:Find:Pt:Bones.long:Doc:XR
C0881817|Views survey:Finding:Point in time:Bones.long:Document:XR
C0881825|Multisection^WO & W contrast Intravenous & W anesthesia:Finding:Point in time:Brain:Document:MRI
C0881825|Brain MRI WO and W contrast IV and W anesthesia
C0881825|Multisection^WO & W contrast IV & W anesthesia:Find:Pt:Brain:Doc:MRI
C0881825|Brain MRI WO+W contr IV+Anesthesia
C0881850|Carot a XRA W contr IA
C0881850|Carotid artery Fluoroscopic angiogram W contrast IA
C0881850|Views^W contrast IA:Find:Pt:Carotid artery:Doc:XR.fluor.angio
C0881850|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery:Document:XR.fluor.angio
C0882527|Chest Flr in Surg
C0882527|Chest Fluoroscopy during surgery
C0882527|View^during surgery:Finding:Point in time:Chest:Document:XR.fluor
C0882527|View^during surgery:Find:Pt:Chest:Doc:XR.fluor
C0881883|Aorta XRA W contr IA
C0881883|Aorta Fluoroscopic angiogram W contrast IA
C0881883|Views^W contrast IA:Find:Pt:Aorta:Doc:XR.fluor.angio
C0881883|Views^W contrast Intra-arterial:Finding:Point in time:Aorta:Document:XR.fluor.angio
C0881893|Colon Fluoroscopy transit Post solid contrast
C0881893|Colon Flr transit p solid contr PO
C0881893|View transit^post solid contrast PO:Find:Pt:Colon:Doc:XR.fluor
C0881893|View transit^post solid contrast Oral:Finding:Point in time:Colon:Document:XR.fluor
C0881971|CT Guidance for injection of Joint space
C0881971|Guidance for injection:Find:Pt:Joint space:Doc:CT
C0881971|Guidance for injection:Finding:Point in time:Joint space:Document:Computerized Tomography
C0881971|Joint space CT Inj guid
C0881989|Multisection:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:XR.tomo
C0881989|Multisection:Find:Pt:Kidney.bilateral:Doc:XR.tomo
C0881989|Kidney - bilateral X-ray tomograph
C0881989|Multisection:Finding:Point in time:Kidney.bilateral:Document:XR.tomo
C0881989|Kdny-Bl XRTomo
C0882013|US Guidance for biopsy of Liver
C0882013|Liver US Bx guid
C0882013|Guidance for biopsy:Finding:Point in time:Liver:Document:Ultrasound
C0882013|Guidance for biopsy:Find:Pt:Liver:Doc:US
C1114564|T-spine XR AP+Lat port
C1114564|Views AP & lateral portable:Find:Pt:Spine.thoracic:Doc:XR
C1114564|Views AP & lateral portable:Finding:Point in time:Spine.thoracic:Document:XR
C1114564|Thoracic spine X-ray AP and lateral portable
C1114568|T-spine XR Obl port
C1114568|View oblique portable:Find:Pt:Spine.thoracic:Doc:XR
C1114568|View oblique portable:Finding:Point in time:Spine.thoracic:Document:XR
C1114568|Thoracic spine X-ray oblique portable
C2608011|View 1 portable:Finding:Point in time:Spine.lumbar:Narrative:XR
C2608011|L-spine XR 1V port
C2608011|View 1 portable:Find:Pt:Spine.lumbar:Doc:XR
C2608011|View 1 portable:Finding:Point in time:Spine.lumbar:Document:XR
C2608011|Lumbar spine X-ray Single view portable
C1114679|Views:Finding:Point in time:Sacrum:Narrative:XR
C1114679|Sacrum X-ray
C1114679|Sacrum XR
C1114679|Views:Finding:Point in time:Sacrum:Document:XR
C1114679|Views:Find:Pt:Sacrum:Doc:XR
C1114686|Cervicocerebral a XRA W contr IA
C1114686|Cervicocerebral artery Fluoroscopic angiogram W contrast IA
C1114686|Views^W contrast IA:Find:Pt:Cervicocerebral artery:Doc:XR.fluor.angio
C1114686|Views^W contrast Intra-arterial:Finding:Point in time:Cervicocerebral artery:Document:XR.fluor.angio
C1116465|Guidance for drainage of abscess:Find:Pt:XXX:Doc:CT
C1116465|CT Guidance for drainage of abscess of Unspecified body region
C1116465|Guidance for drainage of abscess:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1116465|XXX CT Abscess drain guid
C1526824|Ribs Ant+Post-L XR
C1526824|Ribs anterior and posterior - left X-ray
C1526824|Views:Find:Pt:Ribs.anterior+posterior.left:Doc:XR
C1526824|Views:Finding:Point in time:Ribs.anterior+posterior.left:Document:XR
C1543457|Ft-R XR AP+Lat stand
C1543457|Foot - right X-ray AP and lateral standing
C1543457|Views AP & lateral^standing:Finding:Point in time:Foot.right:Document:XR
C1543457|Views AP & lateral^standing:Find:Pt:Foot.right:Doc:XR
C1526025|Radius+Ulna-R XR Obl
C1526025|Radius+Ulna-R XR +Obl
C1526025|Radius - right and Ulna - right X-ray and oblique
C1526025|Radius - right and Ulna - right X-ray oblique
C1526025|Views oblique:Find:Pt:Radius.right+Ulna.right:Doc:XR
C1526025|Views oblique:Finding:Point in time:Radius.right+Ulna.right:Document:XR
C1526025|Views & oblique:Find:Pt:Radius.right+Ulna.right:Doc:XR
C1526025|Views & oblique:Finding:Point in time:Radius.right+Ulna.right:Document:XR
C1543477|Wrist-R XR +Carpal Tunnel
C1543477|Wrist-R XR V1 tunnel.carpal
C1543477|Wrist - right X-ray tunnel.carpal
C1543477|Wrist - right X-ray and carpal tunnel
C1543477|Views & carpal tunnel:Finding:Point in time:Wrist.right:Document:XR
C1543477|View tunnel.carpal:Find:Pt:Wrist.right:Doc:XR
C1543477|View tunnel.carpal:Finding:Point in time:Wrist.right:Document:XR
C1543477|Views & carpal tunnel:Find:Pt:Wrist.right:Doc:XR
C1543493|Deprecated KD-Bl+CS US
C1543493|Multisection:Find:Pt:Kidney.bilateral+Collecting system:Nar:US
C1543493|Deprecated Kidney Bilateral & Collecting system US Multisection
C1543493|Multisection:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:Ultrasound
C1543495|Renal ves-Bl DOP
C1543495|Renal vessels - bilateral US.doppler
C1543495|Multisection:Find:Pt:Renal vessels.bilateral:Doc:US.doppler
C1543495|Multisection:Finding:Point in time:Renal vessels.bilateral:Document:Ultrasound.doppler
C1543784|Hrt RI PF W Stress+W Tc99mMIBI IV
C1543784|Heart Scan perfusion W stress and W Tc-99m Sestamibi IV
C1543784|Views perfusion^W stress & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543784|Views perfusion^W stress & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542847|Thyroid RI W Tc99mMIBI IV
C1542847|Thyroid Scan W Tc-99m Sestamibi IV
C1542847|Views^W Tc-99m Sestamibi Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1542847|Views^W Tc-99m Sestamibi IV:Find:Pt:Thyroid:Doc:Radnuc
C1542905|RI Ltd W In-111 Satmb IV
C1542905|Scan limited W In-111 Satumomab IV
C1542905|Views limited^W In-111 Satumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542905|Views limited^W In-111 Satumomab IV:Find:Pt:^Patient:Doc:Radnuc
C1542858|Joint Scan multiple areas W radionuclide XXX
C1542858|Joint RI Mul Areas W RNC XXX
C1542858|Views multiple areas^W radionuclide XXX:Find:Pt:Joint:Doc:Radnuc
C1542858|Views multiple areas^W radionuclide XXX:Finding:Point in time:Joint:Document:Radnuc
C1542859|Joint SPECT W RNC IV
C1542859|Joint SPECT
C1542859|Multisection^W radionuclide Intravenous:Finding:Point in time:Joint:Document:Radnuc.SPECT
C1542859|Multisection^W radionuclide IV:Find:Pt:Joint:Doc:Radnuc.SPECT
C1543525|Extr v DOP
C1543525|Extremity vein US.doppler
C1543525|Multisection:Finding:Point in time:Extremity vein:Document:Ultrasound.doppler
C1543525|Multisection:Find:Pt:Extremity vein:Doc:US.doppler
C1543148|Fluoroscopy Guidance for needle localization of Unspecified body region
C1543148|XXX Flr Needle local guid
C1543148|Guidance for needle localization:Find:Pt:XXX:Doc:XR.fluor
C1543148|Guidance for needle localization:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1543149|MRI Guidance for needle localization of Unspecified body region
C1543149|XXX MRI Needle local guid
C1543149|Guidance for needle localization:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1543149|Guidance for needle localization:Find:Pt:XXX:Doc:MRI
C1543154|UE MRI WO contr
C1543154|Upper extremity MRI WO contrast
C1543154|Multisection^WO contrast:Find:Pt:Upper extremity:Doc:MRI
C1543154|Multisection^WO contrast:Finding:Point in time:Upper extremity:Document:MRI
C1543579|Extr ves-R DOP
C1543579|Extremity vessels - right US.doppler
C1543579|Multisection:Finding:Point in time:Extremity vessels.right:Document:Ultrasound.doppler
C1543579|Multisection:Find:Pt:Extremity vessels.right:Doc:US.doppler
C1543583|Upper extremity vein - right US.doppler
C1543583|UE v-R DOP
C1543583|Multisection:Finding:Point in time:Upper extremity vein.right:Document:Ultrasound.doppler
C1543583|Multisection:Find:Pt:Upper extremity vein.right:Doc:US.doppler
C1524260|Pelvis+Hip-R XR AP+Lat Frog
C1524260|Pelvis and Hip - right X-ray AP and lateral frog
C1524260|Views AP & lateral frog:Find:Pt:Pelvis+Hip.right:Doc:XR
C1524260|Views AP & lateral frog:Finding:Point in time:Pelvis+Hip.right:Document:XR
C1543720|Hrt SPECT Rest+W RNC IV
C1543720|Heart SPECT at rest and W radionuclide IV
C1543720|Multisection^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543720|Multisection^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543377|LE MRI WO+W contr IV
C1543377|Multisection^WO & W contrast IV:Find:Pt:Lower extremity:Doc:MRI
C1543377|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity:Document:MRI
C1543377|Lower extremity MRI WO and W contrast IV
C1527069|Prostate CT
C1527069|Multisection:Find:Pt:Prostate:Doc:CT
C1527069|Multisection:Finding:Point in time:Prostate:Document:Computerized Tomography
C1524175|Sacrum+Coccyx MRI
C1524175|Sacrum and Coccyx MRI
C1524175|Multisection:Finding:Point in time:Sacrum+Coccyx:Document:MRI
C1524175|Multisection:Find:Pt:Sacrum+Coccyx:Doc:MRI
C1524191|Lower extremity veins MRI angiogram
C1524191|LE vv MRI.Angio
C1524191|Multisection:Finding:Point in time:Lower extremity veins:Document:MRI.angio
C1524191|Multisection:Find:Pt:Lower extremity veins:Doc:MRI.angio
C1524833|Elbow-R MRI WO contr
C1524833|Elbow - right MRI WO contrast
C1524833|Multisection^WO contrast:Finding:Point in time:Elbow.right:Document:MRI
C1524833|Multisection^WO contrast:Find:Pt:Elbow.right:Doc:MRI
C1524835|Lower extremity vessels - bilateral MRI angiogram WO contrast
C1524835|Multisection^WO contrast:Find:Pt:Lower extremity vessels.bilateral:Doc:MRI.angio
C1524835|Multisection^WO contrast:Finding:Point in time:Lower extremity vessels.bilateral:Document:MRI.angio
C1524835|LE ves-Bl MRI.Angio WO contr
C1525101|Temporal bone CT
C1525101|Multisection:Find:Pt:Temporal bone:Doc:CT
C1525101|Multisection:Finding:Point in time:Temporal bone:Document:Computerized Tomography
C1525118|Adrenal vessels MRI angiogram
C1525118|Adrenal ves MRI.Angio
C1525118|Multisection:Find:Pt:Adrenal vessels:Doc:MRI.angio
C1525118|Multisection:Finding:Point in time:Adrenal vessels:Document:MRI.angio
C1524440|Neck ves MRI.Angio
C1524440|Neck vessels MRI angiogram
C1524440|Multisection:Finding:Point in time:Neck vessels:Document:MRI.angio
C1524440|Multisection:Find:Pt:Neck vessels:Doc:MRI.angio
C1524467|SIJ CT W contr IS
C1524467|Multisection^W contrast IS:Find:Pt:Sacroiliac joint:Doc:CT
C1524467|Multisection^W contrast Intrasynovial:Finding:Point in time:Sacroiliac joint:Document:Computerized Tomography
C1524467|Sacroiliac Joint CT W contrast IS
C1525311|Elbow X-ray Jones
C1525311|Elbow XR Jones
C1525311|View Jones:Finding:Point in time:Elbow:Document:XR
C1525311|View Jones:Find:Pt:Elbow:Doc:XR
C1525201|Head vv MRI.Angio W contr IV
C1525201|Head veins MRI angiogram W contrast IV
C1525201|Multisection^W contrast Intravenous:Finding:Point in time:Head veins:Document:MRI.angio
C1525201|Multisection^W contrast IV:Find:Pt:Head veins:Doc:MRI.angio
C1525205|Head vessels CT angiogram W contrast IV
C1525205|Multisection^W contrast IV:Find:Pt:Head>Vessels:Doc:CT.angio
C1525205|Multisection^W contrast Intravenous:Finding:Point in time:Head>Vessels:Document:Computerized Tomography.angio
C1525205|Head vess CT.Angio W contr IV
C1526994|Adrenal gland MRI
C1526994|Adrenal MRI
C1526994|Multisection:Finding:Point in time:Adrenal gland:Document:MRI
C1526994|Multisection:Find:Pt:Adrenal gland:Doc:MRI
C1525458|Humerus XR Transthoracic
C1525458|Humerus X-ray transthoracic
C1525458|View transthoracic:Find:Pt:Humerus:Doc:XR
C1525458|View transthoracic:Finding:Point in time:Humerus:Document:XR
C1525464|Brst-Bl Mam True Lat
C1525464|Breast - bilateral Mammogram true lateral
C1525464|View true lateral:Finding:Point in time:Breast.bilateral:Document:Mam
C1525464|View true lateral:Find:Pt:Breast.bilateral:Doc:Mam
C1524221|Abdomen X-ray upright
C1524221|Abd XR Upr
C1524221|View upright:Finding:Point in time:Abdomen:Document:XR
C1524221|View upright:Find:Pt:Abdomen:Doc:XR
C1524226|Shoulder - left X-ray West Point
C1524226|Should-L XR West Point
C1524226|View West Point:Find:Pt:Shoulder.left:Doc:XR
C1524226|View West Point:Finding:Point in time:Shoulder.left:Document:XR
C1525505|Pelvis+Hip-L XR AP+Lat Frog
C1525505|Pelvis and Hip - left X-ray AP and lateral frog
C1525505|Views AP & lateral frog:Find:Pt:Pelvis+Hip.left:Doc:XR
C1525505|Views AP & lateral frog:Finding:Point in time:Pelvis+Hip.left:Document:XR
C1525539|Should-L XR Outlet+Y
C1525539|Shoulder - left X-ray outlet and Y
C1525539|Views outlet & Y:Find:Pt:Shoulder.left:Doc:XR
C1525539|Views outlet & Y:Finding:Point in time:Shoulder.left:Document:XR
C1525557|Should-L XR Grashey+Ax+Outlet
C1525557|Shoulder - left X-ray Grashey and axillary and outlet
C1525557|Views Grashey & axillary & outlet:Find:Pt:Shoulder.left:Doc:XR
C1525557|Views Grashey & axillary & outlet:Finding:Point in time:Shoulder.left:Document:XR
C1525561|Should-L XR Grashey+Outlet+Serendipity
C1525561|Shoulder - left X-ray Grashey and outlet and Serendipity
C1525561|Views Grashey & outlet & Serendipity:Finding:Point in time:Shoulder.left:Document:XR
C1525561|Views Grashey & outlet & Serendipity:Find:Pt:Shoulder.left:Doc:XR
C1525568|Hip - left X-ray portable
C1525568|Hip-L XR port
C1525568|Views portable:Find:Pt:Hip.left:Doc:XR
C1525568|Views portable:Finding:Point in time:Hip.left:Document:XR
C1525594|Esoph XR W contr PO
C1525594|Esophagus X-ray W contrast PO
C1525594|Views^W contrast PO:Find:Pt:Esophagus:Doc:XR
C1525594|Views^W contrast Oral:Finding:Point in time:Esophagus:Document:XR
C1525685|SC joint-L XR
C1525685|Sternoclavicular joint - left X-ray
C1525685|Views:Find:Pt:Sternoclavicular joint.left:Doc:XR
C1525685|Views:Finding:Point in time:Sternoclavicular joint.left:Document:XR
C1525735|Azygos v XRA W contr IV
C1525735|Azygos vein Fluoroscopic angiogram W contrast IV
C1525735|Views^W contrast IV:Find:Pt:Azygos vein:Doc:XR.fluor.angio
C1525735|Views^W contrast Intravenous:Finding:Point in time:Azygos vein:Document:XR.fluor.angio
C1525770|Wrist - left CT WO contrast
C1525770|Wrist-L CT WO contr
C1525770|Multisection^WO contrast:Finding:Point in time:Wrist.left:Document:Computerized Tomography
C1525770|Multisection^WO contrast:Find:Pt:Wrist.left:Doc:CT
C1525772|Wrist - right CT WO contrast
C1525772|Wrist-R CT WO contr
C1525772|Multisection^WO contrast:Find:Pt:Wrist.right:Doc:CT
C1525772|Multisection^WO contrast:Finding:Point in time:Wrist.right:Document:Computerized Tomography
C1525782|Ankle-L XR Mortise W Stress
C1525782|Ankle - left X-ray Mortise W manual stress
C1525782|View Mortise^W manual stress:Find:Pt:Ankle.left:Doc:XR
C1525782|View Mortise^W manual stress:Finding:Point in time:Ankle.left:Document:XR
C1525792|UE aa-L XRA W contr IA
C1525792|Upper extremity arteries - left Fluoroscopic angiogram W contrast IA
C1525792|Views^W contrast IA:Find:Pt:Upper extremity arteries.left:Doc:XR.fluor.angio
C1525792|Views^W contrast Intra-arterial:Finding:Point in time:Upper extremity arteries.left:Document:XR.fluor.angio
C1525842|TMJ-Bl XR Open+Closed Mouth
C1525842|Temporomandibular joint - bilateral X-ray open and closed mouth
C1525842|Views open & closed mouth:Find:Pt:Temporomandibular joint.bilateral:Doc:XR
C1525842|Views open & closed mouth:Finding:Point in time:Temporomandibular joint.bilateral:Document:XR
C1525864|XXX Flr W contr via Fistula
C1525864|Unspecified body region Fluoroscopy W contrast via fistula
C1525864|Views^W contrast via fistula:Find:Pt:XXX:Doc:XR.fluor
C1525864|Views^W contrast via fistula:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1525870|LE ves XRA W contr IV
C1525870|Lower extremity vessels Fluoroscopic angiogram W contrast IV
C1525870|Views^W contrast Intravenous:Finding:Point in time:Lower extremity vessels:Document:XR.fluor.angio
C1525870|Views^W contrast IV:Find:Pt:Lower extremity vessels:Doc:XR.fluor.angio
C1525883|Ac arch+Carot a-Bl+VA-Bl XRA W contr IA
C1525883|Aortic arch and Carotid artery - bilateral and Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA
C1525883|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery.bilateral+Vertebral artery.bilateral:Document:XR.fluor.angio
C1525883|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery.bilateral+Vertebral artery.bilateral:Doc:XR.fluor.angio
C1525944|Pelvis XR Lat Frog
C1525944|Pelvis X-ray lateral frog
C1525944|View lateral frog:Finding:Point in time:Pelvis:Document:XR
C1525944|View lateral frog:Find:Pt:Pelvis:Doc:XR
C1525825|Finger second - left X-ray
C1525825|Finger.2nd-L XR
C1525825|Views:Finding:Point in time:Finger.second.left:Document:XR
C1525825|Views:Find:Pt:Finger.second.left:Doc:XR
C1525831|Great toe-L XR
C1525831|Great toe - left X-ray
C1525831|Views:Finding:Point in time:Great toe.left:Document:XR
C1525831|Views:Find:Pt:Great toe.left:Doc:XR
C1525835|Breast Mammogram grid
C1525835|Brst Mam Grid
C1525835|Views grid:Finding:Point in time:Breast:Document:Mam
C1525835|Views grid:Find:Pt:Breast:Doc:Mam
C1525953|Acetabulum X-ray 3 views
C1525953|Acetabulum XR 3V
C1525953|Views 3:Find:Pt:Acetabulum:Doc:XR
C1525953|Views 3:Finding:Point in time:Acetabulum:Document:XR
C1525967|SIJ XR Ferguson
C1525967|Sacroiliac Joint X-ray Ferguson
C1525967|View Ferguson:Finding:Point in time:Sacroiliac joint:Document:XR
C1525967|View Ferguson:Find:Pt:Sacroiliac joint:Doc:XR
C1525992|Ankle-R XR stand
C1525992|Ankle - right X-ray standing
C1525992|Views^standing:Find:Pt:Ankle.right:Doc:XR
C1525992|Views^standing:Finding:Point in time:Ankle.right:Document:XR
C1526018|Ft-R XR AP+Lat+Obl
C1526018|Foot - right X-ray AP and lateral and oblique
C1526018|Views AP & lateral & oblique:Finding:Point in time:Foot.right:Document:XR
C1526018|Views AP & lateral & oblique:Find:Pt:Foot.right:Doc:XR
C1526131|Wrist-R XR 2V
C1526131|Wrist - right X-ray 2 views
C1526131|Views 2:Finding:Point in time:Wrist.right:Document:XR
C1526131|Views 2:Find:Pt:Wrist.right:Doc:XR
C1525906|Wrist-R XR PA+Lat+Obl
C1525906|Wrist - right X-ray PA and lateral and oblique
C1525906|Views PA & lateral & oblique:Finding:Point in time:Wrist.right:Document:XR
C1525906|Views PA & lateral & oblique:Find:Pt:Wrist.right:Doc:XR
C1525907|Deprecated Wrist Right X-ray 3 views
C1525907|Views 3:Find:Pt:Wrist.right:Nar:XR
C1525907|Deprecated Wrist-R XR 3V
C1525907|Views 3:Finding:Point in time:Wrist.right:Narrative:XR
C1525907|deprecated VIEWS 3:FINDING:POINT IN TIME:WRIST.RIGHT:NARRATIVE:XR
C1526051|Hip-R XRTomo
C1526051|Hip - right X-ray tomograph
C1526051|Multisection:Find:Pt:Hip.right:Doc:XR.tomo
C1526051|Multisection:Finding:Point in time:Hip.right:Document:XR.tomo
C1525131|Ribs - right X-ray 3 views
C1525131|Ribs-R XR 3V
C1525131|Views 3:Finding:Point in time:Ribs.right:Document:XR
C1525131|Views 3:Find:Pt:Ribs.right:Doc:XR
C1526104|Should-R XR AP+West Point+Outlet
C1526104|Shoulder - right X-ray AP and West Point and outlet
C1526104|Views AP & West Point & outlet:Find:Pt:Shoulder.right:Doc:XR
C1526104|Views AP & West Point & outlet:Finding:Point in time:Shoulder.right:Document:XR
C1524271|SC joint XR 4V
C1524271|Sternoclavicular Joint X-ray 4 views
C1524271|Views 4:Find:Pt:Sternoclavicular joint:Doc:XR
C1524271|Views 4:Finding:Point in time:Sternoclavicular joint:Document:XR
C1526194|US Guidance for biopsy of Breast
C1526194|Brst US Bx guid
C1526194|Guidance for biopsy:Finding:Point in time:Breast:Document:Ultrasound
C1526194|Guidance for biopsy:Find:Pt:Breast:Doc:US
C1526195|Chest US Bx guid
C1526195|US Guidance for biopsy of Chest
C1526195|Guidance for biopsy:Find:Pt:Chest:Doc:US
C1526195|Guidance for biopsy:Finding:Point in time:Chest:Document:Ultrasound
C1526212|Views^W contrast Intrasynovial:Finding:Point in time:Ankle.right:Document:XR.fluor
C1526212|Ankle-R Flr W contr IS
C1526212|Ankle - right Fluoroscopy W contrast IS
C1526212|Views^W contrast IS:Find:Pt:Ankle.right:Doc:XR.fluor
C1526227|Ribs Ant+Post-R XR
C1526227|Ribs anterior and posterior - right X-ray
C1526227|Views:Find:Pt:Ribs.anterior+posterior.right:Doc:XR
C1526227|Views:Finding:Point in time:Ribs.anterior+posterior.right:Document:XR
C1526237|SM v XRA W contr IV
C1526237|Superior mesenteric vein Fluoroscopic angiogram W contrast IV
C1526237|Views^W contrast IV:Find:Pt:Superior mesenteric vein:Doc:XR.fluor.angio
C1526237|Views^W contrast Intravenous:Finding:Point in time:Superior mesenteric vein:Document:XR.fluor.angio
C1526248|Views Broden:Find:Pt:Calcaneus:Doc:XR
C1526248|Deprecated Heel XR Broden
C1526248|Deprecated Calcaneus X-ray Broden
C1526248|Views Broden:Finding:Point in time:Calcaneus:Document:XR
C1524713|Femur - left US
C1524713|Femur-L US
C1524713|Multisection:Finding:Point in time:Femur.left:Document:Ultrasound
C1524713|Multisection:Find:Pt:Femur.left:Doc:US
C1525144|Iliac vessels - right US
C1525144|Iliac ves-R US
C1525144|Multisection:Find:Pt:Iliac vessels.right:Doc:US
C1525144|Multisection:Finding:Point in time:Iliac vessels.right:Document:Ultrasound
C1525150|Finger fifth - right X-ray
C1525150|Finger.5th-R XR
C1525150|Views:Finding:Point in time:Finger.fifth.right:Document:XR
C1525150|Views:Find:Pt:Finger.fifth.right:Doc:XR
C1526322|Spine.epidural space Flr W contr IT
C1526322|Views^W contrast Intrathecal:Finding:Point in time:Spine.epidural space:Document:XR.fluor
C1526322|Views^W contrast IT:Find:Pt:Spine.epidural space:Doc:XR.fluor
C1526322|Spine epidural space Fluoroscopy W contrast IT
C1524481|Ankle-L CT W contr IV
C1524481|Ankle - left CT W contrast IV
C1524481|Multisection^W contrast IV:Find:Pt:Ankle.left:Doc:CT
C1524481|Multisection^W contrast Intravenous:Finding:Point in time:Ankle.left:Document:Computerized Tomography
C1524489|Appendix CT W contr IV
C1524489|Appendix CT W contrast IV
C1524489|Multisection^W contrast IV:Find:Pt:Abdomen+Pelvis>Appendix:Doc:CT
C1524489|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis>Appendix:Document:Computerized Tomography
C1524584|Should CT W contr IV
C1524584|Shoulder CT W contrast IV
C1524584|Multisection^W contrast IV:Find:Pt:Shoulder:Doc:CT
C1524584|Multisection^W contrast Intravenous:Finding:Point in time:Shoulder:Document:Computerized Tomography
C1524306|Fluoroscopy Guidance for biopsy of Spleen
C1524306|Spleen Flr Bx guid
C1524306|Guidance for biopsy:Find:Pt:Spleen:Doc:XR.fluor
C1524306|Guidance for biopsy:Finding:Point in time:Spleen:Document:XR.fluor
C1524594|Lower leg-L CT W contr IV
C1524594|Lower leg - left CT W contrast IV
C1524594|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg.left:Document:Computerized Tomography
C1524594|Multisection^W contrast IV:Find:Pt:Lower leg.left:Doc:CT
C1524601|Multisection^WO & W contrast IV:Find:Pt:Abdomen:Doc:CT
C1524601|Abdomen CT WO and W contrast IV
C1524601|Abd CT WO+W contr IV
C1524601|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524955|Abd XR Obl 1V
C1524955|Abdomen X-ray oblique single view
C1524955|View oblique:Finding:Point in time:Abdomen:Document:XR
C1524955|View oblique:Find:Pt:Abdomen:Doc:XR
C1524959|Finger fourth X-ray oblique single view
C1524959|Finger.4th XR Obl 1V
C1524959|View oblique:Find:Pt:Finger.fourth:Doc:XR
C1524959|View oblique:Finding:Point in time:Finger.fourth:Document:XR
C1526997|Aorta MRI
C1526997|Multisection:Find:Pt:Aorta:Doc:MRI
C1526997|Multisection:Finding:Point in time:Aorta:Document:MRI
C1524630|Finger-L XR 3V
C1524630|Finger - left X-ray 3 views
C1524630|Views 3:Find:Pt:Finger.left:Doc:XR
C1524630|Views 3:Finding:Point in time:Finger.left:Document:XR
C1524648|Elbow - bilateral X-ray 4 views
C1524648|Elbow-Bl XR 4V
C1524648|Views 4:Find:Pt:Elbow.bilateral:Doc:XR
C1524648|Views 4:Finding:Point in time:Elbow.bilateral:Document:XR
C1525013|L-spine XR 2V port
C1525013|Views 2 portable:Find:Pt:Spine.lumbar:Doc:XR
C1525013|Views 2 portable:Finding:Point in time:Spine.lumbar:Document:XR
C1525013|Lumbar spine X-ray 2 views portable
C1525021|Knee - bilateral X-ray 8 views
C1525021|Knee-Bl XR 8V
C1525021|Views 8:Find:Pt:Knee.bilateral:Doc:XR
C1525021|Views 8:Finding:Point in time:Knee.bilateral:Document:XR
C1524352|Internal auditory canal - left CT
C1524352|IAC-L CT
C1524352|Multisection:Find:Pt:Internal auditory canal.left:Doc:CT
C1524352|Multisection:Finding:Point in time:Internal auditory canal.left:Document:Computerized Tomography
C1524358|Elbow - bilateral X-ray tomograph
C1524358|Elbow-Bl XRTomo
C1524358|Multisection:Find:Pt:Elbow.bilateral:Doc:XR.tomo
C1524358|Multisection:Finding:Point in time:Elbow.bilateral:Document:XR.tomo
C1524758|LE.joint-L MRI WO+W contr IV
C1524758|Lower extremity joint - left MRI WO and W contrast IV
C1524758|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.joint.left:Doc:MRI
C1524758|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.joint.left:Document:MRI
C1524759|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.joint.right:Document:MRI
C1524759|LE.joint-R MRI WO+W contr IV
C1524759|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.joint.right:Doc:MRI
C1524759|Lower extremity joint - right MRI WO and W contrast IV
C1524763|Kdny-Bl CT WO+W contr IV
C1524763|Kidney - bilateral CT WO and W contrast IV
C1524763|Multisection^WO & W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:Computerized Tomography
C1524763|Multisection^WO & W contrast IV:Find:Pt:Kidney.bilateral:Doc:CT
C1525030|Elbow-L XR AP+Lat
C1525030|Elbow - left X-ray AP and lateral
C1525030|Views AP & lateral:Finding:Point in time:Elbow.left:Document:XR
C1525030|Views AP & lateral:Find:Pt:Elbow.left:Doc:XR
C1525056|Tib+Fib-Bl XR AP+Lat
C1525056|Tibia - bilateral and Fibula - bilateral X-ray AP and lateral
C1525056|Views AP & lateral:Finding:Point in time:Tibia.bilateral+Fibula.bilateral:Document:XR
C1525056|Views AP & lateral:Find:Pt:Tibia.bilateral+Fibula.bilateral:Doc:XR
C1524416|Upper arm - left CT
C1524416|Upper arm-L CT
C1524416|Multisection:Finding:Point in time:Upper arm.left:Document:Computerized Tomography
C1524416|Multisection:Find:Pt:Upper arm.left:Doc:CT
C1524773|Posterior fossa MRI WO and W contrast IV
C1524773|Multisection^WO & W contrast Intravenous:Finding:Point in time:Posterior fossa:Document:MRI
C1524773|Multisection^WO & W contrast IV:Find:Pt:Posterior fossa:Doc:MRI
C1524773|Post fossa MRI WO+W contr IV
C1830183|US Guidance for aspiration or injection of cyst of Unspecified body region
C1830183|XXX US Asp or Inj of Cyst guid
C1830183|Guidance for aspiration or injection of cyst:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1830183|Guidance for aspiration or injection of cyst:Find:Pt:XXX:Doc:US
C1830229|Head CT W red contr vol IV
C1830229|Head CT W reduced contrast volume IV
C1830229|Multisection^W reduced contrast volume Intravenous:Finding:Point in time:Head:Document:Computerized Tomography
C1830229|Multisection^W reduced contrast volume IV:Find:Pt:Head:Doc:CT
C1830236|Breast - bilateral Mammogram Single view
C1830236|Brst-Bl Mam 1V
C1830236|View 1:Finding:Point in time:Breast.bilateral:Document:Mam
C1830236|View 1:Find:Pt:Breast.bilateral:Doc:Mam
C1830275|Upper extremity vessel graft US.doppler
C1830275|UE ves graft DOP
C1830275|Multisection:Finding:Point in time:Upper extremity vessel graft:Document:Ultrasound.doppler
C1830275|Multisection:Find:Pt:Upper extremity vessel graft:Doc:US.doppler
C1831588|Elbow-Bl XR +Radial Head Capitellar
C1831588|Elbow - bilateral X-ray and radial head capitellar
C1831588|Views & radial head capitellar:Find:Pt:Elbow.bilateral:Doc:XR
C1831588|Views & radial head capitellar:Finding:Point in time:Elbow.bilateral:Document:XR
C1830285|Hrt SPECT Gated Rest+W Tc99mMIBI IV
C1830285|Heart SPECT gated at rest and W Tc-99m Sestamibi IV
C1830285|Multisection gated^at rest & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1830285|Multisection gated^at rest & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1715389|CT Guidance for needle localization of Breast-- WO and W contrast IV
C1715389|Guidance for needle localization^WO & W contrast IV:Find:Pt:Breast:Doc:CT
C1715389|Brst CT Needle local guid WO+W contr IV
C1715389|Guidance for needle localization^WO & W contrast Intravenous:Finding:Point in time:Breast:Document:Computerized Tomography
C1715395|BD+PDs MRI W contr IV
C1715395|Biliary ducts and Pancreatic duct MRI W contrast IV
C1715395|Multisection^W contrast Intravenous:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:MRI
C1715395|Multisection^W contrast IV:Find:Pt:Biliary ducts+Pancreatic duct:Doc:MRI
C1715408|Brain PET
C1715408|Multisection:Find:Pt:Brain:Doc:Radnuc.PET
C1715408|Multisection:Finding:Point in time:Brain:Document:Radnuc.PET
C1645318|Knee-L XR port
C1645318|Knee - left X-ray portable
C1645318|Views portable:Finding:Point in time:Knee.left:Document:XR
C1645318|Views portable:Find:Pt:Knee.left:Doc:XR
C1637277|Hip-L XR AP+Lat+Measure
C1637277|Hip - left X-ray AP and lateral and measurement
C1637277|Views AP & lateral & measurement:Finding:Point in time:Hip.left:Document:XR
C1637277|Views AP & lateral & measurement:Find:Pt:Hip.left:Doc:XR
C1717248|Brain RI During EST
C1717248|Brain Scan during electroconvulsive shock treatment
C1717248|Views^during electroconvulsive shock treatment:Find:Pt:Brain:Doc:Radnuc
C1717248|Views^during electroconvulsive shock treatment:Finding:Point in time:Brain:Document:Radnuc
C1706626|Finger.2nd-L XR GE 3V
C1706626|Finger second - left X-ray GE 3 views
C1706626|Finger second - left Narrative X-ray GE 3 views
C1706626|Views GE 3:Find:Pt:Finger.second.left:Doc:XR
C1706626|Views GE 3:Finding:Point in time:Finger.second.left:Document:XR
C1714921|Pelvis XR 1V or 2V
C1714921|Pelvis X-ray 1 or 2 views
C1714921|Views 1 or 2:Finding:Point in time:Pelvis:Document:XR
C1714921|Views 1 or 2:Find:Pt:Pelvis:Doc:XR
C1706627|Deprecated Finger.2nd-L XR GE 3V
C1706627|Views GE 3:Find:Pt:Finger.second.left:Nar:XR
C1706627|Deprecated Finger second Left X-ray GE 3 views
C1706627|Views GE 3:Finding:Point in time:Finger.second.left:Narrative:XR
C1715122|Wrist - bilateral X-ray tunnel.carpal
C1715122|Wrist-Bl XR Tunnel.carpal
C1715122|Views tunnel.carpal:Finding:Point in time:Wrist.bilateral:Document:XR
C1715122|Views tunnel.carpal:Find:Pt:Wrist.bilateral:Doc:XR
C1638456|Brst-L Mam p wire plac
C1638456|Breast - left Mammogram Post Wire Placement
C1638456|Views^post wire placement:Find:Pt:Breast.left:Doc:Mam
C1638456|Views^post wire placement:Finding:Point in time:Breast.left:Document:Mam
C1635008|Fluoroscopy Guidance for percutaneous drainage of abscess of Unspecified body region
C1635008|XXX Flr PC Abscess Drain guid
C1635008|Guidance for percutaneous drainage of abscess:Find:Pt:XXX:Doc:XR.fluor
C1635008|Guidance for percutaneous drainage of abscess:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1644171|Brst US Bx Excisional guid
C1644171|US Guidance for excisional biopsy of Breast
C1644171|Guidance for biopsy.excisional:Find:Pt:Breast:Doc:US
C1644171|Guidance for biopsy.excisional:Finding:Point in time:Breast:Document:Ultrasound
C1632257|Abd XR AP (Upr+L Lat Decub)
C1632257|Abdomen X-ray AP (upright and left lateral decubitus)
C1632257|Views AP (upright & L-lateral decubitus):Find:Pt:Abdomen:Doc:XR
C1632257|Views AP (upright & L-lateral decubitus):Finding:Point in time:Abdomen:Document:XR
C1626178|Scan whole body
C1626178|RI WB W RNC IV
C1626178|Views whole body^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C1626178|Views whole body^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1631783|Views flow^W radionuclide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1631783|Views flow^W radionuclide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1631783|Kidney - bilateral Scan flow
C1631783|Kdny-Bl RI Flow W RNC IV
C1631259|Guidance for drainage of abscess:Finding:Point in time:Abdomen+Pelvis>Appendix:Document:Computerized Tomography
C1631259|Guidance for drainage of abscess:Find:Pt:Abdomen+Pelvis>Appendix:Doc:CT
C1631259|Appendix CT Abscess drain guid
C1631259|CT Guidance for drainage of abscess of Appendix
C1624696|Clavicle MRI W contr IV
C1624696|Clavicle MRI W contrast IV
C1624696|Multisection^W contrast IV:Find:Pt:Clavicle:Doc:MRI
C1624696|Multisection^W contrast Intravenous:Finding:Point in time:Clavicle:Document:MRI
C2361223|CT Guidance for replacement of percutaneous drainage tube in Abdomen
C2361223|Abd CT Replac of PC drain tube guid
C2361223|Guidance for replacement of percutaneous drainage tube:Find:Pt:Abdomen:Doc:CT
C2361223|Guidance for replacement of percutaneous drainage tube:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1977263|Views:Finding:Point in time:To be specified in another part of the message:Narrative:XR.fluor
C1977263|Unspecified body region Fluoroscopy
C1977263|XXX Flr
C1977263|Views:Find:Pt:XXX:Doc:XR.fluor
C1977263|Views:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1954308|Multisection^WO & W contrast IV:Find:Pt:Brain.temporal:Doc:MRI
C1954308|Brain.temporal MRI WO+W contr IV
C1954308|Brain.temporal MRI WO and W contrast IV
C1954308|Multisection^WO & W contrast Intravenous:Finding:Point in time:Brain.temporal:Document:MRI
C3173624|Renal ves-L XRA W contr
C3173624|Renal vessels - left Fluoroscopic angiogram W contrast
C3173624|Views^W contrast:Find:Pt:Renal vessels.left:Doc:XR.fluor.angio
C3173624|Views^W contrast:Finding:Point in time:Renal vessels.left:Document:XR.fluor.angio
C3262938|Wrist - right CT W contrast IS
C3262938|Multisection^W contrast IS:Find:Pt:Wrist.right:Doc:CT
C3262938|Multisection^W contrast Intrasynovial:Finding:Point in time:Wrist.right:Document:Computerized Tomography
C3262938|Wrist-R CT W contr IS
C3262969|Breast implant - left Mammogram diagnostic
C3262969|Brst implant-L Mam Dx
C3262969|Views diagnostic:Finding:Point in time:Breast implant.left:Document:Mam
C3262969|Views diagnostic:Find:Pt:Breast implant.left:Doc:Mam
C3263008|UE-Bl MRI WO contr
C3263008|Upper extremity - bilateral MRI WO contrast
C3263008|Multisection^WO contrast:Finding:Point in time:Upper extremity.bilateral:Document:MRI
C3263008|Multisection^WO contrast:Find:Pt:Upper extremity.bilateral:Doc:MRI
C3482438|C-spine Flr PC Vertebroplasty guid
C3482438|Guidance for percutaneous vertebroplasty:Find:Pt:Spine.cervical:Doc:XR.fluor
C3482438|Guidance for percutaneous vertebroplasty:Finding:Point in time:Spine.cervical:Document:XR.fluor
C3482438|Fluoroscopy Guidance for percutaneous vertebroplasty of Cervical spine
C3263021|Should-L MRI WO+W contr IS
C3263021|Multisection^WO & W contrast Intrasynovial:Finding:Point in time:Shoulder.left:Document:MRI
C3263021|Multisection^WO & W contrast IS:Find:Pt:Shoulder.left:Doc:MRI
C3263021|Shoulder - left MRI WO and W contrast IS
C3263045|Heart Scan W stress and W Tc-99m Sestamibi IV
C3263045|Hrt RI W Stress+W Tc99mMIBI IV
C3263045|Views^W stress & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C3263045|Views^W stress & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C3263063|Portal v XRA W contr IV
C3263063|Portal vein Fluoroscopic angiogram W contrast IV
C3263063|Views^W contrast Intravenous:Finding:Point in time:Portal vein:Document:XR.fluor.angio
C3263063|Views^W contrast IV:Find:Pt:Portal vein:Doc:XR.fluor.angio
C3263068|Knee - right X-ray Sunrise and tunnel standing
C3263068|Knee-R XR Sunrise+Tunnel stand
C3263068|Views Sunrise & tunnel^standing:Find:Pt:Knee.right:Doc:XR
C3263068|Views Sunrise & tunnel^standing:Finding:Point in time:Knee.right:Document:XR
C3263075|Wrist - right X-ray PA W clenched fist
C3263075|Wrist-R XR PA V1 W clenched fist
C3263075|View PA^W clenched fist:Find:Pt:Wrist.right:Doc:XR
C3263075|View PA^W clenched fist:Finding:Point in time:Wrist.right:Document:XR
C3263077|Shoulder X-ray 4 views
C3263077|Should XR 4V
C3263077|Views 4:Finding:Point in time:Shoulder:Document:XR
C3263077|Views 4:Find:Pt:Shoulder:Doc:XR
C3263204|Urinary bladder US post void
C3263204|Bladder US p vdg
C3263204|Multisection^post void:Finding:Point in time:Urinary bladder:Document:Ultrasound
C3263204|Multisection^post void:Find:Pt:Urinary bladder:Doc:US
C3262880|Acromioclavicular joint - bilateral X-ray WO weight
C3262880|AC joint-Bl XR WO Wt
C3262880|Views^WO weight:Find:Pt:Acromioclavicular joint.bilateral:Doc:XR
C3262880|Views^WO weight:Finding:Point in time:Acromioclavicular joint.bilateral:Document:XR
C3262890|XXX XRA Angpsty W contr
C3262890|Unspecified body region Fluoroscopic angiogram Angioplasty W contrast
C3262890|Angioplasty^W contrast:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor.angio
C3262890|Angioplasty^W contrast:Find:Pt:XXX:Doc:XR.fluor.angio
C3262905|Deprecated Head CT and 3D reconstruction WO contrast
C3262905|Multisection & 3D reconstruction^WO contrast:Finding:Point in time:Head:Document:Computerized Tomography
C3262905|Multisection & 3D reconstruction^WO contrast:Find:Pt:Head:Doc:CT
C3262905|Deprecated Head CT +3DR WO contr
C3262919|Chest CT limited W contrast IV
C3262919|Chest CT Ltd W contr IV
C3262919|Multisection limited^W contrast Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C3262919|Multisection limited^W contrast IV:Find:Pt:Chest:Doc:CT
C2709250|Views:Finding:Point in time:Skull:Narrative:XR
C2709250|Skull X-ray
C2709250|Skull XR
C2709250|Views:Find:Pt:Skull:Doc:XR
C2709250|Views:Finding:Point in time:Skull:Document:XR
C0942189|TO ves-R MRI.Angio W contr IV
C0942189|Thoracic outlet vessels - right MRI angiogram W contrast IV
C0942189|Multisection^W contrast Intravenous:Finding:Point in time:Thoracic outlet vessels.right:Document:MRI.angio
C0942189|Multisection^W contrast IV:Find:Pt:Thoracic outlet vessels.right:Doc:MRI.angio
C0945329|Hand - right MRI
C0945329|Hand-R MRI
C0945329|Multisection:Finding:Point in time:Hand.right:Document:MRI
C0945329|Multisection:Find:Pt:Hand.right:Doc:MRI
C0942304|Mammogram Guidance for needle localization of mass of Breast - right
C0942304|Brst-R Mam Needle local mass guid
C0942304|Guidance for needle localization of mass:Find:Pt:Breast.right:Doc:Mam
C0942304|Guidance for needle localization of mass:Finding:Point in time:Breast.right:Document:Mam
C0942323|Mammogram Guidance for biopsy of Breast - bilateral
C0942323|Brst-Bl Mam Bx guid
C0942323|Guidance for biopsy:Finding:Point in time:Breast.bilateral:Document:Mam
C0942323|Guidance for biopsy:Find:Pt:Breast.bilateral:Doc:Mam
C0942346|Knee-R XR AP+Lat stand
C0942346|Knee - right X-ray AP and lateral standing
C0942346|Views AP & lateral^standing:Finding:Point in time:Knee.right:Document:XR
C0942346|Views AP & lateral^standing:Find:Pt:Knee.right:Doc:XR
C0945348|Patella - left X-ray 2 views
C0945348|Patella-L XR 2V
C0945348|Views 2:Find:Pt:Patella.left:Doc:XR
C0945348|Views 2:Finding:Point in time:Patella.left:Document:XR
C0882206|Multisectional sagittal:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882206|Deprecated Unspecified body region CT Multisectional sagittal
C0882206|Multisectional sagittal:Find:Pt:XXX:Doc:CT
C0882206|Deprecated XXX CT Multisectional sagitta
C0945307|Views^W contrast IS:Find:Pt:Shoulder.right:Doc:XR.fluor
C0945307|Should-R Flr W contr IS
C0945307|Shoulder - right Fluoroscopy W contrast IS
C0945307|Views^W contrast Intrasynovial:Finding:Point in time:Shoulder.right:Document:XR.fluor
C0942107|Knee-L XR stand
C0942107|Knee - left X-ray standing
C0942107|Views^standing:Finding:Point in time:Knee.left:Document:XR
C0942107|Views^standing:Find:Pt:Knee.left:Doc:XR
C0942115|Ft-L XR stand
C0942115|Foot - left X-ray standing
C0942115|Views^standing:Find:Pt:Foot.left:Doc:XR
C0942115|Views^standing:Finding:Point in time:Foot.left:Document:XR
C0942122|Deprecated Heel-R XR
C0942122|Deprecated Calcaneus - right X-ray
C0942122|Views:Find:Pt:Calcaneus.right:Doc:XR
C0942122|Views:Finding:Point in time:Calcaneus.right:Document:XR
C0945311|UE-L XR
C0945311|Upper extremity - left X-ray
C0945311|Views:Finding:Point in time:Upper extremity.left:Document:XR
C0945311|Views:Find:Pt:Upper extremity.left:Doc:XR
C0881793|Artery Fluoroscopic angiogram Embolization W contrast IA
C0881793|Artery XRA Embolization W contr IA
C0881793|Embolization^W contrast Intra-arterial:Finding:Point in time:To be specified in another part of the message artery:Document:XR.fluor.angio
C0881793|Embolization^W contrast IA:Find:Pt:XXX artery:Doc:XR.fluor.angio
C0882520|Head ves MRI.Angio W contr IV
C0882520|Head vessels MRI angiogram W contrast IV
C0882520|Multisection^W contrast Intravenous:Finding:Point in time:Head vessels:Document:MRI.angio
C0882520|Multisection^W contrast IV:Find:Pt:Head vessels:Doc:MRI.angio
C0882522|Guidance for nerve block:Finding:Point in time:Chest>Celiac plexus:Document:Computerized Tomography
C0882522|Guidance for nerve block:Find:Pt:Chest>Celiac plexus:Doc:CT
C0882522|Celiac plexus CT Nerve Block guid
C0882522|CT Guidance for nerve block of Celiac plexus
C0881880|Chest XR AP+AP R-Lat Debuc Port
C0881880|Chest X-ray AP and AP right lateral-decubitus portable
C0881880|Views AP & AP R-lateral-decubitus portable:Find:Pt:Chest:Doc:XR
C0881880|Views AP & AP R-lateral-decubitus portable:Finding:Point in time:Chest:Document:XR
C0881885|TA MRI.Angio
C0881885|Aorta thoracic MRI angiogram
C0881885|Multisection:Find:Pt:Aorta.thoracic:Doc:MRI.angio
C0881885|Multisection:Finding:Point in time:Aorta.thoracic:Document:MRI.angio
C0881951|Head ves DOP
C0881951|Head vessels US.doppler
C0881951|Multisection:Find:Pt:Head vessels:Doc:US.doppler
C0881951|Multisection:Finding:Point in time:Head vessels:Document:Ultrasound.doppler
C0881974|Views^W radionuclide transplant scan:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C0881974|Kidney - bilateral Scan W radionuclide transplant scan
C0881974|Views^W radionuclide transplant scan:Find:Pt:Kidney.bilateral:Doc:Radnuc
C0881974|Kdny-Bl RI W RNC Transplant Scan
C0881984|Multisection^W & WO contrast Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:XR.tomo
C0881984|Multisection^WO & W contrast IV:Find:Pt:Kidney.bilateral:Doc:XR.tomo
C0881984|Multisection^WO & W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:XR.tomo
C0881984|Kdny-Bl XRTomo WO+W contr IV
C0881984|Kidney - bilateral X-ray tomograph WO and W contrast IV
C0881999|View AP:Finding:Point in time:Abdomen:Narrative:XR
C0881999|Abdomen X-ray AP single view
C0881999|Abd XR AP 1V
C0881999|View AP:Find:Pt:Abdomen:Doc:XR
C0881999|View AP:Finding:Point in time:Abdomen:Document:XR
C0882011|Liver CT Bx CN guid
C0882011|CT Guidance for core needle biopsy of Liver
C0882011|Guidance for biopsy.core needle:Find:Pt:Abdomen>Liver:Doc:CT
C0882011|Guidance for biopsy.core needle:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1114482|Neck MRI WO contrast
C1114482|Neck MRI WO contr
C1114482|Multisection^WO contrast:Finding:Point in time:Neck:Document:MRI
C1114482|Multisection^WO contrast:Find:Pt:Neck:Doc:MRI
C1114513|Thyroid Scan
C1114513|Thyroid RI W RNC IV
C1114513|Views^W radionuclide IV:Find:Pt:Thyroid:Doc:Radnuc
C1114513|Views^W radionuclide Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1114513|VIEWS^RADIONUCLIDE.INTRAVENOUS:FINDING:POINT IN TIME:THYROID:NARRATIVE:RADNUC
C1114550|Chest X-ray left lateral
C1114550|Chest XR L-Lat
C1114550|View L-lateral:Find:Pt:Chest:Doc:XR
C1114550|View L-lateral:Finding:Point in time:Chest:Document:XR
C1114610|LE-ves CT.Angio WO+W contr IV
C1114610|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity>Vessels:Document:Computerized Tomography.angio
C1114610|Lower extremity Vessels CT angiogram WO and W contrast IV
C1114610|Multisection^WO & W contrast IV:Find:Pt:Lower extremity>Vessels:Doc:CT.angio
C1114626|SS v+Jugular v XRA W contr IV
C1114626|Sagittal sinus and Jugular veins Fluoroscopic angiogram W contrast IV
C1114626|Views^W contrast IV:Find:Pt:Sagittal sinus vein+Jugular vein:Doc:XR.fluor.angio
C1114626|Views^W contrast Intravenous:Finding:Point in time:Sagittal sinus vein+Jugular vein:Document:XR.fluor.angio
C1114922|IAC CT W contr IV
C1114922|Internal auditory canal CT W contrast IV
C1114922|Multisection^W contrast IV:Find:Pt:Internal auditory canal:Doc:CT
C1114922|Multisection^W contrast Intravenous:Finding:Point in time:Internal auditory canal:Document:Computerized Tomography
C1526823|Ribs upper - left X-ray
C1526823|Ribs upper-L XR
C1526823|Views:Find:Pt:Ribs.upper.left:Doc:XR
C1526823|Views:Finding:Point in time:Ribs.upper.left:Document:XR
C1543458|Ft-R XR AP+Lat+Obl stand
C1543458|Foot - right X-ray AP and lateral and oblique standing
C1543458|Views AP & lateral & oblique^standing:Finding:Point in time:Foot.right:Document:XR
C1543458|Views AP & lateral & oblique^standing:Find:Pt:Foot.right:Doc:XR
C1543746|Liver transplant Scan
C1543746|Liver Transplant RI W RNC IV
C1543746|Views^W radionuclide Intravenous:Finding:Point in time:Liver transplant:Document:Radnuc
C1543746|Views^W radionuclide IV:Find:Pt:Liver transplant:Doc:Radnuc
C1543748|Lung RI W Depreotide+RNC IV
C1543748|Lung Scan W depreotide and W radionuclide IV
C1543748|Views^W depreotide & W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1543748|Views^W depreotide & W radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1543761|Hrt RI PF W DIPY+Tc99mIV
C1543761|Heart Scan perfusion W dipyridamole and W Tc-99m IV
C1543761|Views perfusion^W dipyridamole & W Tc-99m Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543761|Views perfusion^W dipyridamole & W Tc-99m IV:Find:Pt:Heart:Doc:Radnuc
C1543471|Shoulder - right X-ray 3 views and axillary
C1543471|Should-R XR 3V+Ax
C1543471|Views 3 & axillary:Finding:Point in time:Shoulder.right:Document:XR
C1543471|Views 3 & axillary:Find:Pt:Shoulder.right:Doc:XR
C1543483|Sternum XR Lat+R-ant Obl
C1543483|Sternum X-ray lateral and right anterior oblique
C1543483|Views lateral & R-anterior oblique:Find:Pt:Sternum:Doc:XR
C1543483|Views lateral & R-anterior oblique:Finding:Point in time:Sternum:Document:XR
C1543801|RI for Tumor WB W Tc99mMIBI IV
C1543801|Scan for tumor whole body W Tc-99m Sestamibi IV
C1543801|Views for tumor whole body^W Tc-99m Sestamibi Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543801|Views for tumor whole body^W Tc-99m Sestamibi IV:Find:Pt:^Patient:Doc:Radnuc
C1543895|Hrt RI WM W RNC IV
C1543895|Heart Scan wall motion
C1543895|Views wall motion^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543895|Views wall motion^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543931|Hrt RI FP+WM+VV+EF W Stress+W RNC IV
C1543931|Heart Scan first pass and wall motion and ventricular volume and ejection fraction W stress and W radionuclide IV
C1543931|Views first pass & wall motion & ventricular volume & ejection fraction^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543931|Views first pass & wall motion & ventricular volume & ejection fraction^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543947|Hrt RI Gated+WM+EF Rest+W RNC IV
C1543947|Heart Scan gated and wall motion and ejection fraction at rest and W radionuclide IV
C1543947|Views gated & wall motion & ejection fraction^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543947|Views gated & wall motion & ejection fraction^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543949|Hrt RI Gated W Stress+W Tc99mP IV
C1543949|Heart Scan gated W stress and W Tc-99m pertechnetate IV
C1543949|Views gated^W stress & W Tc-99m pertechnetate Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543949|Views gated^W stress & W Tc-99m pertechnetate IV:Find:Pt:Heart:Doc:Radnuc
C1543959|Lung RI VP+Diff W RNC IH+IV
C1543959|Views ventilation & perfusion & differential^W radionuclide Inhalation & W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1543959|Views ventilation & perfusion & differential^W radionuclide IH & W radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1543959|Lung Scan ventilation and perfusion and differential W radionuclide IH and W radionuclide IV
C1543500|Extremity vessels US.doppler limited
C1543500|Extr ves DOP Ltd
C1543500|Multisection limited:Finding:Point in time:Extremity vessels:Document:Ultrasound.doppler
C1543500|Multisection limited:Find:Pt:Extremity vessels:Doc:US.doppler
C1543504|Extremity artery - left US.doppler
C1543504|Extr a-L DOP
C1543504|Multisection:Finding:Point in time:Extremity artery.left:Document:Ultrasound.doppler
C1543504|Multisection:Find:Pt:Extremity artery.left:Doc:US.doppler
C1543507|LE ves-L DOP
C1543507|Lower extremity vessels - left US.doppler
C1543507|Multisection:Finding:Point in time:Lower extremity vessels.left:Document:Ultrasound.doppler
C1543507|Multisection:Find:Pt:Lower extremity vessels.left:Doc:US.doppler
C1543521|Vessels US.doppler
C1543521|Vesl DOP
C1543521|Multisection:Find:Pt:Vessels:Doc:US.doppler
C1543521|Multisection:Finding:Point in time:Vessels:Document:Ultrasound.doppler
C1543160|Multisection:Finding:Point in time:Brachiocephalic artery:Narrative:ULTRASOUND.doppler
C1543160|BrachCeph a DOP
C1543160|Brachiocephalic artery US.doppler
C1543160|Multisection:Finding:Point in time:Brachiocephalic artery:Document:Ultrasound.doppler
C1543160|Multisection:Find:Pt:Brachiocephalic artery:Doc:US.doppler
C1543176|Extr vv XRA W contr IV
C1543176|Extremity veins Fluoroscopic angiogram W contrast IV
C1543176|Views^W contrast Intravenous:Finding:Point in time:Extremity veins:Document:XR.fluor.angio
C1543176|Views^W contrast IV:Find:Pt:Extremity veins:Doc:XR.fluor.angio
C1543186|Pelvis XR AP+Inlet+Outlet+Obl
C1543186|Pelvis X-ray AP and inlet and outlet and oblique
C1543186|Views AP & inlet & outlet & oblique:Find:Pt:Pelvis:Doc:XR
C1543186|Views AP & inlet & outlet & oblique:Finding:Point in time:Pelvis:Document:XR
C1525930|Elbow-R XR Jones
C1525930|Elbow - right X-ray Jones
C1525930|View Jones:Find:Pt:Elbow.right:Doc:XR
C1525930|View Jones:Finding:Point in time:Elbow.right:Document:XR
C1542865|Breast - bilateral FFD mammogram diagnostic
C1542865|Brst-Bl FFDM Dx
C1542865|Views diagnostic:Finding:Point in time:Breast.bilateral:Document:Mam.FFD
C1542865|Views diagnostic:Find:Pt:Breast.bilateral:Doc:Mam.FFD
C1543717|Hrt SPECT for Infarct W Tc99mMIBI IV
C1543717|Heart SPECT for infarct W Tc-99m Sestamibi IV
C1543717|Multisection for infarct^W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543717|Multisection for infarct^W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543721|Views^at rest & W 201 TI IV:Find:Pt:Heart:Nar:Radnuc
C1543721|Deprecated Heart Scintigraphy at rest & W Tl-201 IV
C1543721|Deprecated Hrt RI
C1543721|Views^at rest & W 201 TI Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1543721|Deprecated Hrt RI At Rest+W 201 TI IV
C1526799|Wrist - left X-ray 2 views tunnel.carpal
C1526799|Wrist-L XR 2V Tunnel
C1526799|Views 2 tunnel.carpal:Finding:Point in time:Wrist.left:Document:XR
C1526799|Views 2 tunnel.carpal:Find:Pt:Wrist.left:Doc:XR
C1526805|Lower extremity - left X-ray AP single view standing
C1526805|LE-L XR AP 1V stand
C1526805|View AP^standing:Finding:Point in time:Lower extremity.left:Document:XR
C1526805|View AP^standing:Find:Pt:Lower extremity.left:Doc:XR
C1524429|Knee-L XRTomo
C1524429|Knee - left X-ray tomograph
C1524429|Multisection:Finding:Point in time:Knee.left:Document:XR.tomo
C1524429|Multisection:Find:Pt:Knee.left:Doc:XR.tomo
C1527067|Parathyroid MRI
C1527067|Multisection:Finding:Point in time:Parathyroid:Document:MRI
C1527067|Multisection:Find:Pt:Parathyroid:Doc:MRI
C1524194|IVC MRI.Angio
C1524194|Inferior vena cava MRI angiogram
C1524194|Multisection:Finding:Point in time:Vena cava.inferior:Document:MRI.angio
C1524194|Multisection:Find:Pt:Vena cava.inferior:Doc:MRI.angio
C1524825|Multisection^WO contrast:Find:Pt:Calcaneus.left:Doc:CT
C1524825|Multisection^WO contrast:Finding:Point in time:Calcaneus.left:Document:Computerized Tomography
C1524825|Deprecated Calcaneus - left CT WO contrast
C1524825|Deprecated Heel-L CT WO contr
C1525120|Extr ves MRI.Angio
C1525120|Extremity vessels MRI angiogram
C1525120|Multisection:Finding:Point in time:Extremity vessels:Document:MRI.angio
C1525120|Multisection:Find:Pt:Extremity vessels:Doc:MRI.angio
C1525316|Abd XR Lat Xtable
C1525316|Abdomen X-ray lateral crosstable
C1525316|View lateral crosstable:Find:Pt:Abdomen:Doc:XR
C1525316|View lateral crosstable:Finding:Point in time:Abdomen:Document:XR
C1525324|L-spine XR Lat Xtable port
C1525324|View lateral crosstable portable:Find:Pt:Spine.lumbar:Doc:XR
C1525324|View lateral crosstable portable:Finding:Point in time:Spine.lumbar:Document:XR
C1525324|Lumbar spine X-ray lateral crosstable portable
C1525190|Multisection^W contrast IV:Find:Pt:Head>Arteries:Doc:CT.angio
C1525190|Multisection^W contrast Intravenous:Finding:Point in time:Head>Arteries:Document:Computerized Tomography.angio
C1525190|Head Arteries CT angiogram W contrast IV
C1525190|Head Arteries CT.Angio W contr IV
C1525239|Shoulder vessels - right MRI angiogram WO and W contrast IV
C1525239|Multisection^WO & W contrast IV:Find:Pt:Shoulder vessels.right:Doc:MRI.angio
C1525239|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder vessels.right:Document:MRI.angio
C1525239|Should ves-R MRI.Angio WO+W contr IV
C1525269|Maxillofacial region CT limited
C1525269|Maxillofacial CT Ltd
C1525269|Multisection limited:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1525269|Multisection limited:Find:Pt:Head>Maxillofacial region:Doc:CT
C1525326|Hip - left X-ray lateral frog
C1525326|Hip-L XR Lat Frog
C1525326|View lateral frog:Finding:Point in time:Hip.left:Document:XR
C1525326|View lateral frog:Find:Pt:Hip.left:Doc:XR
C1524683|Abdomen X-ray PA prone
C1524683|Abd XR PA Prone
C1524683|View PA prone:Find:Pt:Abdomen:Doc:XR
C1524683|View PA prone:Finding:Point in time:Abdomen:Document:XR
C1525465|Hip X-ray true lateral
C1525465|Hip XR True Lat
C1525465|View true lateral:Find:Pt:Hip:Doc:XR
C1525465|View true lateral:Finding:Point in time:Hip:Document:XR
C1525466|Hip - left X-ray true lateral
C1525466|Hip-L XR True Lat
C1525466|View true lateral:Finding:Point in time:Hip.left:Document:XR
C1525466|View true lateral:Find:Pt:Hip.left:Doc:XR
C1524222|Shoulder - bilateral X-ray Velpeau axillary
C1524222|Should-Bl XR Velpeau Ax
C1524222|View Velpeau axillary:Find:Pt:Shoulder.bilateral:Doc:XR
C1524222|View Velpeau axillary:Finding:Point in time:Shoulder.bilateral:Document:XR
C1524230|Scapula - bilateral X-ray Y
C1524230|Scapula-Bl XR Y
C1524230|View Y:Find:Pt:Scapula.bilateral:Doc:XR
C1524230|View Y:Finding:Point in time:Scapula.bilateral:Document:XR
C1525494|Should-L XR AP+Ax+Outlet+Zanca
C1525494|Shoulder - left X-ray AP and axillary and outlet and Zanca
C1525494|Views AP & axillary & outlet & Zanca:Find:Pt:Shoulder.left:Doc:XR
C1525494|Views AP & axillary & outlet & Zanca:Finding:Point in time:Shoulder.left:Document:XR
C1525516|Knee-Bl XR AP+Lat+Sunrise+Tunnel
C1525516|Knee - bilateral X-ray AP and lateral and Sunrise and tunnel
C1525516|Views AP & lateral & Sunrise & tunnel:Find:Pt:Knee.bilateral:Doc:XR
C1525516|Views AP & lateral & Sunrise & tunnel:Finding:Point in time:Knee.bilateral:Document:XR
C1525530|Abd XR R-Lat+L-Lat
C1525530|Abdomen X-ray right lateral and left lateral
C1525530|Views R-lateral & L-lateral:Find:Pt:Abdomen:Doc:XR
C1525530|Views R-lateral & L-lateral:Finding:Point in time:Abdomen:Document:XR
C1525578|Popliteal artery - left Fluoroscopic angiogram W contrast IA
C1525578|Popliteal a-L XRA W contr IA
C1525578|Views^W contrast Intra-arterial:Finding:Point in time:Popliteal artery.left:Document:XR.fluor.angio
C1525578|Views^W contrast IA:Find:Pt:Popliteal artery.left:Doc:XR.fluor.angio
C1525607|CT Guidance for biopsy of Bone marrow
C1525607|BM CT Bx guid
C1525607|Guidance for biopsy:Find:Pt:Bone marrow:Doc:CT
C1525607|Guidance for biopsy:Finding:Point in time:Bone marrow:Document:Computerized Tomography
C1525615|Biliary ducts MRI
C1525615|BDs MRI
C1525615|Multisection:Finding:Point in time:Biliary ducts:Document:MRI
C1525615|Multisection:Find:Pt:Biliary ducts:Doc:MRI
C1525644|Soft tissue MRI W contr IV
C1525644|Soft tissue MRI W contrast IV
C1525644|Multisection^W contrast IV:Find:Pt:Soft tissue:Doc:MRI
C1525644|Multisection^W contrast Intravenous:Finding:Point in time:Soft tissue:Document:MRI
C1525800|C-spine CT W contr ID
C1525800|Multisection^W contrast intradisc:Find:Pt:Spine.cervical:Doc:CT
C1525800|Multisection^W contrast intradisc:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C1525800|Cervical spine CT W contrast intradisc
C1525818|LS-spine junc XR Lat Spot
C1525818|Spine Lumbosacral Junction X-ray lateral spot
C1525818|View lateral spot:Find:Pt:Spine.lumbosacral junction:Doc:XR
C1525818|View lateral spot:Finding:Point in time:Spine.lumbosacral junction:Document:XR
C1525965|Sacroiliac Joint X-ray 3 views
C1525965|SIJ XR 3V
C1525965|Views 3:Finding:Point in time:Sacroiliac joint:Document:XR
C1525965|Views 3:Find:Pt:Sacroiliac joint:Doc:XR
C1525978|Acromioclavicular joint - right X-ray AP single view
C1525978|AC joint-R XR AP 1V
C1525978|View AP:Find:Pt:Acromioclavicular joint.right:Doc:XR
C1525978|View AP:Finding:Point in time:Acromioclavicular joint.right:Document:XR
C1526007|Femur - right X-ray 4 views
C1526007|Femur-R XR 4V
C1526007|Views 4:Finding:Point in time:Femur.right:Document:XR
C1526007|Views 4:Find:Pt:Femur.right:Doc:XR
C1526113|Sternoclavicular joint - right X-ray Serendipity
C1526113|SC joint-R XR Serendipity
C1526113|View Serendipity:Finding:Point in time:Sternoclavicular joint.right:Document:XR
C1526113|View Serendipity:Find:Pt:Sternoclavicular joint.right:Doc:XR
C1526057|Knee-R XR 1V
C1526057|Knee - right X-ray Single view
C1526057|View 1:Finding:Point in time:Knee.right:Document:XR
C1526057|View 1:Find:Pt:Knee.right:Doc:XR
C1526103|Shoulder - right X-ray AP single view
C1526103|Should-R XR AP 1V
C1526103|View AP:Finding:Point in time:Shoulder.right:Document:XR
C1526103|View AP:Find:Pt:Shoulder.right:Doc:XR
C1526146|Sinuses XR 3V
C1526146|Sinuses X-ray 3 views
C1526146|Views 3:Finding:Point in time:Sinuses:Document:XR
C1526146|Views 3:Find:Pt:Sinuses:Doc:XR
C1526161|Skull XR Lat+Towne
C1526161|Skull X-ray lateral and Towne
C1526161|Views lateral & Towne:Finding:Point in time:Skull:Document:XR
C1526161|Views lateral & Towne:Find:Pt:Skull:Doc:XR
C1526193|Abd US Bx guid
C1526193|US Guidance for biopsy of Abdomen
C1526193|Guidance for biopsy:Find:Pt:Abdomen:Doc:US
C1526193|Guidance for biopsy:Finding:Point in time:Abdomen:Document:Ultrasound
C1526200|Salivary gland US Bx guid
C1526200|US Guidance for biopsy of Salivary gland
C1526200|Guidance for biopsy:Find:Pt:Salivary gland:Doc:US
C1526200|Guidance for biopsy:Finding:Point in time:Salivary gland:Document:Ultrasound
C1526213|Carot a+VA-R XRA W contr IA
C1526213|Carotid artery+Vertebral artery - right Fluoroscopic angiogram W contrast IA
C1526213|Views^W contrast IA:Find:Pt:Carotid artery+Vertebral artery.right:Doc:XR.fluor.angio
C1526213|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Vertebral artery.right:Document:XR.fluor.angio
C1526223|Orbit vv-R XRA W contr IV
C1526223|Orbit veins - right Fluoroscopic angiogram W contrast IV
C1526223|Views^W contrast Intravenous:Finding:Point in time:Orbit veins.right:Document:XR.fluor.angio
C1526223|Views^W contrast IV:Find:Pt:Orbit veins.right:Doc:XR.fluor.angio
C1526304|Breast specimen - left Mammogram
C1526304|Brst specimen-L Mam
C1526304|Views:Find:Pt:Breast specimen.left:Doc:Mam
C1526304|Views:Finding:Point in time:Breast specimen.left:Document:Mam
C1526323|Kidney XR W contr retro
C1526323|Views^W contrast retrograde:Finding:Point in time:Kidney:Document:XR
C1526323|Kidney X-ray W contrast retrograde
C1526323|Views^W contrast retrograde:Find:Pt:Kidney:Doc:XR
C1524857|Forearm CT WO contr
C1524857|Forearm CT WO contrast
C1524857|Multisection^WO contrast:Find:Pt:Forearm:Doc:CT
C1524857|Multisection^WO contrast:Finding:Point in time:Forearm:Document:Computerized Tomography
C1524150|Should-L CT WO contr
C1524150|Shoulder - left CT WO contrast
C1524150|Multisection^WO contrast:Finding:Point in time:Shoulder.left:Document:Computerized Tomography
C1524150|Multisection^WO contrast:Find:Pt:Shoulder.left:Doc:CT
C1524548|LE.joint-L MRI W contr IV
C1524548|Lower extremity joint - left MRI W contrast IV
C1524548|Multisection^W contrast IV:Find:Pt:Lower extremity.joint.left:Doc:MRI
C1524548|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.joint.left:Document:MRI
C1524938|Humerus XR 1V
C1524938|Humerus X-ray Single view
C1524938|View 1:Finding:Point in time:Humerus:Document:XR
C1524938|View 1:Find:Pt:Humerus:Doc:XR
C0881863|Chest X-ray AP portable single view
C0881863|Chest XR AP V1 port
C0881863|View AP portable:Find:Pt:Chest:Doc:XR
C0881863|View AP portable:Finding:Point in time:Chest:Document:XR
C1524941|Femur XR Lat
C1524941|Femur X-ray lateral
C1524941|View lateral:Finding:Point in time:Femur:Document:XR
C1524941|View lateral:Find:Pt:Femur:Doc:XR
C1524286|CT Guidance for aspiration of cyst of Unspecified body region
C1524286|XXX CT Cyst Asp guid
C1524286|Guidance for aspiration of cyst:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1524286|Guidance for aspiration of cyst:Find:Pt:XXX:Doc:CT
C1524605|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Aorta.abdominal:Doc:CT
C1524605|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Aorta.abdominal:Document:Computerized Tomography
C1524605|Abdominal Aorta CT WO and W contrast IV
C1524605|Abd Aorta CT WO+W contr IV
C1524615|Lower extremity - bilateral MRI WO and W contrast IV
C1524615|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.bilateral:Doc:MRI
C1524615|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.bilateral:Document:MRI
C1524615|LE-Bl MRI WO+W contr IV
C1524621|Ankle-Bl XR 3V
C1524621|Ankle - bilateral X-ray 3 views
C1524621|Views 3:Find:Pt:Ankle.bilateral:Doc:XR
C1524621|Views 3:Finding:Point in time:Ankle.bilateral:Document:XR
C1524952|Knee XR Lat
C1524952|Knee X-ray lateral
C1524952|View lateral:Finding:Point in time:Knee:Document:XR
C1524952|View lateral:Find:Pt:Knee:Doc:XR
C1524962|Ft XR Obl 1V
C1524962|Foot X-ray oblique single view
C1524962|View oblique:Find:Pt:Foot:Doc:XR
C1524962|View oblique:Finding:Point in time:Foot:Document:XR
C1524969|Hand X-ray PA
C1524969|Hand XR PA V1
C1524969|View PA:Find:Pt:Hand:Doc:XR
C1524969|View PA:Finding:Point in time:Hand:Document:XR
C1524317|Kidney CT Drain guid
C1524317|CT Guidance for drainage of Kidney
C1524317|Guidance for drainage:Finding:Point in time:Kidney:Document:Computerized Tomography
C1524317|Guidance for drainage:Find:Pt:Kidney:Doc:CT
C1524319|CT Guidance for drainage of Lymph node
C1524319|LN CT Drain guid
C1524319|Guidance for drainage:Finding:Point in time:Lymph node:Document:Computerized Tomography
C1524319|Guidance for drainage:Find:Pt:Lymph node:Doc:CT
C1524328|CT Guidance for localization of Breast - right
C1524328|Brst-R CT Localization guid
C1524328|Guidance for localization:Find:Pt:Breast.right:Doc:CT
C1524328|Guidance for localization:Finding:Point in time:Breast.right:Document:Computerized Tomography
C1524330|Pelvis CT Nerve Block guid
C1524330|CT Guidance for nerve block of Pelvis
C1524330|Guidance for nerve block:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1524330|Guidance for nerve block:Find:Pt:Pelvis:Doc:CT
C1524332|Spine CT PC Vertebroplasty guid
C1524332|CT Guidance for percutaneous vertebroplasty of Spine
C1524332|Guidance for percutaneous vertebroplasty:Finding:Point in time:Spine:Document:Computerized Tomography
C1524332|Guidance for percutaneous vertebroplasty:Find:Pt:Spine:Doc:CT
C1524337|CT Guidance for placement of tube in Chest
C1524337|Chest CT Tube plac guid
C1524337|Guidance for placement of tube:Find:Pt:Chest:Doc:CT
C1524337|Guidance for placement of tube:Finding:Point in time:Chest:Document:Computerized Tomography
C1524632|Foot - bilateral X-ray 3 views
C1524632|Ft-Bl XR 3V
C1524632|Views 3:Finding:Point in time:Foot.bilateral:Document:XR
C1524632|Views 3:Find:Pt:Foot.bilateral:Doc:XR
C1524646|Chest X-ray 4 views
C1524646|Chest XR 4V
C1524646|Views 4:Find:Pt:Chest:Doc:XR
C1524646|Views 4:Finding:Point in time:Chest:Document:XR
C1524659|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.right:Doc:MRI
C1524659|Lower extremity - right MRI WO and W contrast IV
C1524659|LE-R MRI WO+W contr IV
C1524659|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.right:Document:MRI
C1524660|Multisection^WO & W contrast IV:Find:Pt:Upper extremity:Doc:CT
C1524660|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity:Document:Computerized Tomography
C1524660|UE CT WO+W contr IV
C1524660|Upper extremity CT WO and W contrast IV
C1524662|Upper extremity - right CT WO and W contrast IV
C1524662|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.right:Doc:CT
C1524662|UE-R CT WO+W contr IV
C1524662|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.right:Document:Computerized Tomography
C1524363|Esophagus CT
C1524363|Esoph CT
C1524363|Multisection:Finding:Point in time:Esophagus:Document:Computerized Tomography
C1524363|Multisection:Find:Pt:Esophagus:Doc:CT
C1524370|LE-L CT
C1524370|Lower extremity - left CT
C1524370|Multisection:Finding:Point in time:Lower extremity.left:Document:Computerized Tomography
C1524370|Multisection:Find:Pt:Lower extremity.left:Doc:CT
C1524730|Foot - left MRI WO and W contrast IV
C1524730|Multisection^WO & W contrast IV:Find:Pt:Foot.left:Doc:MRI
C1524730|Multisection^WO & W contrast Intravenous:Finding:Point in time:Foot.left:Document:MRI
C1524730|Ft-L MRI WO+W contr IV
C1524795|Multisection^WO & W contrast IV:Find:Pt:Lower leg.left:Doc:MRI
C1524795|Lower leg-L MRI WO+W contr IV
C1524795|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower leg.left:Document:MRI
C1524795|Lower leg - left MRI WO and W contrast IV
C1830192|Guidance for drainage^WO & W contrast IV:Find:Pt:XXX:Doc:CT
C1830192|Guidance for drainage^WO & W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1830192|CT Guidance for drainage of Unspecified body region-- WO and W contrast IV
C1830192|XXX CT Drain guid WO+W contr IV
C1830194|CT Guidance for drainage of Unspecified body region-- WO contrast
C1830194|XXX CT Drain guid WO contr
C1830194|Guidance for drainage^WO contrast:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1830194|Guidance for drainage^WO contrast:Find:Pt:XXX:Doc:CT
C1830221|Orbit+Face CT W contr IV
C1830221|Orbit and Face CT W contrast IV
C1830221|Multisection^W contrast IV:Find:Pt:Head>Orbit+Face:Doc:CT
C1830221|Multisection^W contrast Intravenous:Finding:Point in time:Head>Orbit+Face:Document:Computerized Tomography
C1830266|Celiac plexus CT Ablation guid
C1830266|CT Guidance for ablation of tissue of Celiac plexus
C1830266|Guidance for ablation of tissue:Finding:Point in time:Chest>Celiac plexus:Document:Computerized Tomography
C1830266|Guidance for ablation of tissue:Find:Pt:Chest>Celiac plexus:Doc:CT
C1715378|CT Guidance for fine needle aspiration of Prostate
C1715378|Prostate CT FNA Asp
C1715378|Guidance for aspiration.fine needle:Find:Pt:Prostate:Doc:CT
C1715378|Guidance for aspiration.fine needle:Finding:Point in time:Prostate:Document:Computerized Tomography
C1715398|Lower extremity vessels MRI angiogram WO and W contrast IV
C1715398|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity vessels:Document:MRI.angio
C1715398|Multisection^WO & W contrast IV:Find:Pt:Lower extremity vessels:Doc:MRI.angio
C1715398|LE ves MRI.Angio WO+W contr IV
C1715431|Multisection & 3D reconstruction:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1715431|Multisection & 3D reconstruction:Find:Pt:XXX:Doc:US
C1715431|Deprecated Unspecified body region US and 3D reconstruction
C1715431|Deprecated XXX US +3DR
C1717317|Ft XR GE 3V
C1717317|Foot X-ray GE 3 views
C1717317|Views GE 3:Finding:Point in time:Foot:Document:XR
C1717317|Views GE 3:Find:Pt:Foot:Doc:XR
C1715457|Hand X-ray GE 3 Portable views
C1715457|Hand XR GE 3V Port
C1715457|Views GE 3 portable:Finding:Point in time:Hand:Document:XR
C1715457|Views GE 3 portable:Find:Pt:Hand:Doc:XR
C1715466|C+T+L-spine XR port
C1715466|Spine Cervical and Thoracic and Lumbar X-ray portable
C1715466|Views portable:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:XR
C1715466|Views portable:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:XR
C1715474|PD Flr Endo guid W contr retro
C1715474|Fluoroscopy Guidance for endoscopy of Pancreatic duct-- W contrast retrograde
C1715474|Guidance for endoscopy^W contrast retrograde:Finding:Point in time:Pancreatic duct:Document:XR.fluor
C1715474|Guidance for endoscopy^W contrast retrograde:Find:Pt:Pancreatic duct:Doc:XR.fluor
C1715482|Fluoroscopy Guidance for procedure of Joint space
C1715482|Joint space Flr Procedure guid
C1715482|Guidance for procedure:Find:Pt:Joint space:Doc:XR.fluor
C1715482|Guidance for procedure:Finding:Point in time:Joint space:Document:XR.fluor
C1715487|Colon Fluoroscopy W barium contrast PR
C1715487|Colon Flr W Ba PR
C1715487|Views^W barium contrast PR:Find:Pt:Colon:Doc:XR.fluor
C1715487|Views^W barium contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C1715496|Views:Finding:Point in time:Trachea:Narrative:XR
C1715496|Trachea X-ray
C1715496|Trachea XR
C1715496|Views:Finding:Point in time:Trachea:Document:XR
C1715496|Views:Find:Pt:Trachea:Doc:XR
C1634501|Brst Flr Bx needle guid
C1634501|Fluoroscopy Guidance for needle biopsy of Breast
C1634501|Guidance for biopsy.needle:Finding:Point in time:Breast:Document:XR.fluor
C1634501|Guidance for biopsy.needle:Find:Pt:Breast:Doc:XR.fluor
C1714816|Joint XR Lat W Stress
C1714816|Joint X-ray lateral W manual stress
C1714816|Views lateral^W manual stress:Find:Pt:Joint:Doc:XR
C1714816|Views lateral^W manual stress:Finding:Point in time:Joint:Document:XR
C1714906|Axilla-R MRI W contr IV
C1714906|Axilla - right MRI W contrast IV
C1714906|Multisection^W contrast IV:Find:Pt:Axilla.right:Doc:MRI
C1714906|Multisection^W contrast Intravenous:Finding:Point in time:Axilla.right:Document:MRI
C1714922|Sinuses X-ray 1 or 2 views
C1714922|Sinuses XR 1V or 2V
C1714922|Views 1 or 2:Find:Pt:Sinuses:Doc:XR
C1714922|Views 1 or 2:Finding:Point in time:Sinuses:Document:XR
C1714941|Carotid artery - unilateral US
C1714941|Carot a-UL US
C1714941|Multisection:Finding:Point in time:Carotid artery.unilateral:Document:Ultrasound
C1714941|Multisection:Find:Pt:Carotid artery.unilateral:Doc:US
C1714950|Chest and Abdomen X-ray AP upright and AP chest
C1714950|Chest+Abd XR AP Upr+AP Chst
C1714950|Views AP upright & AP chest:Find:Pt:Chest+Abdomen:Doc:XR
C1714950|Views AP upright & AP chest:Finding:Point in time:Chest+Abdomen:Document:XR
C1717262|Guidance for deep biopsy:Find:Pt:Bone:Doc:US
C1717262|Bone US Guidance for deep biopsy
C1717262|Guidance for deep biopsy:Finding:Point in time:Bone:Document:Ultrasound
C1717262|US Guidance for deep biopsy of Bone
C1714954|Guidance for deep biopsy:Find:Pt:Bone:Doc:CT
C1714954|Bone CT Guidance for deep biopsy
C1714954|CT Guidance for deep biopsy of Bone
C1714954|Guidance for deep biopsy:Finding:Point in time:Bone:Document:Computerized Tomography
C1715107|Spine Cervicothoracic Junction X-ray
C1715107|CTJ XR
C1715107|Views:Find:Pt:Spine.cervicothoracic junction:Doc:XR
C1715107|Views:Finding:Point in time:Spine.cervicothoracic junction:Document:XR
C1630191|Skull X-ray stereo
C1630191|Skull XR Stereo
C1630191|View stereo:Finding:Point in time:Skull:Document:XR
C1630191|View stereo:Find:Pt:Skull:Doc:XR
C1634492|Pelvis+Hip-L XR 2V
C1634492|Pelvis and Hip - left X-ray 2 views
C1634492|Views 2:Finding:Point in time:Pelvis+Hip.left:Document:XR
C1634492|Views 2:Find:Pt:Pelvis+Hip.left:Doc:XR
C1632229|Scrotum+Test RI Flow W RNC IV
C1632229|Scrotum and Testicle Scan flow
C1632229|Views flow^W radionuclide Intravenous:Finding:Point in time:Scrotum+Testicle:Document:Radnuc
C1632229|Views flow^W radionuclide IV:Find:Pt:Scrotum+Testicle:Doc:Radnuc
C1624134|US Guidance for injection of Pleural space
C1624134|Pl space US Inj guid
C1624134|Guidance for injection:Finding:Point in time:Chest>Pleural space:Document:Ultrasound
C1624134|Guidance for injection:Find:Pt:Chest>Pleural space:Doc:US
C1624700|C-spine XR Ltd
C1624700|Views limited:Find:Pt:Spine.cervical:Doc:XR
C1624700|Views limited:Finding:Point in time:Spine.cervical:Document:XR
C1624700|Cervical spine X-ray limited
C1977322|Hrt SPECT Rest+W Tc99mMIBI IV
C1977322|Heart SPECT at rest and W Tc-99m Sestamibi IV
C1977322|Multisection^at rest & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1977322|Multisection^at rest & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1954309|Skull.base XR 1V
C1954309|Skull.base X-ray Single view
C1954309|View 1:Find:Pt:Skull.base:Doc:XR
C1954309|View 1:Finding:Point in time:Skull.base:Document:XR
C1953946|Skull.base MRI W contr IV
C1953946|Skull.base MRI W contrast IV
C1953946|Multisection^W contrast Intravenous:Finding:Point in time:Skull.base:Document:MRI
C1953946|Multisection^W contrast IV:Find:Pt:Skull.base:Doc:MRI
C1953956|Multisection^WO & W contrast IT:Find:Pt:Spine.cervical:Doc:MRI
C1953956|Multisection^WO & W contrast Intrathecal:Finding:Point in time:Spine.cervical:Document:MRI
C1953956|C-spine MRI WO+W contr IT
C1953956|Cervical spine MRI WO and W contrast IT
C1953971|Views:Finding:Point in time:Larynx:Narrative:XR.fluor
C1953971|Larynx Flr
C1953971|Larynx Fluoroscopy
C1953971|Views:Finding:Point in time:Larynx:Document:XR.fluor
C1953971|Views:Find:Pt:Larynx:Doc:XR.fluor
C2925713|Hrt MRI W Stress
C2925713|Heart MRI W stress
C2925713|Multisection^W stress:Finding:Point in time:Heart:Document:MRI
C2925713|Multisection^W stress:Find:Pt:Heart:Doc:MRI
C3533905|Multisection screening:Finding:Point in time:Breast.right:Document:Mam.FFD.tomosynthesis
C3533905|Brst-R FFDM-DBT Screening
C3533905|Breast - right FFD mammogram-tomosynthesis screening
C3533905|Multisection screening:Find:Pt:Breast.right:Doc:Mam.FFD.tomosynthesis
C3533793|Multisection^WO contrast:Find:Pt:Chest+Abdomen+Pelvis:Doc:CT
C3533793|Chest and Abdomen and Pelvis CT WO contrast
C3533793|Chest+Abd+Pelvis CT WO contr
C3533793|Multisection^WO contrast:Finding:Point in time:Chest+Abdomen+Pelvis:Document:Computerized Tomography
C3262929|Multisection^W contrast IS:Find:Pt:Knee.left:Doc:CT
C3262929|Knee - left CT W contrast IS
C3262929|Multisection^W contrast Intrasynovial:Finding:Point in time:Knee.left:Document:Computerized Tomography
C3262929|Knee-L CT W contr IS
C3262967|Knee - left X-ray AP and lateral and right oblique and left oblique
C3262967|Knee-L XR AP+Lat+R-Obl+L-Obl
C3262967|Views AP & lateral & R-oblique & L-oblique:Finding:Point in time:Knee.left:Document:XR
C3262967|Views AP & lateral & R-oblique & L-oblique:Find:Pt:Knee.left:Doc:XR
C3262978|Brst implant XR Screening
C3262978|Breast implant X-ray screening
C3262978|Views screening:Finding:Point in time:Breast implant:Document:XR
C3262978|Views screening:Find:Pt:Breast implant:Doc:XR
C3262471|Finger - left MRI W contrast IV
C3262471|Finger-L MRI W contr IV
C3262471|Multisection^W contrast IV:Find:Pt:Finger.left:Doc:MRI
C3262471|Multisection^W contrast Intravenous:Finding:Point in time:Finger.left:Document:MRI
C3262472|Finger - left MRI WO contrast
C3262472|Finger-L MRI WO contr
C3262472|Multisection^WO contrast:Find:Pt:Finger.left:Doc:MRI
C3262472|Multisection^WO contrast:Finding:Point in time:Finger.left:Document:MRI
C3263025|Pelvis MRI limited
C3263025|Pelvis MRI Ltd
C3263025|Multisection limited:Find:Pt:Pelvis:Doc:MRI
C3263025|Multisection limited:Finding:Point in time:Pelvis:Document:MRI
C3263072|Patella-R XR 1V
C3263072|Patella - right X-ray Single view
C3263072|View 1:Finding:Point in time:Patella.right:Document:XR
C3263072|View 1:Find:Pt:Patella.right:Doc:XR
C3263092|US Guidance for aspiration of Breast - left
C3263092|Brst-L US Asp guid
C3263092|Guidance for aspiration:Finding:Point in time:Breast.left:Document:Ultrasound
C3263092|Guidance for aspiration:Find:Pt:Breast.left:Doc:US
C3262885|Knee - bilateral X-ray 4 views standing
C3262885|Knee-Bl XR 4V stand
C3262885|Views 4^standing:Find:Pt:Knee.bilateral:Doc:XR
C3262885|Views 4^standing:Finding:Point in time:Knee.bilateral:Document:XR
C3262913|Shoulder - bilateral CT WO contrast
C3262913|Should-Bl CT WO contr
C3262913|Multisection^WO contrast:Find:Pt:Shoulder.bilateral:Doc:CT
C3262913|Multisection^WO contrast:Finding:Point in time:Shoulder.bilateral:Document:Computerized Tomography
C0942161|Radius+Ulna-R XR
C0942161|Radius - right and Ulna - right X-ray
C0942161|Views:Finding:Point in time:Radius.right+Ulna.right:Document:XR
C0942161|Views:Find:Pt:Radius.right+Ulna.right:Doc:XR
C0942177|Toes-L XR
C0942177|Toes - left X-ray
C0942177|Views:Find:Pt:Toes.left:Doc:XR
C0942177|Views:Finding:Point in time:Toes.left:Document:XR
C0942200|Thigh - bilateral MRI WO and W contrast IV
C0942200|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thigh.bilateral:Document:MRI
C0942200|Thigh-Bl MRI WO+W contr IV
C0942200|Multisection^WO & W contrast IV:Find:Pt:Thigh.bilateral:Doc:MRI
C0942211|Wrist-R MRI WO+W contr IV
C0942211|Multisection^WO & W contrast IV:Find:Pt:Wrist.right:Doc:MRI
C0942211|Wrist - right MRI WO and W contrast IV
C0942211|Multisection^WO & W contrast Intravenous:Finding:Point in time:Wrist.right:Document:MRI
C0942220|Carotid artery - bilateral US
C0942220|Carot a-Bl US
C0942220|Multisection:Finding:Point in time:Carotid artery.bilateral:Document:Ultrasound
C0942220|Multisection:Find:Pt:Carotid artery.bilateral:Doc:US
C0942228|Extremity - left CT
C0942228|Extr-L CT
C0942228|Multisection:Find:Pt:Extremity.left:Doc:CT
C0942228|Multisection:Finding:Point in time:Extremity.left:Document:Computerized Tomography
C0942262|Shoulder - left US
C0942262|Should-L US
C0942262|Multisection:Finding:Point in time:Shoulder.left:Document:Ultrasound
C0942262|Multisection:Find:Pt:Shoulder.left:Doc:US
C0942279|Knee-R XR Merchants
C0942279|Knee - right X-ray Merchants
C0942279|View Merchants:Finding:Point in time:Knee.right:Document:XR
C0942279|View Merchants:Find:Pt:Knee.right:Doc:XR
C0942307|CT Guidance for injection of Sacroiliac joint - left
C0942307|SIJ-L CT Inj guid
C0942307|Guidance for injection:Finding:Point in time:Sacroiliac joint.left:Document:Computerized Tomography
C0942307|Guidance for injection:Find:Pt:Sacroiliac joint.left:Doc:CT
C0942316|US Guidance for drainage of Kidney - left
C0942316|Kidney-L US Drain guid
C0942316|Guidance for drainage:Finding:Point in time:Kidney.left:Document:Ultrasound
C0942316|Guidance for drainage:Find:Pt:Kidney.left:Doc:US
C0942320|Mammogram Guidance for core needle percutaneous biopsy of Breast - bilateral
C0942320|Brst-Bl Mam PC Bx CN guid
C0942320|Guidance for percutaneous biopsy.core needle:Find:Pt:Breast.bilateral:Doc:Mam
C0942320|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast.bilateral:Document:Mam
C0945342|Wrist+Hand-L XR Bone Age
C0945342|Wrist - left and Hand - left X-ray bone age
C0945342|Views bone age:Find:Pt:Wrist.left+Hand.left:Doc:XR
C0945342|Views bone age:Finding:Point in time:Wrist.left+Hand.left:Document:XR
C0942347|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Brachiocephalic artery.bilateral:Narrative:XR.fluor.angio
C0942347|Angioplasty^W contrast IA:Find:Pt:Brachiocephalic artery.bilateral:Nar:XR.fluor.angio
C0942347|Deprecated Brachiocephalic artery - bilateral Fluoroscopic angiogram Angioplasty W contrast IA
C0942347|Deprecated BrachCeph a-Bl XRA Angpsty W
C0882049|CT Guidance for aspiration of Pancreas
C0882049|Pancreas CT Asp guid
C0882049|Guidance for aspiration:Find:Pt:Abdomen>Pancreas:Doc:CT
C0882049|Guidance for aspiration:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C0882062|Pelvis+Hip MRI
C0882062|Pelvis and Hip MRI
C0882062|Multisection:Find:Pt:Pelvis+Hip:Doc:MRI
C0882062|Multisection:Finding:Point in time:Pelvis+Hip:Document:MRI
C0882070|Popliteal a XRA PTA of ves W contr IA
C0882070|Popliteal artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C0882070|Percutaneous transluminal angioplasty of vessel^W contrast IA:Find:Pt:Popliteal artery:Doc:XR.fluor.angio
C0882070|Percutaneous transluminal angioplasty of vessel^W contrast Intra-arterial:Finding:Point in time:Popliteal artery:Document:XR.fluor.angio
C0882095|Sinus tract Fluoroscopy W contrast intra sinus tract
C0882095|Sinus tr Flr W contr intra ST
C0882095|Views^W contrast intra sinus tract:Find:Pt:Sinus tract:Doc:XR.fluor
C0882095|Views^W contrast intra sinus tract:Finding:Point in time:Sinus tract:Document:XR.fluor
C0882120|C-spine XR 3V
C0882120|Views 3:Finding:Point in time:Spine.cervical:Document:XR
C0882120|Views 3:Find:Pt:Spine.cervical:Doc:XR
C0882120|Cervical spine X-ray 3 views
C0882144|T+L-spine XR 2V
C0882144|Spine Thoracic and Lumbar X-ray 2 views
C0882144|Views 2:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C0882144|Views 2:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C0882149|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Spleen:Document:Computerized Tomography
C0882149|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Spleen:Doc:CT
C0882149|Spleen CT WO and W contrast IV
C0882149|Spleen CT WO+W contr IV
C0882150|Spleen US
C0882150|Multisection:Find:Pt:Spleen:Doc:US
C0882150|Multisection:Finding:Point in time:Spleen:Document:Ultrasound
C0882189|Wrist MRI
C0882189|Multisection:Finding:Point in time:Wrist:Narrative:MRI
C0882189|Multisection:Finding:Point in time:Wrist:Document:MRI
C0882189|Multisection:Find:Pt:Wrist:Doc:MRI
C0882226|Kidney arteries Fluoroscopic angiogram W contrast IA
C0882226|Kidney aa XRA W contr IA
C0882226|Views^W contrast Intra-arterial:Finding:Point in time:Kidney arteries:Document:XR.fluor.angio
C0882226|Views^W contrast IA:Find:Pt:Kidney arteries:Doc:XR.fluor.angio
C0942092|Salivary gland - right Fluoroscopy W contrast intra salivary duct
C0942092|Salivary gland-R Flr W contr intra SD
C0942092|Views^W contrast intra salivary duct:Finding:Point in time:Salivary gland.right:Document:XR.fluor
C0942092|Views^W contrast intra salivary duct:Find:Pt:Salivary gland.right:Doc:XR.fluor
C0942134|Femur - bilateral X-ray
C0942134|Femur-Bl XR
C0942134|Views:Find:Pt:Femur.bilateral:Doc:XR
C0942134|Views:Finding:Point in time:Femur.bilateral:Document:XR
C0881818|Brachiocephalic artery Fluoroscopic angiogram Angioplasty W contrast IA
C0881818|BrachCeph a XRA Angpsty W contr IA
C0881818|Angioplasty^W contrast IA:Find:Pt:Brachiocephalic artery:Doc:XR.fluor.angio
C0881818|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Brachiocephalic artery:Document:XR.fluor.angio
C0881834|Mammogram Guidance for aspiration of Breast
C0881834|Brst Mam Asp guid
C0881834|Guidance for aspiration:Finding:Point in time:Breast:Document:Mam
C0881834|Guidance for aspiration:Find:Pt:Breast:Doc:Mam
C0881838|Brst Mam Bx Str Guid
C0881838|Mammogram Guidance for stereotactic biopsy of Breast
C0881838|Guidance for stereotactic biopsy:Finding:Point in time:Breast:Document:Mam
C0881838|Guidance for stereotactic biopsy:Find:Pt:Breast:Doc:Mam
C0881845|Views:Find:Pt:Calcaneus:Doc:XR
C0881845|Deprecated Calcaneus X-ray
C0881845|Deprecated Heel XR
C0881845|Views:Finding:Point in time:Calcaneus:Document:XR
C0881856|Centl v XRA Cath plac guid W contr IV
C0881856|Fluoroscopic angiogram Guidance for placement of catheter in Central vein-- W contrast IV
C0881856|Guidance for placement of catheter^W contrast IV:Find:Pt:Central vein:Doc:XR.fluor.angio
C0881856|Guidance for placement of catheter^W contrast Intravenous:Finding:Point in time:Central vein:Document:XR.fluor.angio
C0881859|Multisection^W contrast Intravenous:Finding:Point in time:Chest:Narrative:COMPUTERIZED TOMOGRAPHY
C0881859|Chest CT W contr IV
C0881859|Chest CT W contrast IV
C0881859|Multisection^W contrast IV:Find:Pt:Chest:Doc:CT
C0881859|Multisection^W contrast Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C0881870|Chest XR AP+PA Upr
C0881870|Views AP & PA upright:Find:Pt:Chest:Doc:XR
C0881870|Views AP & PA upright:Finding:Point in time:Chest:Document:XR
C0881870|Chest X-ray AP and PA upright
C0881878|Chest XR AP R-Lat Debuc Port
C0881878|Chest X-ray AP right lateral-decubitus portable
C0881878|View AP R-lateral-decubitus portable:Finding:Point in time:Chest:Document:XR
C0881878|View AP R-lateral-decubitus portable:Find:Pt:Chest:Doc:XR
C0882528|Lower Extremity Joint MRI
C0882528|LE.joint MRI
C0882528|Multisection:Find:Pt:Lower extremity.joint:Doc:MRI
C0882528|Multisection:Finding:Point in time:Lower extremity.joint:Document:MRI
C0881914|Extr CT W contr IV
C0881914|Extremity CT W contrast IV
C0881914|Multisection^W contrast Intravenous:Finding:Point in time:Extremity:Document:Computerized Tomography
C0881914|Multisection^W contrast IV:Find:Pt:Extremity:Doc:CT
C0881933|GI RI W Tc99mRBC IV
C0881933|Gastrointestine Scan W Tc-99m tagged RBC IV
C0881933|Views^W Tc-99m tagged RBC Intravenous:Finding:Point in time:Gastrointestine:Document:Radnuc
C0881933|Views^W Tc-99m tagged RBC IV:Find:Pt:Gastrointestine:Doc:Radnuc
C0881936|Ileal conduit X-ray Loopogram
C0881936|Ileal conduit XR Loopogram
C0881936|Loopogram:Find:Pt:Ileal conduit:Doc:XR
C0881936|Loopogram:Finding:Point in time:Ileal conduit:Document:XR
C0881943|Multisection:Finding:Point in time:Head:Narrative:COMPUTERIZED TOMOGRAPHY
C0881943|Head CT
C0881943|Multisection:Find:Pt:Head:Doc:CT
C0881943|Multisection:Finding:Point in time:Head:Document:Computerized Tomography
C0882540|Liver CT W contr IV
C0882540|Liver CT W contrast IV
C0882540|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C0882540|Multisection^W contrast IV:Find:Pt:Abdomen>Liver:Doc:CT
C1114489|C-spine MRI WO contr
C1114489|Multisection^WO contrast:Finding:Point in time:Spine.cervical:Document:MRI
C1114489|Multisection^WO contrast:Find:Pt:Spine.cervical:Doc:MRI
C1114489|Cervical spine MRI WO contrast
C1114504|Forearm MRI WO+W contr IV
C1114504|Multisection^WO & W contrast Intravenous:Finding:Point in time:Forearm:Document:MRI
C1114504|Multisection^WO & W contrast IV:Find:Pt:Forearm:Doc:MRI
C1114504|Forearm MRI WO and W contrast IV
C1114561|Should XR 5V
C1114561|Shoulder X-ray 5 views
C1114561|Views 5:Find:Pt:Shoulder:Doc:XR
C1114561|Views 5:Finding:Point in time:Shoulder:Document:XR
C1114589|Ft XR 2V
C1114589|Foot X-ray 2 views
C1114589|Views 2:Finding:Point in time:Foot:Document:XR
C1114589|Views 2:Find:Pt:Foot:Doc:XR
C1114590|Ft XR W forced dorsiflex
C1114590|Foot X-ray W forced dorsiflexion
C1114590|Views^W forced dorsiflexion:Find:Pt:Foot:Doc:XR
C1114590|Views^W forced dorsiflexion:Finding:Point in time:Foot:Document:XR
C1114949|C+T+L-spine Flr W contr IT
C1114949|Spine Cervical and Thoracic and Lumbar Fluoroscopy W contrast IT
C1114949|Views^W contrast Intrathecal:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:XR.fluor
C1114949|Views^W contrast IT:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:XR.fluor
C1114949|VIEWS^W CONTRAST.XXX INTRATHECAL:FINDING:POINT IN TIME:SPINAL CORD.CERVICAL AND THORACIC AND LUMBAR:NARRATIVE:XR.FLUOR
C1114657|Carot ves+Neck ves MRI.Angio
C1114657|Carotid vessels and Neck Vessels MRI angiogram
C1114657|Multisection:Finding:Point in time:Carotid vessels+Neck vessels:Document:MRI.angio
C1114657|Multisection:Find:Pt:Carotid vessels+Neck vessels:Doc:MRI.angio
C2713072|Deprecated US.doppler
C2713072|Deprecated Abdominal vessels US.doppler Multisection
C2713072|Multisection:Find:Pt:Vessels.abdomen:Nar:US.doppler
C2713072|Multisection:Finding:Point in time:Vessels.abdomen:Narrative:Ultrasound.doppler
C1114440|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Liver:Doc:CT
C1114440|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1114440|Liver CT WO+W contr IV
C1114440|Liver CT WO and W contrast IV
C1114444|Multisection^WO & W contrast IV:Find:Pt:Pelvis:Doc:CT
C1114444|Pelvis CT WO and W contrast IV
C1114444|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1114444|Pelvis CT WO+W contr IV
C1114452|LE CT W contr IV
C1114452|Lower extremity CT W contrast IV
C1114452|Multisection^W contrast IV:Find:Pt:Lower extremity:Doc:CT
C1114452|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity:Document:Computerized Tomography
C1526829|Kidney-L Flr W contr RU
C1526829|Views^W contrast retrograde via urethra:Finding:Point in time:Kidney.left:Document:XR.fluor
C1526829|Kidney - left Fluoroscopy W contrast retrograde via urethra
C1526829|Views^W contrast retrograde via urethra:Find:Pt:Kidney.left:Doc:XR.fluor
C1543426|Chest XR Lat+PA W insp+exp
C1543426|Chest X-ray lateral and PA W inspiration and expiration
C1543426|Views lateral & PA^W inspiration & expiration:Find:Pt:Chest:Doc:XR
C1543426|Views lateral & PA^W inspiration & expiration:Finding:Point in time:Chest:Document:XR
C1543446|Chest Flr Tube plac guid
C1543446|Fluoroscopy Guidance for placement of tube in Chest
C1543446|Guidance for placement of tube:Finding:Point in time:Chest:Document:XR.fluor
C1543446|Guidance for placement of tube:Find:Pt:Chest:Doc:XR.fluor
C1543450|Scapula XR Lat+Outlet
C1543450|Scapula X-ray lateral and outlet
C1543450|Views lateral & outlet:Finding:Point in time:Scapula:Document:XR
C1543450|Views lateral & outlet:Find:Pt:Scapula:Doc:XR
C2713301|Knee-R XR 2V+Obl
C2713301|Knee - right X-ray 2 views and oblique
C2713301|Views 2 & oblique:Find:Pt:Knee.right:Doc:XR
C2713301|Views 2 & oblique:Finding:Point in time:Knee.right:Document:XR
C1543469|Knee-R XR +Sunrise
C1543469|Knee - right X-ray and Sunrise
C1543469|Views & Sunrise:Find:Pt:Knee.right:Doc:XR
C1543469|Views & Sunrise:Finding:Point in time:Knee.right:Document:XR
C1543780|Hrt RI PF Rest+W RNC IV
C1543780|Heart Scan perfusion at rest and W radionuclide IV
C1543780|Views perfusion^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543780|Views perfusion^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543782|Views perfusion^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1543782|Hrt RI PF W Stress+W RNC IV
C1543782|Heart Scan perfusion W stress and W radionuclide IV
C1543782|Views perfusion^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543782|Views perfusion^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543788|Hrt SPECT PF W Stress+W Tc99mMIBI IV
C1543788|Heart SPECT perfusion W stress and W Tc-99m Sestamibi IV
C1543788|Multisection perfusion^W stress & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543788|Multisection perfusion^W stress & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1542975|Spleen Scan
C1542975|Spleen RI W RNC IV
C1542975|Views^W radionuclide Intravenous:Finding:Point in time:Spleen:Narrative:Radnuc
C1542975|Views^W radionuclide Intravenous:Finding:Point in time:Spleen:Document:Radnuc
C1542975|Views^W radionuclide IV:Find:Pt:Spleen:Doc:Radnuc
C1543811|Stomach Scan for gastric emptying W radionuclide PO
C1543811|Stom RI GE W RNC PO
C1543811|Views for gastric emptying^W radionuclide Oral:Finding:Point in time:Stomach:Document:Radnuc
C1543811|Views for gastric emptying^W radionuclide PO:Find:Pt:Stomach:Doc:Radnuc
C1543855|Bone SPECT Ltd W RNC IV
C1543855|Bone SPECT limited
C1543855|Multisection limited^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1543855|Multisection limited^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1543858|Bone SPECT whole body
C1543858|Bone SPECT WB W RNC IV
C1543858|Multisection whole body^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1543858|Multisection whole body^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1542906|SPECT W In-111 Satmb IV
C1542906|SPECT W In-111 Satumomab IV
C1542906|Multisection^W In-111 Satumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1542906|Multisection^W In-111 Satumomab IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543898|Liver+Spleen SPECT W RNC IV
C1543898|Liver and Spleen SPECT
C1543898|Multisection^W radionuclide Intravenous:Finding:Point in time:Liver+Spleen:Document:Radnuc.SPECT
C1543898|Multisection^W radionuclide IV:Find:Pt:Liver+Spleen:Doc:Radnuc.SPECT
C1543923|Bone RI 3 Phase Mul Areas W RNC IV
C1543923|Bone Scan 3 views phase multiple areas
C1543923|Views 3 phase multiple areas^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543923|Views 3 phase multiple areas ^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543580|Femoral vessels - right US.doppler
C1543580|Fem ves-R DOP
C1543580|Multisection:Find:Pt:Femoral vessels.right:Doc:US.doppler
C1543580|Multisection:Finding:Point in time:Femoral vessels.right:Document:Ultrasound.doppler
C1526350|Bone density:Mass Aeric:Point in time:Hip:Quantitative:XR.DXA
C1526350|Hip DXA Bone density
C1526350|Bone density:MAric:Pt:Hip:Qn:XR.DXA
C1526350|Hip DXA BDM
C1543168|Hip Fluoroscopy during surgery
C1543168|Hip Flr in Surg
C1543168|View^during surgery:Find:Pt:Hip:Doc:XR.fluor
C1543168|View^during surgery:Finding:Point in time:Hip:Document:XR.fluor
C1543586|Lymphatics pelvic Fluoroscopy W contrast intra lymphatic
C1543586|Lymph Pelvic Flr W contr IL
C1543586|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.pelvic:Document:XR.fluor
C1543586|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.pelvic:Doc:XR.fluor
C1543260|XXX US VA guid
C1543260|US Guidance for vascular access of Unspecified body region
C1543260|Guidance for vascular access:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1543260|Guidance for vascular access:Find:Pt:XXX:Doc:US
C1524258|Should-R XR AP+Ax+Y
C1524258|Shoulder - right X-ray AP and axillary and Y
C1524258|Views AP & axillary & Y:Find:Pt:Shoulder.right:Doc:XR
C1524258|Views AP & axillary & Y:Finding:Point in time:Shoulder.right:Document:XR
C1526810|Brst-L Mam Mag+Spot
C1526810|Breast - left Mammogram magnification and spot
C1526810|Views magnification & spot:Find:Pt:Breast.left:Doc:Mam
C1526810|Views magnification & spot:Finding:Point in time:Breast.left:Document:Mam
C1524438|Posterior fossa MRI
C1524438|Post fossa MRI
C1524438|Multisection:Finding:Point in time:Posterior fossa:Document:MRI
C1524438|Multisection:Find:Pt:Posterior fossa:Doc:MRI
C1527073|Spleen MRI
C1527073|Multisection:Finding:Point in time:Spleen:Narrative:MRI
C1527073|Multisection:Find:Pt:Spleen:Doc:MRI
C1527073|Multisection:Finding:Point in time:Spleen:Document:MRI
C1524819|Appendix CT WO contrast
C1524819|Appendix CT WO contr
C1524819|Multisection^WO contrast:Find:Pt:Abdomen+Pelvis>Appendix:Doc:CT
C1524819|Multisection^WO contrast:Finding:Point in time:Abdomen+Pelvis>Appendix:Document:Computerized Tomography
C1524828|Elbow CT WO contrast
C1524828|Elbow CT WO contr
C1524828|Multisection^WO contrast:Find:Pt:Elbow:Doc:CT
C1524828|Multisection^WO contrast:Finding:Point in time:Elbow:Document:Computerized Tomography
C1525175|Knee vessels MRI angiogram
C1525175|Knee ves MRI.Angio
C1525175|Multisection:Finding:Point in time:Knee vessels:Document:MRI.angio
C1525175|Multisection:Find:Pt:Knee vessels:Doc:MRI.angio
C1525188|Multisection^W contrast IS:Find:Pt:Joint:Doc:MRI
C1525188|Multisection^W contrast Intrasynovial:Finding:Point in time:Joint:Document:MRI
C1525188|Joint MRI W contr IS
C1525188|Joint MRI W contrast IS
C1525288|Orbit+Face MRI WO contr
C1525288|Orbit and Face MRI WO contrast
C1525288|Multisection^WO contrast:Find:Pt:Orbit+Face:Doc:MRI
C1525288|Multisection^WO contrast:Finding:Point in time:Orbit+Face:Document:MRI
C1525258|Mastoid X-ray 5 views
C1525258|Mastoid XR 5V
C1525258|Views 5:Find:Pt:Mastoid:Doc:XR
C1525258|Views 5:Finding:Point in time:Mastoid:Document:XR
C1525337|Breast - left Mammogram magnification
C1525337|Brst-L Mam Mag
C1525337|View magnification:Find:Pt:Breast.left:Doc:Mam
C1525337|View magnification:Finding:Point in time:Breast.left:Document:Mam
C1524688|Knee - bilateral X-ray Rosenberg standing
C1524688|Knee-Bl XR Rosenberg stand
C1524688|View Rosenberg^standing:Find:Pt:Knee.bilateral:Doc:XR
C1524688|View Rosenberg^standing:Finding:Point in time:Knee.bilateral:Document:XR
C1525473|Fetal X-ray
C1525473|Fet XR
C1525473|Views:Finding:Point in time:^Fetus:Document:XR
C1525473|Views:Find:Pt:^Fetus:Doc:XR
C1525477|Ribs-L XR 2V
C1525477|Ribs - left X-ray 2 views
C1525477|Views 2:Find:Pt:Ribs.left:Doc:XR
C1525477|Views 2:Finding:Point in time:Ribs.left:Document:XR
C1525496|Abd XR AP(sup+Lat Decub)
C1525496|Abdomen X-ray AP (supine and lateral-decubitus)
C1525496|Views AP (supine & lateral-decubitus):Finding:Point in time:Abdomen:Document:XR
C1525496|Views AP (supine & lateral-decubitus):Find:Pt:Abdomen:Doc:XR
C1525519|Abd XR AP+Obl
C1525519|Abdomen X-ray AP and oblique
C1525519|Views AP & oblique:Finding:Point in time:Abdomen:Document:XR
C1525519|Views AP & oblique:Find:Pt:Abdomen:Doc:XR
C1525528|Should-L XR Ax+Y
C1525528|Shoulder - left X-ray axillary and Y
C1525528|Views axillary & Y:Find:Pt:Shoulder.left:Doc:XR
C1525528|Views axillary & Y:Finding:Point in time:Shoulder.left:Document:XR
C1525563|Face XR Lat+Caldwell+Waters
C1525563|Facial bones X-ray lateral and Caldwell and Waters
C1525563|Views lateral & Caldwell & Waters:Finding:Point in time:Facial bones:Document:XR
C1525563|Views lateral & Caldwell & Waters:Find:Pt:Facial bones:Doc:XR
C1525613|Brain Stem+Nerves.cranial MRI
C1525613|Brain Stem and Nerves.cranial MRI
C1525613|Multisection:Find:Pt:Brain stem+Nerves.cranial:Doc:MRI
C1525613|Multisection:Finding:Point in time:Brain stem+Nerves.cranial:Document:MRI
C1525749|Wrist-Bl CT
C1525749|Wrist - bilateral CT
C1525749|Multisection:Find:Pt:Wrist.bilateral:Doc:CT
C1525749|Multisection:Finding:Point in time:Wrist.bilateral:Document:Computerized Tomography
C1525871|GB XR W contr+Fatty Meal PO
C1525871|Gallbladder X-ray W contrast and fatty meal PO
C1525871|Views^W contrast & fatty meal PO:Find:Pt:Gallbladder:Doc:XR
C1525871|Views^W contrast & fatty meal Oral:Finding:Point in time:Gallbladder:Document:XR
C1525885|Ac arch+Carot a.com-L XRA W contr IA
C1525885|Aortic arch and Carotid artery.common - left Fluoroscopic angiogram W contrast IA
C1525885|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery.common.left:Document:XR.fluor.angio
C1525885|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery.common.left:Doc:XR.fluor.angio
C1525819|LS-spine junc XR Lat Spot stand
C1525819|Spine Lumbosacral Junction X-ray lateral spot standing
C1525819|View lateral spot^standing:Finding:Point in time:Spine.lumbosacral junction:Document:XR
C1525819|View lateral spot^standing:Find:Pt:Spine.lumbosacral junction:Doc:XR
C1525828|Toe 5th-L XR
C1525828|Toe fifth - left X-ray
C1525828|Views:Finding:Point in time:Toe.fifth.left:Document:XR
C1525828|Views:Find:Pt:Toe.fifth.left:Doc:XR
C1525964|Sacroiliac Joint Fluoroscopy W contrast IS
C1525964|SIJ Flr W contr IS
C1525964|Views^W contrast Intrasynovial:Finding:Point in time:Sacroiliac joint:Document:XR.fluor
C1525964|Views^W contrast IS:Find:Pt:Sacroiliac joint:Doc:XR.fluor
C1526134|Should XR AP 1V
C1526134|Shoulder X-ray AP single view
C1526134|View AP:Finding:Point in time:Shoulder:Document:XR
C1526134|View AP:Find:Pt:Shoulder:Doc:XR
C1526037|Hip - right X-ray 2 views
C1526037|Hip-R XR 2V
C1526037|Views 2:Finding:Point in time:Hip.right:Document:XR
C1526037|Views 2:Find:Pt:Hip.right:Doc:XR
C1526073|Knee-R XR Obl
C1526073|Knee - right X-ray oblique
C1526073|Views oblique:Find:Pt:Knee.right:Doc:XR
C1526073|Views oblique:Finding:Point in time:Knee.right:Document:XR
C1526076|Knee-R XRTomo
C1526076|Knee - right X-ray tomograph
C1526076|Multisection:Find:Pt:Knee.right:Doc:XR.tomo
C1526076|Multisection:Finding:Point in time:Knee.right:Document:XR.tomo
C1526092|Scapula-R XR 2V
C1526092|Scapula - right X-ray 2 views
C1526092|Views 2:Finding:Point in time:Scapula.right:Document:XR
C1526092|Views 2:Find:Pt:Scapula.right:Doc:XR
C1526144|Sinuses XR Caldwell+Waters
C1526144|Sinuses X-ray Caldwell and Waters
C1526144|Views Caldwell & Waters:Find:Pt:Sinuses:Doc:XR
C1526144|Views Caldwell & Waters:Finding:Point in time:Sinuses:Document:XR
C1526148|Sinuses X-ray 5 views
C1526148|Sinuses XR 5V
C1526148|Views 5:Find:Pt:Sinuses:Doc:XR
C1526148|Views 5:Finding:Point in time:Sinuses:Document:XR
C1526153|Sinuses XR SMV
C1526153|Sinuses X-ray submentovertex
C1526153|View submentovertex:Find:Pt:Sinuses:Doc:XR
C1526153|View submentovertex:Finding:Point in time:Sinuses:Document:XR
C1526185|T-spine XR 2V
C1526185|Views 2:Finding:Point in time:Spine.thoracic:Document:XR
C1526185|Views 2:Find:Pt:Spine.thoracic:Doc:XR
C1526185|Thoracic spine X-ray 2 views
C1526188|T-spine XR AP+Lat+Obl
C1526188|Views AP & lateral & oblique:Finding:Point in time:Spine.thoracic:Document:XR
C1526188|Views AP & lateral & oblique:Find:Pt:Spine.thoracic:Doc:XR
C1526188|Thoracic spine X-ray AP and lateral and oblique
C1524703|Wrist X-ray 2 views
C1524703|Wrist XR 2V
C1524703|Views 2:Find:Pt:Wrist:Doc:XR
C1524703|Views 2:Finding:Point in time:Wrist:Document:XR
C1524712|Kidney US Ltd
C1524712|Kidney US limited
C1524712|Multisection limited:Find:Pt:Kidney:Doc:US
C1524712|Multisection limited:Finding:Point in time:Kidney:Document:Ultrasound
C1526275|Lower extremity artery US.doppler limited
C1526275|LE a DOP Ltd
C1526275|Multisection limited:Finding:Point in time:Lower extremity artery:Document:Ultrasound.doppler
C1526275|Multisection limited:Find:Pt:Lower extremity artery:Doc:US.doppler
C1508087|Breast - bilateral Mammogram W air
C1508087|Brst-Bl Mam W Air
C1508087|Views^W air:Finding:Point in time:Breast.bilateral:Document:Mam
C1508087|Views^W air:Find:Pt:Breast.bilateral:Doc:Mam
C1526321|C-spine+L-spine Flr W contr IT
C1526321|Spine Cervical and Spine Lumbar Fluoroscopy W contrast IT
C1526321|Views^W contrast IT:Find:Pt:Spine.cervical+Spine.lumbar:Doc:XR.fluor
C1526321|Views^W contrast Intrathecal:Finding:Point in time:Spine.cervical+Spine.lumbar:Document:XR.fluor
C1524504|Elbow-L MRI W contr IV
C1524504|Elbow - left MRI W contrast IV
C1524504|Multisection^W contrast Intravenous:Finding:Point in time:Elbow.left:Document:MRI
C1524504|Multisection^W contrast IV:Find:Pt:Elbow.left:Doc:MRI
C1524904|Prostate MRI WO contr
C1524904|Prostate MRI WO contrast
C1524904|Multisection^WO contrast:Finding:Point in time:Prostate:Document:MRI
C1524904|Multisection^WO contrast:Find:Pt:Prostate:Doc:MRI
C1524145|Sacrum MRI WO contrast
C1524145|Sacrum MRI WO contr
C1524145|Multisection^WO contrast:Finding:Point in time:Sacrum:Document:MRI
C1524145|Multisection^WO contrast:Find:Pt:Sacrum:Doc:MRI
C1524919|Portal vein MRI angiogram WO contrast
C1524919|Portal v MRI.Angio WO contr
C1524919|Multisection^WO contrast:Finding:Point in time:Portal vein:Document:MRI.angio
C1524919|Multisection^WO contrast:Find:Pt:Portal vein:Doc:MRI.angio
C1524575|TO-R MRI W contr IV
C1524575|Thoracic outlet - right MRI W contrast IV
C1524575|Multisection^W contrast Intravenous:Finding:Point in time:Thoracic outlet.right:Document:MRI
C1524575|Multisection^W contrast IV:Find:Pt:Thoracic outlet.right:Doc:MRI
C1524576|Post fossa CT W contr IV
C1524576|Posterior fossa CT W contrast IV
C1524576|Multisection^W contrast IV:Find:Pt:Posterior fossa:Doc:CT
C1524576|Multisection^W contrast Intravenous:Finding:Point in time:Posterior fossa:Document:Computerized Tomography
C1524942|Finger.5th XR Lat
C1524942|Finger fifth X-ray lateral
C1524942|View lateral:Find:Pt:Finger.fifth:Doc:XR
C1524942|View lateral:Finding:Point in time:Finger.fifth:Document:XR
C1524288|Chest Flr Bronch guid
C1524288|Fluoroscopy Guidance for bronchoscopy of Chest
C1524288|Guidance for bronchoscopy:Find:Pt:Chest:Doc:XR.fluor
C1524288|Guidance for bronchoscopy:Finding:Point in time:Chest:Document:XR.fluor
C1524298|Fluoroscopy Guidance for biopsy of Kidney
C1524298|Kidney Flr Bx guid
C1524298|Guidance for biopsy:Finding:Point in time:Kidney:Document:XR.fluor
C1524298|Guidance for biopsy:Find:Pt:Kidney:Doc:XR.fluor
C1524589|Sinuses CT W contr IV
C1524589|Sinuses CT W contrast IV
C1524589|Multisection^W contrast IV:Find:Pt:Head>Sinuses:Doc:CT
C1524589|Multisection^W contrast Intravenous:Finding:Point in time:Head>Sinuses:Document:Computerized Tomography
C1524618|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.right:Document:Computerized Tomography
C1524618|Lower extremity - right CT WO and W contrast IV
C1524618|LE-R CT WO+W contr IV
C1524618|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.right:Doc:CT
C1524980|Humerus-L XR
C1524980|Humerus - left X-ray
C1524980|Views:Find:Pt:Humerus.left:Doc:XR
C1524980|Views:Finding:Point in time:Humerus.left:Document:XR
C1524636|Knee - bilateral X-ray 3 views
C1524636|Knee-Bl XR 3V
C1524636|Views 3:Find:Pt:Knee.bilateral:Doc:XR
C1524636|Views 3:Finding:Point in time:Knee.bilateral:Document:XR
C1525003|Finger XR 2V
C1525003|Finger X-ray 2 views
C1525003|Views 2:Finding:Point in time:Finger:Document:XR
C1525003|Views 2:Find:Pt:Finger:Doc:XR
C1525031|LE XR AP+Lat
C1525031|Lower extremity X-ray AP and lateral
C1525031|Views AP & lateral:Find:Pt:Lower extremity:Doc:XR
C1525031|Views AP & lateral:Finding:Point in time:Lower extremity:Document:XR
C1524403|Hip XRTomo
C1524403|Hip X-ray tomograph
C1524403|Multisection:Find:Pt:Hip:Doc:XR.tomo
C1524403|Multisection:Finding:Point in time:Hip:Document:XR.tomo
C1524409|Hip - left MRI
C1524409|Hip-L MRI
C1524409|Multisection:Find:Pt:Hip.left:Doc:MRI
C1524409|Multisection:Finding:Point in time:Hip.left:Document:MRI
C1524786|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C1524786|Multisection^WO & W contrast IV:Find:Pt:Spine.cervical:Doc:CT
C1524786|C-spine CT WO+W contr IV
C1524786|Cervical spine CT WO and W contrast IV
C1830187|Mammogram Guidance for needle biopsy of Breast
C1830187|Brst Mam Bx needle guid
C1830187|Guidance for biopsy.needle:Find:Pt:Breast:Doc:Mam
C1830187|Guidance for biopsy.needle:Finding:Point in time:Breast:Document:Mam
C1830237|Brst-L Mam 1V
C1830237|Breast - left Mammogram Single view
C1830237|View 1:Finding:Point in time:Breast.left:Document:Mam
C1830237|View 1:Find:Pt:Breast.left:Doc:Mam
C1830267|SPECT Guidance for biopsy of Bone
C1830267|Bone SPECT Bx guid W RNC IV
C1830267|Guidance for biopsy^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1830267|Guidance for biopsy^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1830268|CT Guidance for needle biopsy of Adrenal gland
C1830268|Adrenal CT Bx needle guid
C1830268|Guidance for biopsy.needle:Find:Pt:Abdomen>Adrenal gland:Doc:CT
C1830268|Guidance for biopsy.needle:Finding:Point in time:Abdomen>Adrenal gland:Document:Computerized Tomography
C1715397|Heart MRI limited cine for function
C1715397|Hrt MRI limited cine for function
C1715397|Multisection limited cine for function:Finding:Point in time:Heart:Document:MRI
C1715397|Multisection limited cine for function:Find:Pt:Heart:Doc:MRI
C1715424|US Guidance for ablation of tissue of Kidney
C1715424|Kidney US Ablation guid
C1715424|Guidance for ablation of tissue:Find:Pt:Kidney:Doc:US
C1715424|Guidance for ablation of tissue:Finding:Point in time:Kidney:Document:Ultrasound
C1715489|Multisection:Find:Pt:Bone:Doc:CT
C1715489|Bone CT
C1715489|Multisection:Finding:Point in time:Bone:Document:Computerized Tomography
C1648949|Ribs-L+Chest XR +PA Chst
C1648949|Ribs - left and Chest X-ray and PA chest
C1648949|Views & PA chest:Finding:Point in time:Ribs.left+Chest:Document:XR
C1648949|Views & PA chest:Find:Pt:Ribs.left+Chest:Doc:XR
C1631816|L-spine XR AP W R+L-bending
C1631816|Views AP^W R-bending & W L-bending:Find:Pt:Spine.lumbar:Doc:XR
C1631816|Views AP^W R-bending & W L-bending:Finding:Point in time:Spine.lumbar:Document:XR
C1631816|Lumbar spine X-ray AP W right bending and W left bending
C1714801|Ribs - bilateral and Chest X-ray lateral and PA chest
C1714801|Views lateral & PA chest:Find:Pt:Ribs.bilateral+Chest:Doc:XR
C1714801|Views lateral & PA chest:Finding:Point in time:Ribs.bilateral+Chest:Document:XR
C1714801|Ribs-Bl+Chest XR Lat+PA Chst
C1714819|Thumb - right X-ray GE 3 views
C1714819|Thumb-R XR GE 3V
C1714819|Views GE 3:Finding:Point in time:Thumb.right:Document:XR
C1714819|Views GE 3:Find:Pt:Thumb.right:Doc:XR
C1714930|Deprecated Eye US Bleeding local guid
C1714930|Guidance for localization of bleeding site:Find:Pt:Eye:Nar:US
C1714930|Deprecated US Guidance for localization of bleeding site of Eye
C1714930|Guidance for localization of bleeding site:Finding:Point in time:Eye:Narrative:Ultrasound
C1714937|Pelvis XR GE 3V
C1714937|Pelvis X-ray GE 3 views
C1714937|Views GE 3:Find:Pt:Pelvis:Doc:XR
C1714937|Views GE 3:Finding:Point in time:Pelvis:Document:XR
C1714783|Pulmonary system CT
C1714783|Pulm CT
C1714783|Multisection:Find:Pt:Pulmonary system:Doc:CT
C1714783|Multisection:Finding:Point in time:Pulmonary system:Document:Computerized Tomography
C1715035|Thyroid Scan spot
C1715035|Thyroid RI Spot W RNC IV
C1715035|View spot^W radionuclide IV:Find:Pt:Thyroid:Doc:Radnuc
C1715035|View spot^W radionuclide Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1636060|Ft.Sesamoids XR AP+Lat
C1636060|Foot sesamoid bones X-ray AP and lateral
C1636060|Views AP & lateral:Finding:Point in time:Foot.sesamoid bones:Document:XR
C1636060|Views AP & lateral:Find:Pt:Foot.sesamoid bones:Doc:XR
C1634998|Brst-Bl Mam p wire plac
C1634998|Breast - bilateral Mammogram Post Wire Placement
C1634998|Views^post wire placement:Finding:Point in time:Breast.bilateral:Document:Mam
C1634998|Views^post wire placement:Find:Pt:Breast.bilateral:Doc:Mam
C1635010|Knee - right X-ray 2 views and (views standing)
C1635010|Knee-R XR 2V+(views Stand)
C1635010|Views 2 & (views^standing):Finding:Point in time:Knee.right:Document:XR
C1635010|Views 2 & (views^standing):Find:Pt:Knee.right:Doc:XR
C1624665|Ribs-R+Chest XR +PA Chst
C1624665|Ribs - right and Chest X-ray and PA chest
C1624665|Views & PA chest:Finding:Point in time:Ribs.right+Chest:Document:XR
C1624665|Views & PA chest:Find:Pt:Ribs.right+Chest:Doc:XR
C1638468|LE ves graft-R DOP
C1638468|Lower extremity vessel graft - right US.doppler
C1638468|Multisection:Find:Pt:Lower extremity vessel graft.right:Doc:US.doppler
C1638468|Multisection:Finding:Point in time:Lower extremity vessel graft.right:Document:Ultrasound.doppler
C1640450|Iliac graft US.doppler limited
C1640450|Iliac Graft DOP Ltd
C1640450|Multisection limited:Find:Pt:Iliac graft:Doc:US.doppler
C1640450|Multisection limited:Finding:Point in time:Iliac graft:Document:Ultrasound.doppler
C1631784|Thyroid RI +Uptake W I-123 IV
C1631784|Thyroid Scan and uptake W I-123 IV
C1631784|Views & uptake^W I-123 IV:Find:Pt:Thyroid:Doc:Radnuc
C1631784|Views & uptake^W I-123 Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1630177|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space:Document:Computerized Tomography
C1630177|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space:Doc:CT
C1630177|CT Guidance for drainage of abscess of Pleural space
C1630177|Pl space CT Abscess drain guid
C3484380|Uterus MRI
C3484380|Multisection:Finding:Point in time:Uterus:Narrative:MRI
C3484380|Multisection:Find:Pt:Uterus:Doc:MRI
C3484380|Multisection:Finding:Point in time:Uterus:Document:MRI
C1633448|Clavicle MRI WO contrast
C1633448|Clavicle MRI WO contr
C1633448|Multisection^WO contrast:Finding:Point in time:Clavicle:Document:MRI
C1633448|Multisection^WO contrast:Find:Pt:Clavicle:Doc:MRI
C1632338|Head+Neck ves MRI.Angio
C1632338|Head vessels and Neck vessels MRI angiogram
C1632338|Multisection:Finding:Point in time:Head vessels+Neck vessels:Document:MRI.angio
C1632338|Multisection:Find:Pt:Head vessels+Neck vessels:Doc:MRI.angio
C1978439|Brst RI W Tl-201 IV
C1978439|Breast Scan W Tl-201 IV
C1978439|Views^W Tl-201 Intravenous:Finding:Point in time:Breast:Document:Radnuc
C1978439|Views^W Tl-201 IV:Find:Pt:Breast:Doc:Radnuc
C1953042|T-spine XR Obl
C1953042|Views oblique:Finding:Point in time:Spine.thoracic:Document:XR
C1953042|Views oblique:Find:Pt:Spine.thoracic:Doc:XR
C1953042|Thoracic spine X-ray oblique
C1953941|Fluoroscopy Guidance for injection of Salivary gland - bilateral
C1953941|Salivary gland-Bl Flr Inj guid
C1953941|Guidance for injection:Find:Pt:Salivary gland.bilateral:Doc:XR.fluor
C1953941|Guidance for injection:Finding:Point in time:Salivary gland.bilateral:Document:XR.fluor
C1952713|Brst implant-Bl Mam Screening
C1952713|Breast implant - bilateral Mammogram screening
C1952713|Views screening:Find:Pt:Breast implant.bilateral:Doc:Mam
C1952713|Views screening:Finding:Point in time:Breast implant.bilateral:Document:Mam
C2925711|Brain Functional MRI
C2925711|Brain fMRI
C2925711|Multisection:Finding:Point in time:Brain:Document:MRI.function
C2925711|Multisection:Find:Pt:Brain:Doc:MRI.function
C3533560|Guidance for facet joint denervation:Find:Pt:Spine.lumbar:Doc:XR.fluor
C3533560|L-spine Flr FJ DN guid
C3533560|Guidance for facet joint denervation:Finding:Point in time:Spine.lumbar:Document:XR.fluor
C3533560|Fluoroscopy Guidance for facet joint denervation of Lumbar spine
C3533804|Multisection^WO & W contrast IV:Find:Pt:Toes.left:Doc:MRI
C3533804|Multisection^WO & W contrast Intravenous:Finding:Point in time:Toes.left:Document:MRI
C3533804|Toes-L MRI WO+W contr IV
C3533804|Toes - left MRI WO and W contrast IV
C3262957|Iliac artery Fluoroscopic angiogram Atherectomy W contrast
C3262957|Iliac a XRA Atherect W contr
C3262957|Atherectomy^W contrast:Finding:Point in time:Iliac artery:Document:XR.fluor.angio
C3262957|Atherectomy^W contrast:Find:Pt:Iliac artery:Doc:XR.fluor.angio
C3266952|Hip-L XR +Danelius Miller
C3266952|Hip - left X-ray and Danelius Miller
C3266952|Views & Danelius Miller:Finding:Point in time:Hip.left:Document:XR
C3266952|Views & Danelius Miller:Find:Pt:Hip.left:Doc:XR
C3263039|Fluoroscopy Guidance for needle biopsy of Muscle
C3263039|Muscle Flr Bx needle guid
C3263039|Guidance for biopsy.needle:Find:Pt:Muscle:Doc:XR.fluor
C3263039|Guidance for biopsy.needle:Finding:Point in time:Muscle:Document:XR.fluor
C3261710|T-spine XR stand
C3261710|Views^standing:Finding:Point in time:Spine.thoracic:Document:XR
C3261710|Views^standing:Find:Pt:Spine.thoracic:Doc:XR
C3261710|Thoracic spine X-ray standing
C3263095|Renal vessels US
C3263095|Renal ves US
C3263095|Multisection:Find:Pt:Renal vessels:Doc:US
C3263095|Multisection:Finding:Point in time:Renal vessels:Document:Ultrasound
C3263207|US Guidance for cordocentesis
C3263207|Cordocentesis guid US
C3263207|Guidance for cordocentesis:Finding:Point in time:Umbilical cord^Fetus:Document:Ultrasound
C3263207|Guidance for cordocentesis:Find:Pt:Umbilical cord^fetus:Doc:US
C3263209|LE vv-L US
C3263209|Lower extremity veins - left US
C3263209|Multisection:Finding:Point in time:Lower extremity veins.left:Document:Ultrasound
C3263209|Multisection:Find:Pt:Lower extremity veins.left:Doc:US
C3263210|L-spine US
C3263210|Multisection:Finding:Point in time:Spine.lumbar:Document:Ultrasound
C3263210|Multisection:Find:Pt:Spine.lumbar:Doc:US
C3263210|Lumbar spine US
C3262884|Knee-Bl XR 2V+Tunnel
C3262884|Knee - bilateral X-ray 2 views and tunnel
C3262884|Views 2 & tunnel:Find:Pt:Knee.bilateral:Doc:XR
C3262884|Views 2 & tunnel:Finding:Point in time:Knee.bilateral:Document:XR
C3262903|C-spine XR 5V W FE
C3262903|Views 5^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C3262903|Views 5^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C3262903|Cervical spine X-ray 5 views W flexion and W extension
C0942150|Acromioclavicular joint - right X-ray
C0942150|AC joint-R XR
C0942150|Views:Find:Pt:Acromioclavicular joint.right:Doc:XR
C0942150|Views:Finding:Point in time:Acromioclavicular joint.right:Document:XR
C0942155|Optic foramen - left X-ray
C0942155|Optic foramen-L XR
C0942155|Views:Find:Pt:Optic foramen.left:Doc:XR
C0942155|Views:Finding:Point in time:Optic foramen.left:Document:XR
C0942169|Shoulder - right X-ray
C0942169|Should-R XR
C0942169|Views:Find:Pt:Shoulder.right:Doc:XR
C0942169|Views:Finding:Point in time:Shoulder.right:Document:XR
C0942179|Wrist-Bl XR
C0942179|Wrist - bilateral X-ray
C0942179|Views:Find:Pt:Wrist.bilateral:Doc:XR
C0942179|Views:Finding:Point in time:Wrist.bilateral:Document:XR
C0947255|TO ves-L MRI.Angio W contr IV
C0947255|Thoracic outlet vessels - left MRI angiogram W contrast IV
C0947255|Multisection^W contrast Intravenous:Finding:Point in time:Thoracic outlet vessels.left:Document:MRI.angio
C0947255|Multisection^W contrast IV:Find:Pt:Thoracic outlet vessels.left:Doc:MRI.angio
C0942196|Multisection^WO & W contrast IV:Find:Pt:Thoracic outlet.right:Doc:MRI
C0942196|TO-R MRI WO+W contr IV
C0942196|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thoracic outlet.right:Document:MRI
C0942196|Thoracic outlet - right MRI WO and W contrast IV
C0942205|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee.right:Document:MRI
C0942205|Knee-R MRI WO+W contr IV
C0942205|Multisection^WO & W contrast IV:Find:Pt:Knee.right:Doc:MRI
C0942205|Knee - right MRI WO and W contrast IV
C0942241|Ft-R MRI
C0942241|Foot - right MRI
C0942241|Multisection:Find:Pt:Foot.right:Doc:MRI
C0942241|Multisection:Finding:Point in time:Foot.right:Document:MRI
C0942252|Knee-L MRI
C0942252|Knee - left MRI
C0942252|Multisection:Find:Pt:Knee.left:Doc:MRI
C0942252|Multisection:Finding:Point in time:Knee.left:Document:MRI
C0942365|Ankle - left X-ray 2 views
C0942365|Ankle-L XR 2V
C0942365|Views 2:Find:Pt:Ankle.left:Doc:XR
C0942365|Views 2:Finding:Point in time:Ankle.left:Document:XR
C0942370|Humerus-L XR 2V
C0942370|Humerus - left X-ray 2 views
C0942370|Views 2:Find:Pt:Humerus.left:Doc:XR
C0942370|Views 2:Finding:Point in time:Humerus.left:Document:XR
C0942376|Hip - bilateral X-ray Single view
C0942376|Hip-Bl XR 1V
C0942376|View 1:Find:Pt:Hip.bilateral:Doc:XR
C0942376|View 1:Finding:Point in time:Hip.bilateral:Document:XR
C0882128|Bone density:MAric:Pt:Spine.lumbar:Qn:XR.DXA
C0882128|Bone density:Mass Aeric:Point in time:Spine.lumbar:Quantitative:XR.DXA
C0882128|L-spine DXA BDM
C0882128|Lumbar spine DXA Bone density
C0882147|Spine CT W contr IV
C0882147|Spine CT W contrast IV
C0882147|Multisection^W contrast Intravenous:Finding:Point in time:Spine:Document:Computerized Tomography
C0882147|Multisection^W contrast IV:Find:Pt:Spine:Doc:CT
C0882161|Scrotum+Test RI W Tc99mP IV
C0882161|Scrotum and Testicle Scan W Tc-99m pertechnetate IV
C0882161|Views^W Tc-99m pertechnetate Intravenous:Finding:Point in time:Scrotum+Testicle:Document:Radnuc
C0882161|Views^W Tc-99m pertechnetate IV:Find:Pt:Scrotum+Testicle:Doc:Radnuc
C0882187|Views^W radionuclide Intravenous:Finding:Point in time:Bone:Narrative:Radnuc
C0882187|Bone RI W RNC IV
C0882187|Bone Scan
C0882187|Views^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C0882187|Views^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C0882192|Wrist US
C0882192|Multisection:Find:Pt:Wrist:Doc:US
C0882192|Multisection:Finding:Point in time:Wrist:Document:Ultrasound
C0882562|Multisection sagittal & coronal:Find:Pt:XXX:Doc:CT
C0882562|Multisection sagittal & coronal:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0882562|Deprecated XXX CT Sagittal+Coronal
C0882562|Deprecated Unspecified body region CT sagittal and coronal
C0942145|Acetabulum - bilateral X-ray
C0942145|Acetabulum-Bl XR
C0942145|Views:Finding:Point in time:Acetabulum.bilateral:Document:XR
C0942145|Views:Find:Pt:Acetabulum.bilateral:Doc:XR
C0881787|Appendix US
C0881787|Multisection:Find:Pt:Appendix:Doc:US
C0881787|Multisection:Finding:Point in time:Appendix:Document:Ultrasound
C0881790|AVF XRA W contr IA
C0881790|AV fistula Fluoroscopic angiogram W contrast IA
C0881790|Views^W contrast Intra-arterial:Finding:Point in time:AV fistula:Document:XR.fluor.angio
C0881790|Views^W contrast IA:Find:Pt:AV fistula:Doc:XR.fluor.angio
C0881816|Bones SPECT W RNC IV
C0881816|Bones SPECT
C0881816|Multisection^W radionuclide IV:Find:Pt:Bones:Doc:Radnuc.SPECT
C0881816|Multisection^W radionuclide Intravenous:Finding:Point in time:Bones:Document:Radnuc.SPECT
C0881827|Multisection:Finding:Point in time:Brain:Narrative:MRI
C0881827|Brain MRI
C0881827|Multisection:Finding:Point in time:Brain:Document:MRI
C0881827|Multisection:Find:Pt:Brain:Doc:MRI
C0881843|Brst Mam Ltd
C0881843|Breast Mammogram limited
C0881843|Views limited:Finding:Point in time:Breast:Document:Mam
C0881843|Views limited:Find:Pt:Breast:Doc:Mam
C0881846|Cent CV a XRA Cath plac guid in art
C0881846|Fluoroscopic angiogram Guidance for placement of catheter in artery in Central cardiovascular artery
C0881846|Guidance for placement of catheter in artery:Find:Pt:Cardiovascular.central artery:Doc:XR.fluor.angio
C0881846|Guidance for placement of catheter in artery:Finding:Point in time:Cardiovascular.central artery:Document:XR.fluor.angio
C0881875|Chest X-ray PA upright
C0881875|Chest XR 1V PA Upr
C0881875|View PA upright:Find:Pt:Chest:Doc:XR
C0881875|View PA upright:Finding:Point in time:Chest:Document:XR
C0881886|Pleural space Fluoroscopy W contrast intra pleural space
C0881886|Pl space Flr W contr intra PS
C0881886|Views^W contrast intra pleural space:Finding:Point in time:Chest>Pleural space:Document:XR.fluor
C0881886|Views^W contrast intra pleural space:Find:Pt:Chest>Pleural space:Doc:XR.fluor
C0881905|Esoph Flr Dilation guid
C0881905|Fluoroscopy Guidance for dilation of Esophagus
C0881905|Guidance for dilation:Finding:Point in time:Esophagus:Document:XR.fluor
C0881905|Guidance for dilation:Find:Pt:Esophagus:Doc:XR.fluor
C0881912|Upper extremity MRI
C0881912|UE MRI
C0881912|Multisection:Find:Pt:Upper extremity:Doc:MRI
C0881912|Multisection:Finding:Point in time:Upper extremity:Document:MRI
C0881913|Upper extremity X-ray
C0881913|UE XR
C0881913|Views:Find:Pt:Upper extremity:Doc:XR
C0881913|Views:Finding:Point in time:Upper extremity:Document:XR
C0882163|Multisection:Finding:Point in time:Thigh:Narrative:MRI
C0882163|Thigh MRI
C0882163|Multisection:Find:Pt:Thigh:Doc:MRI
C0882163|Multisection:Finding:Point in time:Thigh:Document:MRI
C0881930|Forearm MRI
C0881930|Multisection:Find:Pt:Forearm:Doc:MRI
C0881930|Multisection:Finding:Point in time:Forearm:Document:MRI
C0881985|deprecated KD-Bl+CS XRTomo 1V
C0881985|View 1:Find:Pt:Kidney.bilateral+Collecting system:Nar:XR.tomo
C0881985|deprecated Kidney - bilateral & Collecting system X-ray tomograph Single view
C0881985|View 1:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:XR.tomo
C1114487|MRI Guidance for radiation treatment of Unspecified body region-- WO contrast
C1114487|XXX MRI RT guid WO contr
C1114487|Guidance for radiation treatment^WO contrast:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1114487|Guidance for radiation treatment^WO contrast:Find:Pt:XXX:Doc:MRI
C1114490|Abd MRI WO contr
C1114490|Abdomen MRI WO contrast
C1114490|Multisection^WO contrast:Finding:Point in time:Abdomen:Document:MRI
C1114490|Multisection^WO contrast:Find:Pt:Abdomen:Doc:MRI
C1114506|Multisection^WO & W contrast IV:Find:Pt:Hand:Doc:MRI
C1114506|Hand MRI WO+W contr IV
C1114506|Hand MRI WO and W contrast IV
C1114506|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hand:Document:MRI
C1114547|View AP lateral-decubitus:Finding:Point in time:Chest:Narrative:XR
C1114547|Chest XR AP Lat Decub
C1114547|Chest X-ray AP lateral-decubitus
C1114547|View AP lateral-decubitus:Find:Pt:Chest:Doc:XR
C1114547|View AP lateral-decubitus:Finding:Point in time:Chest:Document:XR
C1114619|FT Flr Cath guid transcervical
C1114619|Fluoroscopy Guidance for catheterization of Fallopian tubes-- transcervical
C1114619|Guidance for catheterization^transcervical:Find:Pt:Fallopian tubes:Doc:XR.fluor
C1114619|Guidance for catheterization^transcervical:Finding:Point in time:Fallopian tubes:Document:XR.fluor
C1114421|Pituitary and Sella turcica CT WO contrast
C1114421|Multisection^WO contrast:Find:Pt:Head>Pituitary+Sella turcica:Doc:CT
C1114421|Multisection^WO contrast:Finding:Point in time:Head>Pituitary+Sella turcica:Document:Computerized Tomography
C1114421|Head Pit+Slla turc CT WO contr
C1114460|Fluoroscopy Guidance for biopsy of Lung
C1114460|Lung Flr Bx guid
C1114460|Guidance for biopsy:Finding:Point in time:Lung:Document:XR.fluor
C1114460|Guidance for biopsy:Find:Pt:Lung:Doc:XR.fluor
C1114468|SVC XRA W contr IV
C1114468|Superior vena cava Fluoroscopic angiogram W contrast IV
C1114468|Views^W contrast Intravenous:Finding:Point in time:Vena cava.superior:Document:XR.fluor.angio
C1114468|Views^W contrast IV:Find:Pt:Vena cava.superior:Doc:XR.fluor.angio
C1543436|Ribs upper ant+post-L XR
C1543436|Ribs upper anterior and posterior - left X-ray
C1543436|Views:Finding:Point in time:Ribs.upper.anterior+posterior.left:Document:XR
C1543436|Views:Find:Pt:Ribs.upper.anterior+posterior.left:Doc:XR
C1543453|Ankle-R XR AP+Lat+Obl W Stress
C1543453|Ankle - right X-ray AP and lateral and oblique W manual stress
C1543453|Views AP & lateral & oblique^W manual stress:Find:Pt:Ankle.right:Doc:XR
C1543453|Views AP & lateral & oblique^W manual stress:Finding:Point in time:Ankle.right:Document:XR
C1744693|Deprecated Views perfusion^at rest & W stress & W 99m Tc Sestamibi IV:Find:Pt:Heart:Nar:Radnuc
C1744693|Deprecated Heart Scintigraphy perfusion at rest & W stress & W Tc-99m Sestamibi IV
C1744693|Views perfusion^at rest & W stress & W 99m Tc Sestamibi IV:Find:Pt:Heart:Nar:Radnuc
C1744693|Deprecated Hrt RI PF
C1744693|Views perfusion^at rest & W stress & W 99m Tc Sestamibi Intravenous:Finding:Point in time:Heart:Narrative:Radnuc
C1543459|Knee-R XR 2V+Sunrise
C1543459|Knee - right X-ray 2 views and Sunrise
C1543459|Views 2 & Sunrise:Find:Pt:Knee.right:Doc:XR
C1543459|Views 2 & Sunrise:Finding:Point in time:Knee.right:Document:XR
C1543798|Views^W Tc-99m Mertiatide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1543798|Views^W Tc-99m Mertiatide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1543798|Kidney - bilateral Scan W Tc-99m Mertiatide IV
C1543798|Kdny-Bl RI W Tc99mMAG3 IV
C1542977|Scrotum+Test RI W Tc99mDTPA IV
C1542977|Scrotum and Testicle Scan W Tc-99m DTPA IV
C1542977|Views^W Tc-99m DTPA IV:Find:Pt:Scrotum+Testicle:Doc:Radnuc
C1542977|Views^W Tc-99m DTPA Intravenous:Finding:Point in time:Scrotum+Testicle:Document:Radnuc
C1542926|Heart Scan flow
C1542926|Hrt RI Flow W RNC IV
C1542926|Views flow^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542926|Views flow^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543905|Bone RI 3 Phase W RNC IV
C1543905|Bone Scan 3 views phase
C1543905|Views 3 phase^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543905|Views 3 phase^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543943|Hrt RI Gated Rest+W RNC IV
C1543943|Heart Scan gated at rest and W radionuclide IV
C1543943|Views gated^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543943|Views gated^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543946|Hrt RI Gated Rest+stress+W RNC IV
C1543946|Heart Scan gated at rest and W stress and W radionuclide IV
C1543946|Views gated^at rest & W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543946|Views gated^at rest & W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543957|Lung RI V+EQ+WO W RNC IH
C1543957|Lung Scan ventilation and equilibrium and washout W radionuclide IH
C1543957|Views ventilation & equilibrium & washout^W radionuclide Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1543957|Views ventilation & equilibrium & washout^W radionuclide IH:Find:Pt:Lung:Doc:Radnuc
C1543503|Carotid artery - left US.doppler
C1543503|Carot a-L DOP
C1543503|Multisection:Finding:Point in time:Carotid artery.left:Document:Ultrasound.doppler
C1543503|Multisection:Find:Pt:Carotid artery.left:Doc:US.doppler
C1543198|Should XR AP+Transthoracic
C1543198|Shoulder X-ray AP and transthoracic
C1543198|Views AP & transthoracic:Finding:Point in time:Shoulder:Document:XR
C1543198|Views AP & transthoracic:Find:Pt:Shoulder:Doc:XR
C1543588|Hip-R XR +Danelius Miller
C1543588|Hip - right X-ray and Danelius Miller
C1543588|Views & Danelius Miller:Finding:Point in time:Hip.right:Document:XR
C1543588|Views & Danelius Miller:Find:Pt:Hip.right:Doc:XR
C1525928|Hand-R XR Brewerton
C1525928|Hand - right X-ray Brewerton
C1525928|View Brewerton:Finding:Point in time:Hand.right:Document:XR
C1525928|View Brewerton:Find:Pt:Hand.right:Doc:XR
C1543735|SPECT W Ga-67 IV
C1543735|Multisection^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc.SPECT
C1543735|Multisection^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc.SPECT
C1526802|Ft-L XR 2V
C1526802|Foot - left X-ray 2 views
C1526802|Views 2:Finding:Point in time:Foot.left:Document:XR
C1526802|Views 2:Find:Pt:Foot.left:Doc:XR
C1524436|Multisection:Finding:Point in time:Thoracic outlet:Narrative:COMPUTERIZED TOMOGRAPHY
C1524436|Thoracic outlet CT
C1524436|TO CT
C1524436|Multisection:Finding:Point in time:Thoracic outlet:Document:Computerized Tomography
C1524436|Multisection:Find:Pt:Thoracic outlet:Doc:CT
C1524848|Thigh - left MRI WO contrast
C1524848|Thigh-L MRI WO contr
C1524848|Multisection^WO contrast:Find:Pt:Thigh.left:Doc:MRI
C1524848|Multisection^WO contrast:Finding:Point in time:Thigh.left:Document:MRI
C1527065|Ovary MRI
C1527065|Multisection:Finding:Point in time:Ovary:Narrative:MRI
C1527065|Multisection:Finding:Point in time:Ovary:Document:MRI
C1527065|Multisection:Find:Pt:Ovary:Doc:MRI
C1525110|LE vv-L MRI.Angio
C1525110|Lower extremity veins - left MRI angiogram
C1525110|Multisection:Finding:Point in time:Lower extremity veins.left:Document:MRI.angio
C1525110|Multisection:Find:Pt:Lower extremity veins.left:Doc:MRI.angio
C1525177|Knee vessels - right MRI angiogram
C1525177|Knee ves-R MRI.Angio
C1525177|Multisection:Find:Pt:Knee vessels.right:Doc:MRI.angio
C1525177|Multisection:Finding:Point in time:Knee vessels.right:Document:MRI.angio
C1525183|Should ves-R MRI.Angio
C1525183|Shoulder vessels - right MRI angiogram
C1525183|Multisection:Find:Pt:Shoulder vessels.right:Doc:MRI.angio
C1525183|Multisection:Finding:Point in time:Shoulder vessels.right:Document:MRI.angio
C1525187|Joint CT W contrast IS
C1525187|Multisection^W contrast Intrasynovial:Finding:Point in time:Joint:Document:Computerized Tomography
C1525187|Joint CT W contr IS
C1525187|Multisection^W contrast IS:Find:Pt:Joint:Doc:CT
C1524453|Pelvis CT Ltd W contr IV
C1524453|Pelvis CT limited W contrast IV
C1524453|Multisection limited^W contrast Intravenous:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1524453|Multisection limited^W contrast IV:Find:Pt:Pelvis:Doc:CT
C1525309|View Harris:Finding:Point in time:Calcaneus.left:Document:XR
C1525309|Deprecated Calcaneus - left X-ray Harris
C1525309|Deprecated Heel-L XR Harris
C1525309|View Harris:Find:Pt:Calcaneus.left:Doc:XR
C1525193|UE joint-Bl MRI W contr IV
C1525193|Upper extremity joint - bilateral MRI W contrast IV
C1525193|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.joint.bilateral:Document:MRI
C1525193|Multisection^W contrast IV:Find:Pt:Upper extremity.joint.bilateral:Doc:MRI
C1525200|LE.R-veins CT W contr IV
C1525200|Lower extremity - right Veins CT W contrast IV
C1525200|Multisection^W contrast IV:Find:Pt:Lower extremity.right>Veins:Doc:CT
C1525200|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.right>Veins:Document:Computerized Tomography
C1525481|Wrist-Bl XR 4V
C1525481|Wrist - bilateral X-ray 4 views
C1525481|Views 4:Finding:Point in time:Wrist.bilateral:Document:XR
C1525481|Views 4:Find:Pt:Wrist.bilateral:Doc:XR
C1525486|Hip X-ray AP portable
C1525486|Hip XR AP ports
C1525486|Views AP portable:Find:Pt:Hip:Doc:XR
C1525486|Views AP portable:Finding:Point in time:Hip:Document:XR
C1525491|Should-Bl XR AP+Ax
C1525491|Shoulder - bilateral X-ray AP and axillary
C1525491|Views AP & axillary:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525491|Views AP & axillary:Find:Pt:Shoulder.bilateral:Doc:XR
C1524253|L-spine XR AP+Lat+Spot
C1524253|Views AP & lateral & spot:Find:Pt:Spine.lumbar:Doc:XR
C1524253|Views AP & lateral & spot:Finding:Point in time:Spine.lumbar:Document:XR
C1524253|Lumbar spine X-ray AP and lateral and spot
C1525511|Knee XR AP+Lat+Sunrise+Tunnel
C1525511|Knee X-ray AP and lateral and Sunrise and tunnel
C1525511|Views AP & lateral & Sunrise & tunnel:Find:Pt:Knee:Doc:XR
C1525511|Views AP & lateral & Sunrise & tunnel:Finding:Point in time:Knee:Document:XR
C1525552|Mastoid XR Stenver+Arcelin
C1525552|Mastoid X-ray Stenver and Arcelin
C1525552|Views Stenver & Arcelin:Find:Pt:Mastoid:Doc:XR
C1525552|Views Stenver & Arcelin:Finding:Point in time:Mastoid:Document:XR
C1525630|Great vessel MRI
C1525630|Great ves MRI
C1525630|Multisection:Find:Pt:Great vessel:Doc:MRI
C1525630|Multisection:Finding:Point in time:Great vessel:Document:MRI
C1525660|Brain+IAC MRI WO contr
C1525660|Brain and Internal auditory canal MRI WO contrast
C1525660|Multisection^WO contrast:Find:Pt:Brain+Internal auditory canal:Doc:MRI
C1525660|Multisection^WO contrast:Finding:Point in time:Brain+Internal auditory canal:Document:MRI
C1525700|Bones XR Bone Age
C1525700|Bones X-ray bone age
C1525700|Views bone age:Finding:Point in time:Bones:Document:XR
C1525700|Views bone age:Find:Pt:Bones:Doc:XR
C1525717|Carot a+VA XRA W contr IA
C1525717|Carotid artery and Vertebral artery Fluoroscopic angiogram W contrast IA
C1525717|Views^W contrast IA:Find:Pt:Carotid artery+Vertebral artery:Doc:XR.fluor.angio
C1525717|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Vertebral artery:Document:XR.fluor.angio
C1525752|Wrist-R CT
C1525752|Wrist - right CT
C1525752|Multisection:Finding:Point in time:Wrist.right:Document:Computerized Tomography
C1525752|Multisection:Find:Pt:Wrist.right:Doc:CT
C1525890|Nasal bones XRTomo
C1525890|Nasal bones X-ray tomograph
C1525890|Multisection:Finding:Point in time:Nasal bones:Document:XR.tomo
C1525890|Multisection:Find:Pt:Nasal bones:Doc:XR.tomo
C1525805|C-spine ves MRI.Angio W contr IV
C1525805|Cervical Spine vessels MRI angiogram W contrast IV
C1525805|Multisection^W contrast IV:Find:Pt:Spine.cervical vessels:Doc:MRI.angio
C1525805|Multisection^W contrast Intravenous:Finding:Point in time:Spine.cervical vessels:Document:MRI.angio
C1525823|Finger.4th-L XR
C1525823|Finger fourth - left X-ray
C1525823|Views:Find:Pt:Finger.fourth.left:Doc:XR
C1525823|Views:Finding:Point in time:Finger.fourth.left:Document:XR
C1525837|Mastoid-Bl XR Law+Mayer+Stenver+Towne
C1525837|Mastoid - bilateral X-ray law and Mayer and Stenver and Towne
C1525837|Views law & Mayer & Stenver & Towne:Find:Pt:Mastoid.bilateral:Doc:XR
C1525837|Views law & Mayer & Stenver & Towne:Finding:Point in time:Mastoid.bilateral:Document:XR
C1525984|Ankle-R XR AP+Lat+Obl
C1525984|Ankle - right X-ray AP and lateral and oblique
C1525984|Views AP & lateral & oblique:Find:Pt:Ankle.right:Doc:XR
C1525984|Views AP & lateral & oblique:Finding:Point in time:Ankle.right:Document:XR
C1525991|Ankle - right X-ray 2 views standing
C1525991|Ankle-R XR 2V stand
C1525991|Views 2^standing:Find:Pt:Ankle.right:Doc:XR
C1525991|Views 2^standing:Finding:Point in time:Ankle.right:Document:XR
C1526023|Radius+Ulna-R XR 2V
C1526023|Radius - right and Ulna - right X-ray 2 views
C1526023|Views 2:Finding:Point in time:Radius.right+Ulna.right:Document:XR
C1526023|Views 2:Find:Pt:Radius.right+Ulna.right:Doc:XR
C1525909|Should XR AP+Lat+Ax
C1525909|Shoulder X-ray AP and lateral and axillary
C1525909|Views AP & lateral & axillary:Find:Pt:Shoulder:Doc:XR
C1525909|Views AP & lateral & axillary:Finding:Point in time:Shoulder:Document:XR
C1526036|Views^standing:Find:Pt:Calcaneus.right:Doc:XR
C1526036|Deprecated Heel-R XR stand
C1526036|Deprecated Calcaneus - right X-ray standing
C1526036|Views^standing:Finding:Point in time:Calcaneus.right:Document:XR
C1526055|Iliac artery - right Fluoroscopic angiogram W contrast IA
C1526055|Iliac a-R XRA W contr IA
C1526055|Views^W contrast IA:Find:Pt:Iliac artery.right:Doc:XR.fluor.angio
C1526055|Views^W contrast Intra-arterial:Finding:Point in time:Iliac artery.right:Document:XR.fluor.angio
C1526075|Knee-R XR Sunrise+Tunnel
C1526075|Knee - right X-ray Sunrise and tunnel
C1526075|Views Sunrise & tunnel:Finding:Point in time:Knee.right:Document:XR
C1526075|Views Sunrise & tunnel:Find:Pt:Knee.right:Doc:XR
C1526101|Should-R XR 6V
C1526101|Shoulder - right X-ray 6 views
C1526101|Views 6:Find:Pt:Shoulder.right:Doc:XR
C1526101|Views 6:Finding:Point in time:Shoulder.right:Document:XR
C1526158|Sinuses X-ray tomograph
C1526158|Sinuses XRTomo
C1526158|Multisection:Finding:Point in time:Sinuses:Document:XR.tomo
C1526158|Multisection:Find:Pt:Sinuses:Doc:XR.tomo
C1526203|Zygomatic arch X-ray 3 views
C1526203|Zygomatic arch XR 3V
C1526203|Views 3:Find:Pt:Zygomatic arch:Doc:XR
C1526203|Views 3:Finding:Point in time:Zygomatic arch:Document:XR
C1526214|Carot a+Cerebral a-R XRA W contr IA
C1526214|Carotid artery and Cerebral artery - right Fluoroscopic angiogram W contrast IA
C1526214|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery+Cerebral artery.right:Document:XR.fluor.angio
C1526214|Views^W contrast IA:Find:Pt:Carotid artery+Cerebral artery.right:Doc:XR.fluor.angio
C1526235|Splenic v XRA W contr IV
C1526235|Splenic vein Fluoroscopic angiogram W contrast IV
C1526235|Views^W contrast IV:Find:Pt:Splenic vein:Doc:XR.fluor.angio
C1526235|Views^W contrast Intravenous:Finding:Point in time:Splenic vein:Document:XR.fluor.angio
C1526246|Lumbar Spine vessels MRI angiogram WO contrast
C1526246|L-spine ves MRI.Angio WO contr
C1526246|Multisection^WO contrast:Find:Pt:Spine.lumbar vessels:Doc:MRI.angio
C1526246|Multisection^WO contrast:Finding:Point in time:Spine.lumbar vessels:Document:MRI.angio
C1526293|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast implant.right:Document:MRI
C1526293|Brst implant-R MRI WO+W contr IV
C1526293|Breast implant - right MRI WO and W contrast IV
C1526293|Multisection^WO & W contrast IV:Find:Pt:Breast implant.right:Doc:MRI
C1526294|Breast implant - left MRI WO contrast
C1526294|Brst implant-L MRI WO contr
C1526294|Multisection^WO contrast:Finding:Point in time:Breast implant.left:Document:MRI
C1526294|Multisection^WO contrast:Find:Pt:Breast implant.left:Doc:MRI
C1526349|Wrist XR 6V
C1526349|Wrist X-ray 6 views
C1526349|Views 6:Finding:Point in time:Wrist:Document:XR
C1526349|Views 6:Find:Pt:Wrist:Doc:XR
C1524499|IAC MRI W contr IV
C1524499|Internal auditory canal MRI W contrast IV
C1524499|Multisection^W contrast Intravenous:Finding:Point in time:Internal auditory canal:Document:MRI
C1524499|Multisection^W contrast IV:Find:Pt:Internal auditory canal:Doc:MRI
C1524927|Ankle XR 1V
C1524927|Ankle X-ray Single view
C1524927|View 1:Find:Pt:Ankle:Doc:XR
C1524927|View 1:Finding:Point in time:Ankle:Document:XR
C1524551|SIJ CT W contr IV
C1524551|Sacroiliac Joint CT W contrast IV
C1524551|Multisection^W contrast Intravenous:Finding:Point in time:Sacroiliac joint:Document:Computerized Tomography
C1524551|Multisection^W contrast IV:Find:Pt:Sacroiliac joint:Doc:CT
C1524574|TO-L MRI W contr IV
C1524574|Thoracic outlet - left MRI W contrast IV
C1524574|Multisection^W contrast Intravenous:Finding:Point in time:Thoracic outlet.left:Document:MRI
C1524574|Multisection^W contrast IV:Find:Pt:Thoracic outlet.left:Doc:MRI
C1524203|Clavicle X-ray AP single view
C1524203|Clavicle XR AP 1V
C1524203|View AP:Finding:Point in time:Clavicle:Document:XR
C1524203|View AP:Find:Pt:Clavicle:Doc:XR
C1524204|Lower extremity X-ray AP single view
C1524204|LE XR AP 1V
C1524204|View AP:Find:Pt:Lower extremity:Doc:XR
C1524204|View AP:Finding:Point in time:Lower extremity:Document:XR
C1524207|Finger fourth X-ray AP single view
C1524207|Finger.4th XR AP 1V
C1524207|View AP:Find:Pt:Finger.fourth:Doc:XR
C1524207|View AP:Finding:Point in time:Finger.fourth:Document:XR
C1524284|Guidance for drainage of abscess:Find:Pt:XXX:Doc:XR.fluor
C1524284|XXX Flr Abscess drain guid
C1524284|Fluoroscopy Guidance for drainage of abscess of Unspecified body region
C1524284|Guidance for drainage of abscess:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1524300|CT Guidance for biopsy of Lymph node
C1524300|LN CT Bx guid
C1524300|Guidance for biopsy:Find:Pt:Lymph node:Doc:CT
C1524300|Guidance for biopsy:Finding:Point in time:Lymph node:Document:Computerized Tomography
C1524323|CT Guidance for drainage of Chest-- WO contrast
C1524323|Chest CT Drain guid WO contr
C1524323|Guidance for drainage^WO contrast:Find:Pt:Chest:Doc:CT
C1524323|Guidance for drainage^WO contrast:Finding:Point in time:Chest:Document:Computerized Tomography
C1524639|Ribs - bilateral X-ray 3 views
C1524639|Ribs-Bl XR 3V
C1524639|Views 3:Finding:Point in time:Ribs.bilateral:Document:XR
C1524639|Views 3:Find:Pt:Ribs.bilateral:Doc:XR
C1524993|Clavicle XR 2V
C1524993|Clavicle X-ray 2 views
C1524993|Views 2:Find:Pt:Clavicle:Doc:XR
C1524993|Views 2:Finding:Point in time:Clavicle:Document:XR
C1524355|Clavicle CT
C1524355|Multisection:Finding:Point in time:Clavicle:Document:Computerized Tomography
C1524355|Multisection:Find:Pt:Clavicle:Doc:CT
C1524374|Lower extremity - right MRI
C1524374|LE-R MRI
C1524374|Multisection:Finding:Point in time:Lower extremity.right:Document:MRI
C1524374|Multisection:Find:Pt:Lower extremity.right:Doc:MRI
C1524386|Ft-Bl CT
C1524386|Foot - bilateral CT
C1524386|Multisection:Find:Pt:Foot.bilateral:Doc:CT
C1524386|Multisection:Finding:Point in time:Foot.bilateral:Document:Computerized Tomography
C1524390|Forearm - bilateral CT
C1524390|Forearm-Bl CT
C1524390|Multisection:Find:Pt:Forearm.bilateral:Doc:CT
C1524390|Multisection:Finding:Point in time:Forearm.bilateral:Document:Computerized Tomography
C1524734|Multisection^WO & W contrast IV:Find:Pt:Forearm.left:Doc:CT
C1524734|Forearm-L CT WO+W contr IV
C1524734|Forearm - left CT WO and W contrast IV
C1524734|Multisection^WO & W contrast Intravenous:Finding:Point in time:Forearm.left:Document:Computerized Tomography
C1524744|Deprecated Calcaneus CT WO and W contrast IV
C1524744|Multisection^WO & W contrast Intravenous:Finding:Point in time:Calcaneus:Document:Computerized Tomography
C1524744|Deprecated Heel CT WO+W contr IV
C1524744|Multisection^WO & W contrast IV:Find:Pt:Calcaneus:Doc:CT
C1524753|Upper arm - left CT WO and W contrast IV
C1524753|Upper arm-L CT WO+W contr IV
C1524753|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper arm.left:Document:Computerized Tomography
C1524753|Multisection^WO & W contrast IV:Find:Pt:Upper arm.left:Doc:CT
C1525032|Femur XR AP+Lat
C1525032|Femur X-ray AP and lateral
C1525032|Views AP & lateral:Find:Pt:Femur:Doc:XR
C1525032|Views AP & lateral:Finding:Point in time:Femur:Document:XR
C1525035|Ft-Bl XR AP+Lat
C1525035|Foot - bilateral X-ray AP and lateral
C1525035|Views AP & lateral:Find:Pt:Foot.bilateral:Doc:XR
C1525035|Views AP & lateral:Finding:Point in time:Foot.bilateral:Document:XR
C1524401|Multisection:Find:Pt:Calcaneus:Doc:CT
C1524401|Deprecated Calcaneus CT
C1524401|Deprecated Heel CT
C1524401|Multisection:Finding:Point in time:Calcaneus:Document:Computerized Tomography
C1524673|L-spine XR AP+Lat+Obl
C1524673|Views AP & lateral & oblique:Find:Pt:Spine.lumbar:Doc:XR
C1524673|Views AP & lateral & oblique:Finding:Point in time:Spine.lumbar:Document:XR
C1524673|Lumbar spine X-ray AP and lateral and oblique
C1830181|Deprecated Bone density:Mass Aeric:Point in time:Radius.right+Ulna.right:Quantitative:XR.DEXA
C1830181|Bone density:MAric:Pt:Radius.right+Ulna.right:Qn:XR.DEXA
C1830181|Deprecated Radius+Ulna-R DEXA BDM
C1830181|Bone density:Mass Aeric:Point in time:Radius.right+Ulna.right:Quantitative:XR.DEXA
C1830181|Deprecated Radius & Ulna right DEXA Bone density
C1830184|Mammogram Guidance for fine needle aspiration of Breast - right
C1830184|Brst-R Mam FNA Asp
C1830184|Guidance for aspiration.fine needle:Find:Pt:Breast.right:Doc:Mam
C1830184|Guidance for aspiration.fine needle:Finding:Point in time:Breast.right:Document:Mam
C1830212|Multisection^WO & W contrast Intravenous:Finding:Point in time:Parotid gland:Document:Computerized Tomography
C1830212|Parotid gland CT WO+W contr IV
C1830212|Multisection^WO & W contrast IV:Find:Pt:Parotid gland:Doc:CT
C1830212|Parotid gland CT WO and W contrast IV
C1830083|US Guidance for needle biopsy of Ovary
C1830083|Ovary US Bx needle guid
C1830083|Guidance for biopsy.needle:Finding:Point in time:Ovary:Document:Ultrasound
C1830083|Guidance for biopsy.needle:Find:Pt:Ovary:Doc:US
C1830277|Brst Mam FNA Asp
C1830277|Mammogram Guidance for fine needle aspiration of Breast
C1830277|Guidance for aspiration.fine needle:Finding:Point in time:Breast:Document:Mam
C1830277|Guidance for aspiration.fine needle:Find:Pt:Breast:Doc:Mam
C1715401|Aorta MRI.Angio WO+W contr IV
C1715401|Multisection^WO & W contrast Intravenous:Finding:Point in time:Aorta:Document:MRI.angio
C1715401|Aorta MRI angiogram WO and W contrast IV
C1715401|Multisection^WO & W contrast IV:Find:Pt:Aorta:Doc:MRI.angio
C1717320|T+L-spine XR Scoli 1V
C1717320|View scoliosis:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1717320|View scoliosis:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1717320|Spine Thoracic and Lumbar X-ray scoliosis single view
C1645314|Maxillofacial CT
C1645314|Maxillofacial region CT
C1645314|Multisection:Find:Pt:Head>Maxillofacial region:Doc:CT
C1645314|Multisection:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1634508|Brain+Pituitary+ST MRI
C1634508|Brain and Pituitary and Sella turcica MRI
C1634508|Multisection:Find:Pt:Brain+Pituitary+Sella turcica:Doc:MRI
C1634508|Multisection:Finding:Point in time:Brain+Pituitary+Sella turcica:Document:MRI
C1714795|C+T-spine MRI
C1714795|Spine Cervical and Spine Thoracic MRI
C1714795|Multisection:Finding:Point in time:Spine.cervical+Spine.thoracic:Document:MRI
C1714795|Multisection:Find:Pt:Spine.cervical+Spine.thoracic:Doc:MRI
C1714811|BD+PDs Flr Endo guid 15m P contr retro
C1714811|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 15 minutes post contrast retrograde
C1714811|Guidance for endoscopy^15 minutes post contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1714811|Guidance for endoscopy^15M post contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1714812|BD+PDs Flr Endo guid 30M P contr retro
C1714812|Fluoroscopy Guidance for endoscopy of Biliary ducts and Pancreatic duct-- 30 minutes post contrast retrograde
C1714812|Guidance for endoscopy^30 minutes post contrast retrograde:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:XR.fluor
C1714812|Guidance for endoscopy^30M post contrast retrograde:Find:Pt:Biliary ducts+Pancreatic duct:Doc:XR.fluor
C1714529|XXX US RT fields plac guid
C1714529|US Guidance for placement of radiation therapy fields in Unspecified body region
C1714529|Guidance for placement of radiation therapy fields:Find:Pt:XXX:Doc:US
C1714529|Guidance for placement of radiation therapy fields:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1705864|Finger.3rd-L XR GE 3V
C1705864|Finger third - left X-ray GE 3 views
C1705864|Finger third - left Narrative X-ray GE 3 views
C1705864|Views GE 3:Find:Pt:Finger.third.left:Doc:XR
C1705864|Views GE 3:Finding:Point in time:Finger.third.left:Document:XR
C1714786|Liver MRI WO+W Ferumoxides IV
C1714786|Liver MRI WO and W ferumoxides IV
C1714786|Multisection^WO & W ferumoxides Intravenous:Finding:Point in time:Liver:Document:MRI
C1714786|Multisection^WO & W ferumoxides IV:Find:Pt:Liver:Doc:MRI
C1715025|Liver+Spleen RI Flow W RNC IV
C1715025|Liver and Spleen Scan flow
C1715025|Views flow^W radionuclide IV:Find:Pt:Liver+Spleen:Doc:Radnuc
C1715025|Views flow^W radionuclide Intravenous:Finding:Point in time:Liver+Spleen:Document:Radnuc
C1715102|Multisection^WO & W contrast Intravenous:Finding:Point in time:Kidney:Document:MRI
C1715102|Multisection^WO & W contrast IV:Find:Pt:Kidney:Doc:MRI
C1715102|Kidney MRI WO+W contr IV
C1715102|Kidney MRI WO and W contrast IV
C1645331|T+L-spine XR Scoli AP 1V sitting
C1645331|View scoliosis AP^sitting:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1645331|Spine Thoracic and Lumbar X-ray scoliosis AP sitting
C1645331|View scoliosis AP^sitting:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1644170|Neck X-ray AP single view
C1644170|Neck XR AP 1V
C1644170|View AP:Find:Pt:Neck:Doc:XR
C1644170|View AP:Finding:Point in time:Neck:Document:XR
C1638465|T-spine XR AP W+WO R-bending
C1638465|Views AP^W R-bending & WO bending:Find:Pt:Spine.thoracic:Doc:XR
C1638465|Views AP^W R-bending & WO bending:Finding:Point in time:Spine.thoracic:Document:XR
C1638465|Thoracic spine X-ray AP W right bending and WO bending
C1639533|Kidney ves Transplant DOP
C1639533|Kidney vessels transplant US.doppler
C1639533|Multisection:Finding:Point in time:Kidney vessels transplant:Document:Ultrasound.doppler
C1639533|Multisection:Find:Pt:Kidney vessels transplant:Doc:US.doppler
C1626767|Brst US Screening
C1626767|Breast US screening
C1626767|Multisection screening:Finding:Point in time:Breast:Document:Ultrasound
C1626767|Multisection screening:Find:Pt:Breast:Doc:US
C1627300|Breast - right FFD mammogram diagnostic
C1627300|Brst-R FFDM Dx
C1627300|Views diagnostic:Find:Pt:Breast.right:Doc:Mam.FFD
C1627300|Views diagnostic:Finding:Point in time:Breast.right:Document:Mam.FFD
C1632268|C-spine MRI W FE
C1632268|Multisection^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:MRI
C1632268|Multisection^W flexion & W extension:Find:Pt:Spine.cervical:Doc:MRI
C1632268|Cervical spine MRI W flexion and W extension
C1624129|Colon Fluoroscopy W gastrografin PR
C1624129|Colon Flr W Gastrografin PR
C1624129|Views^W gastrografin Rectal:Finding:Point in time:Colon:Document:XR.fluor
C1624129|Views^W gastrografin PR:Find:Pt:Colon:Doc:XR.fluor
C1639939|UGI Flr W Ba PO
C1639939|Gastrointestine upper Fluoroscopy W barium contrast PO
C1639939|Views^W barium contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1639939|Views^W barium contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1633389|Ribs - bilateral X-ray 2 views
C1633389|Ribs-Bl XR 2V
C1633389|Views 2:Find:Pt:Ribs.bilateral:Doc:XR
C1633389|Views 2:Finding:Point in time:Ribs.bilateral:Document:XR
C1642086|Hip-R XR AP+Lat port
C1642086|Hip - right X-ray AP and lateral portable
C1642086|Views AP & lateral portable:Find:Pt:Hip.right:Doc:XR
C1642086|Views AP & lateral portable:Finding:Point in time:Hip.right:Document:XR
C1643247|Ribs - right X-ray portable
C1643247|Ribs-R XR port
C1643247|Views portable:Find:Pt:Ribs.right:Doc:XR
C1643247|Views portable:Finding:Point in time:Ribs.right:Document:XR
C1630176|Ankle - bilateral X-ray 6 views
C1630176|Ankle-Bl XR 6V
C1630176|Views 6:Finding:Point in time:Ankle.bilateral:Document:XR
C1630176|Views 6:Find:Pt:Ankle.bilateral:Doc:XR
C1632782|Spine XR W FE
C1632782|Spine X-ray W flexion and W extension
C1632782|Views^W flexion & W extension:Finding:Point in time:Spine:Document:XR
C1632782|Views^W flexion & W extension:Find:Pt:Spine:Doc:XR
C1623596|T+L-spine XR
C1623596|Spine Thoracic and Lumbar X-ray
C1623596|Views:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1623596|Views:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1625218|C+T+L-spine MRI
C1625218|Spine Cervical and Thoracic and Lumbar MRI
C1625218|Multisection:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:MRI
C1625218|Multisection:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:MRI
C3174373|SS v+Jugular v-R XRA W contr IV
C3174373|Sagittal sinus and Jugular veins - right Fluoroscopic angiogram W contrast IV
C3174373|Views^W contrast Intravenous:Finding:Point in time:Sagittal sinus vein.right+Jugular vein.right:Document:XR.fluor.angio
C3174373|Views^W contrast IV:Find:Pt:Sagittal sinus vein.right+Jugular vein.right:Doc:XR.fluor.angio
C3262951|Fluoroscopy Guidance for needle biopsy of Salivary gland
C3262951|Salivary gland Flr Bx needle guid
C3262951|Guidance for biopsy.needle:Finding:Point in time:Salivary gland:Document:XR.fluor
C3262951|Guidance for biopsy.needle:Find:Pt:Salivary gland:Doc:XR.fluor
C3262999|Hand - bilateral MRI WO contrast
C3262999|Hand-Bl MRI WO contr
C3262999|Multisection^WO contrast:Find:Pt:Hand.bilateral:Doc:MRI
C3262999|Multisection^WO contrast:Finding:Point in time:Hand.bilateral:Document:MRI
C3483136|C-spine Flr Inj guid
C3483136|Guidance for injection:Find:Pt:Spine.cervical:Doc:XR.fluor
C3483136|Guidance for injection:Finding:Point in time:Spine.cervical:Document:XR.fluor
C3483136|Fluoroscopy Guidance for injection of Cervical spine
C3483138|T-spine Flr Inj guid
C3483138|Guidance for injection:Finding:Point in time:Spine.thoracic:Document:XR.fluor
C3483138|Guidance for injection:Find:Pt:Spine.thoracic:Doc:XR.fluor
C3483138|Fluoroscopy Guidance for injection of Thoracic spine
C3482442|T-spine US
C3482442|Multisection:Finding:Point in time:Spine.thoracic:Document:Ultrasound
C3482442|Multisection:Find:Pt:Spine.thoracic:Doc:US
C3482442|Thoracic spine US
C3263020|Guidance for biopsy.needle:Finding:Point in time:Chest>Pleura:Document:MRI
C3263020|Chest Pleura MRI Bx needle guid
C3263020|Guidance for biopsy.needle:Find:Pt:Chest>Pleura:Doc:MRI
C3263020|MRI Guidance for needle biopsy of Chest Pleura
C3263038|Fluoroscopy Guidance for needle biopsy of Chest
C3263038|Chest Flr Bx needle guid
C3263038|Guidance for biopsy.needle:Find:Pt:Chest:Doc:XR.fluor
C3263038|Guidance for biopsy.needle:Finding:Point in time:Chest:Document:XR.fluor
C3263203|Epididymis US Bx guid
C3263203|US Guidance for biopsy of Epididymis
C3263203|Guidance for biopsy:Finding:Point in time:Epididymis:Document:Ultrasound
C3263203|Guidance for biopsy:Find:Pt:Epididymis:Doc:US
C3263212|Upper extremity veins US
C3263212|UE vv US
C3263212|Multisection:Finding:Point in time:Upper extremity veins:Document:Ultrasound
C3263212|Multisection:Find:Pt:Upper extremity veins:Doc:US
C0487982|Chest X-ray Diameter.anterior-posterior W expiration
C0487982|Chest XR Diam AP W Exp
C0487982|Diameter.anterior-posterior^W expiration:Len:Pt:Chest:Qn:XR
C0487982|Diameter.anterior-posterior^W expiration:Length:Point in time:Chest:Quantitative:XR
C0487983|Diameter.anterior-posterior^W inspiration:Len:Pt:Chest:Qn:XR
C0487983|Chest XR Diam AP W Insp
C0487983|Chest X-ray Diameter.anterior-posterior W inspiration
C0487983|Diameter.anterior-posterior^W inspiration:Length:Point in time:Chest:Quantitative:XR
C0944157|Spine CT
C0944157|Multisection:Finding:Point in time:Spine:Narrative:Computerized Tomography
C0944157|Multisection:Finding:Point in time:Spine:Document:Computerized Tomography
C0944157|Multisection:Find:Pt:Spine:Doc:CT
C0942159|Radius+Ulna-L XR
C0942159|Radius - left and Ulna.left X-ray
C0942159|Views:Find:Pt:Radius.left+Ulna.left:Doc:XR
C0942159|Views:Finding:Point in time:Radius.left+Ulna.left:Document:XR
C0945317|Zygomatic arch-R XR
C0945317|Zygomatic arch - right X-ray
C0945317|Views:Finding:Point in time:Zygomatic arch.right:Document:XR
C0945317|Views:Find:Pt:Zygomatic arch.right:Doc:XR
C0945321|Multisection^WO & W contrast IV:Find:Pt:Thoracic outlet.bilateral:Doc:MRI
C0945321|Thoracic outlet - bilateral MRI WO and W contrast IV
C0945321|Multisection^WO & W contrast Intravenous:Finding:Point in time:Thoracic outlet.bilateral:Document:MRI
C0945321|TO-Bl MRI WO+W contr IV
C0942227|Extremity - left US
C0942227|Extr-L US
C0942227|Multisection:Find:Pt:Extremity.left:Doc:US
C0942227|Multisection:Finding:Point in time:Extremity.left:Document:Ultrasound
C0942321|Mammogram Guidance for core needle percutaneous biopsy of Breast - left
C0942321|Brst-L Mam PC Bx CN guid
C0942321|Guidance for percutaneous biopsy.core needle:Finding:Point in time:Breast.left:Document:Mam
C0942321|Guidance for percutaneous biopsy.core needle:Find:Pt:Breast.left:Doc:Mam
C0942343|Knee-R XR AP+PA stand
C0942343|Knee - right X-ray AP and PA standing
C0942343|Views AP & PA^standing:Find:Pt:Knee.right:Doc:XR
C0942343|Views AP & PA^standing:Finding:Point in time:Knee.right:Document:XR
C0942348|Brachiocephalic artery - left Fluoroscopic angiogram Angioplasty W contrast IA
C0942348|BrachCeph a-L XRA Angpsty W contr IA
C0942348|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Brachiocephalic artery.left:Document:XR.fluor.angio
C0942348|Angioplasty^W contrast IA:Find:Pt:Brachiocephalic artery.left:Doc:XR.fluor.angio
C0882035|Neck MRI W contr IV
C0882035|Neck MRI W contrast IV
C0882035|Multisection^W contrast Intravenous:Finding:Point in time:Neck:Document:MRI
C0882035|Multisection^W contrast IV:Find:Pt:Neck:Doc:MRI
C0882041|Orbit-Bl CT
C0882041|Orbit - bilateral CT
C0882041|Multisection:Find:Pt:Head>Orbit.bilateral:Doc:CT
C0882041|Multisection:Finding:Point in time:Head>Orbit.bilateral:Document:Computerized Tomography
C0882059|Pelvis US Drain guid
C0882059|US Guidance for drainage of Pelvis
C0882059|Guidance for drainage:Finding:Point in time:Pelvis:Document:Ultrasound
C0882059|Guidance for drainage:Find:Pt:Pelvis:Doc:US
C0882170|Tibl a XRA Angpsty W contr IA
C0882170|Tibial artery Fluoroscopic angiogram Angioplasty W contrast IA
C0882170|Angioplasty^W contrast IA:Find:Pt:Tibial artery:Doc:XR.fluor.angio
C0882170|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibial artery:Document:XR.fluor.angio
C0882180|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein
C0882180|Centl v XRA LT per cath plac guid
C0882180|Guidance for placement of longterm peripheral catheter:Finding:Point in time:Central vein:Document:XR.fluor.angio
C0882180|Guidance for placement of longterm peripheral catheter:Find:Pt:Central vein:Doc:XR.fluor.angio
C0882222|Vessel Fluoroscopic angiogram Removal of foreign body from vascular space
C0882222|Removal of foreign body from vascular space:Finding:Point in time:Vessel:Document:XR.fluor.angio
C0882222|Removal of foreign body from vascular space:Find:Pt:Vessel:Doc:XR.fluor.angio
C0882222|Vesl XRA FB rem from VS
C0942116|Ft-R XR stand
C0942116|Foot - right X-ray standing
C0942116|Views^standing:Finding:Point in time:Foot.right:Document:XR
C0942116|Views^standing:Find:Pt:Foot.right:Doc:XR
C0942142|Foot - left X-ray
C0942142|Ft-L XR
C0942142|Views:Find:Pt:Foot.left:Doc:XR
C0942142|Views:Finding:Point in time:Foot.left:Document:XR
C0881976|Multisection^W contrast IV:Find:Pt:Kidney.bilateral+Collecting system:Nar:CT
C0881976|Deprecated KD-Bl+CS CT W contr IV
C0881976|Multisection^W contrast Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:Computerized Tomography
C0881976|Deprecated Kidney - bilateral and Collecting system CT W contrast IV
C0881980|Views^W contrast via nephrostomy tube:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C0881980|Views^W contrast via nephrostomy tube:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C0881980|Kidney - bilateral Fluoroscopy W contrast via nephrostomy tube
C0881980|Kdny-Bl Flr W contr via NT
C2608057|Views^W contrast Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:XR
C2608057|Views^W contrast IV:Find:Pt:Kidney.bilateral:Doc:XR
C2608057|Kidney - bilateral X-ray W contrast IV
C2608057|Views^W contrast Intravenous:Finding:Point in time:Kidney.bilateral:Document:XR
C2608057|Kdny-Bl XR W contr IV
C1114543|C-spine.odontoidaxis XR AP V1 port
C1114543|Spine Cervical Odontoid and Cervical axis X-ray AP portable single view
C1114543|View AP portable:Finding:Point in time:Spine.cervical.odontoid+Spine.cervical.axis:Document:XR
C1114543|View AP portable:Find:Pt:Spine.cervical.odontoid+Spine.cervical.axis:Doc:XR
C1114577|Pelvis X-ray portable
C1114577|Pelvis XR port
C1114577|Views portable:Finding:Point in time:Pelvis:Document:XR
C1114577|Views portable:Find:Pt:Pelvis:Doc:XR
C1114620|Carotid artery.external - bilateral Fluoroscopic angiogram W contrast IA
C1114620|Carot a.ext-Bl XRA W contr IA
C1114620|Views^W contrast IA:Find:Pt:Carotid artery.external.bilateral:Doc:XR.fluor.angio
C1114620|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.external.bilateral:Document:XR.fluor.angio
C1526820|Carot a.Int-L XRA W contr IA
C1526820|Carotid artery.internal - left Fluoroscopic angiogram W contrast IA
C1526820|Views^W contrast IA:Find:Pt:Carotid artery.internal.left:Doc:XR.fluor.angio
C1526820|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.internal.left:Document:XR.fluor.angio
C1543424|Should-Bl XR AP+Ax+Outlet+30 Deg Cau
C1543424|Shoulder - bilateral X-ray AP and axillary and outlet and 30 degree caudal angle
C1543424|Views AP & axillary & outlet & 30 degree caudal angle:Find:Pt:Shoulder.bilateral:Doc:XR
C1543424|Views AP & axillary & outlet & 30 degree caudal angle:Finding:Point in time:Shoulder.bilateral:Document:XR
C1543755|Hrt RI PF W DBM+RNC IV
C1543755|Heart Scan perfusion W dobutamine and W radionuclide IV
C1543755|Views perfusion^W dobutamine & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543755|Views perfusion^W dobutamine & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543760|Hrt RI PF W DPY+RNC IV
C1543760|Heart Scan perfusion W dipyridamole and W radionuclide IV
C1543760|Views perfusion^W dipyridamole & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543760|Views perfusion^W dipyridamole & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543463|Knee - right X-ray 3 views and Sunrise
C1543463|Knee-R XR 3V+Sunrise
C1543463|Views 3 & Sunrise:Find:Pt:Knee.right:Doc:XR
C1543463|Views 3 & Sunrise:Finding:Point in time:Knee.right:Document:XR
C1543484|T-spine XR 5V+Obl
C1543484|Views 5 & oblique:Finding:Point in time:Spine.thoracic:Document:XR
C1543484|Views 5 & oblique:Find:Pt:Spine.thoracic:Doc:XR
C1543484|Thoracic spine X-ray 5 views and oblique
C1542848|Thyroid RI W Tc99mIV
C1542848|Thyroid Scan W Tc-99m IV
C1542848|Views^W Tc-99m IV:Find:Pt:Thyroid:Doc:Radnuc
C1542848|Views^W Tc-99m Intravenous:Finding:Point in time:Thyroid:Document:Radnuc
C1542904|RI Delayed W In-111 Satmb IV
C1542904|Scan delayed W In-111 Satumomab IV
C1542904|Views delayed^W In-111 Satumomab IV:Find:Pt:^Patient:Doc:Radnuc
C1542904|Views delayed^W In-111 Satumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542922|Hrt RI FP Rest+W RNC IV
C1542922|Heart Scan first pass at rest and W radionuclide IV
C1542922|Views first pass^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1542922|Views first pass^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543935|Hrt SPECT Gated+EF W RNC IV
C1543935|Heart SPECT gated and ejection fraction
C1543935|Multisection gated & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543935|Multisection gated & ejection fraction^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543936|Hrt RI Gated W Tc99mMIBI IV
C1543936|Heart Scan gated W Tc-99m Sestamibi IV
C1543936|Views gated^W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543936|Views gated^W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543965|Scrotum+Test RI Static+Flow W RNC IV
C1543965|Scrotum and Testicle Scan static and flow
C1543965|Views static & flow^W radionuclide IV:Find:Pt:Scrotum+Testicle:Doc:Radnuc
C1543965|Views static & flow^W radionuclide Intravenous:Finding:Point in time:Scrotum+Testicle:Document:Radnuc
C1543496|Lower extremity vein - bilateral US.doppler
C1543496|LE v-Bl DOP
C1543496|Multisection:Find:Pt:Lower extremity vein.bilateral:Doc:US.doppler
C1543496|Multisection:Finding:Point in time:Lower extremity vein.bilateral:Document:Ultrasound.doppler
C1543163|Extremity artery US.doppler
C1543163|Extr a DOP
C1543163|Multisection:Finding:Point in time:Extremity artery:Document:Ultrasound.doppler
C1543163|Multisection:Find:Pt:Extremity artery:Doc:US.doppler
C1543196|Toes XR AP+Obl
C1543196|Toes X-ray AP and oblique
C1543196|Views AP & oblique:Finding:Point in time:Toes:Document:XR
C1543196|Views AP & oblique:Find:Pt:Toes:Doc:XR
C1543599|Vein US.doppler limited
C1543599|Vein DOP Ltd
C1543599|Multisection limited:Finding:Point in time:Vein:Document:Ultrasound.doppler
C1543599|Multisection limited:Find:Pt:Vein:Doc:US.doppler
C1526752|Hip-R XR port
C1526752|Hip - right X-ray portable
C1526752|Views portable:Find:Pt:Hip.right:Doc:XR
C1526752|Views portable:Finding:Point in time:Hip.right:Document:XR
C1524435|Maxilla CT
C1524435|Multisection:Find:Pt:Maxilla:Doc:CT
C1524435|Multisection:Finding:Point in time:Maxilla:Document:Computerized Tomography
C1524849|Femur - right CT WO contrast
C1524849|Femur-R CT WO contr
C1524849|Multisection^WO contrast:Finding:Point in time:Femur.right:Document:Computerized Tomography
C1524849|Multisection^WO contrast:Find:Pt:Femur.right:Doc:CT
C1524457|Multisection limited^WO & W contrast Intravenous:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524457|Multisection limited^WO & W contrast IV:Find:Pt:Abdomen:Doc:CT
C1524457|Abdomen CT limited WO and W contrast IV
C1524457|Abd CT Ltd WO+W contr IV
C1525297|Hand XR Ball Catcher
C1525297|Hand X-ray Ball Catcher
C1525297|View Ball Catcher:Find:Pt:Hand:Doc:XR
C1525297|View Ball Catcher:Finding:Point in time:Hand:Document:XR
C1525240|Temporal bone CT WO contr
C1525240|Temporal bone CT WO contrast
C1525240|Multisection^WO contrast:Finding:Point in time:Temporal bone:Document:Computerized Tomography
C1525240|Multisection^WO contrast:Find:Pt:Temporal bone:Doc:CT
C1525250|Neck vv MRI.Angio WO contr
C1525250|Neck veins MRI angiogram WO contrast
C1525250|Multisection^WO contrast:Find:Pt:Neck veins:Doc:MRI.angio
C1525250|Multisection^WO contrast:Finding:Point in time:Neck veins:Document:MRI.angio
C1525277|Knee - bilateral X-ray 2 views standing
C1525277|Knee-Bl XR 2V stand
C1525277|Views 2^standing:Finding:Point in time:Knee.bilateral:Document:XR
C1525277|Views 2^standing:Find:Pt:Knee.bilateral:Doc:XR
C1525497|Hip XR AP+Lat Xtable
C1525497|Hip X-ray AP and lateral crosstable
C1525497|Views AP & lateral crosstable:Find:Pt:Hip:Doc:XR
C1525497|Views AP & lateral crosstable:Finding:Point in time:Hip:Document:XR
C1525504|Hip-L XR AP+Lat Frog
C1525504|Hip - left X-ray AP and lateral frog
C1525504|Views AP & lateral frog:Finding:Point in time:Hip.left:Document:XR
C1525504|Views AP & lateral frog:Find:Pt:Hip.left:Doc:XR
C1524247|C-spine XR AP+Lat+Obl+Odont
C1524247|Views AP & lateral & oblique & odontoid:Finding:Point in time:Spine.cervical:Document:XR
C1524247|Views AP & lateral & oblique & odontoid:Find:Pt:Spine.cervical:Doc:XR
C1524247|Cervical spine X-ray AP and lateral and oblique and odontoid
C1524249|L-spine XR AP+Lat+Obl+Spot
C1524249|Views AP & lateral & oblique & spot:Find:Pt:Spine.lumbar:Doc:XR
C1524249|Views AP & lateral & oblique & spot:Finding:Point in time:Spine.lumbar:Document:XR
C1524249|Lumbar spine X-ray AP and lateral and oblique and spot
C1525522|Should-L XR AP+Stryker Notch
C1525522|Shoulder - left X-ray AP and Stryker Notch
C1525522|Views AP & Stryker Notch:Finding:Point in time:Shoulder.left:Document:XR
C1525522|Views AP & Stryker Notch:Find:Pt:Shoulder.left:Doc:XR
C1525549|Chest XR PA+R-Obl+L-Obl
C1525549|Chest X-ray PA and right oblique and left oblique
C1525549|Views PA & R-oblique & L-oblique:Finding:Point in time:Chest:Document:XR
C1525549|Views PA & R-oblique & L-oblique:Find:Pt:Chest:Doc:XR
C1525571|Coronary arteries Fluoroscopic angiogram W contrast IA
C1525571|Coronary aa XRA W contr IA
C1525571|Views^W contrast Intra-arterial:Finding:Point in time:Coronary arteries:Document:XR.fluor.angio
C1525571|Views^W contrast IA:Find:Pt:Coronary arteries:Doc:XR.fluor.angio
C1525575|Iliac a-L XRA W contr IA
C1525575|Iliac artery - left Fluoroscopic angiogram W contrast IA
C1525575|Views^W contrast Intra-arterial:Finding:Point in time:Iliac artery.left:Document:XR.fluor.angio
C1525575|Views^W contrast IA:Find:Pt:Iliac artery.left:Doc:XR.fluor.angio
C1525597|Ankle X-ray standing
C1525597|Ankle XR stand
C1525597|Views^standing:Finding:Point in time:Ankle:Document:XR
C1525597|Views^standing:Find:Pt:Ankle:Doc:XR
C1525636|SC joint CT W contr IV
C1525636|Sternoclavicular Joint CT W contrast IV
C1525636|Multisection^W contrast Intravenous:Finding:Point in time:Sternoclavicular joint:Document:Computerized Tomography
C1525636|Multisection^W contrast IV:Find:Pt:Sternoclavicular joint:Doc:CT
C1525639|TMJ-Bl MRI W contr IV
C1525639|Temporomandibular joint - bilateral MRI W contrast IV
C1525639|Multisection^W contrast IV:Find:Pt:Temporomandibular joint.bilateral:Doc:MRI
C1525639|Multisection^W contrast Intravenous:Finding:Point in time:Temporomandibular joint.bilateral:Document:MRI
C1525690|L-spine+Sacrum+Coccyx XR
C1525690|Spine Lumbar and Sacrum and Coccyx X-ray
C1525690|Views:Find:Pt:Spine.lumbar+Sacrum+Coccyx:Doc:XR
C1525690|Views:Finding:Point in time:Spine.lumbar+Sacrum+Coccyx:Document:XR
C1525738|LE vv-Bl XRA W contr IV
C1525738|Lower extremity veins - bilateral Fluoroscopic angiogram W contrast IV
C1525738|Views^W contrast Intravenous:Finding:Point in time:Lower extremity veins.bilateral:Document:XR.fluor.angio
C1525738|Views^W contrast IV:Find:Pt:Lower extremity veins.bilateral:Doc:XR.fluor.angio
C1525767|Wrist MRI WO contr
C1525767|Wrist MRI WO contrast
C1525767|Multisection^WO contrast:Finding:Point in time:Wrist:Document:MRI
C1525767|Multisection^WO contrast:Find:Pt:Wrist:Doc:MRI
C1525774|AC joint XR 10 Deg Ceph Angle
C1525774|Acromioclavicular Joint X-ray 10 degree cephalic angle
C1525774|View 10 degree cephalic angle:Finding:Point in time:Acromioclavicular joint:Document:XR
C1525774|View 10 degree cephalic angle:Find:Pt:Acromioclavicular joint:Doc:XR
C1525851|Wrist-L XR Ulnar+Radial Deviation
C1525851|Wrist - left X-ray ulnar deviation and radial deviation
C1525851|Views ulnar deviation & radial deviation:Find:Pt:Wrist.left:Doc:XR
C1525851|Views ulnar deviation & radial deviation:Finding:Point in time:Wrist.left:Document:XR
C1525879|Pelvis+Hip-Bl XR +Lat Frog
C1525879|Pelvis and Hip - bilateral X-ray and lateral frog
C1525879|Views & lateral frog:Finding:Point in time:Pelvis+Hip.bilateral:Document:XR
C1525879|Views & lateral frog:Find:Pt:Pelvis+Hip.bilateral:Doc:XR
C1524137|Ac arch+Carot a+VA XRA W contr IA
C1524137|Aortic arch and Carotid artery and Vertebral artery Fluoroscopic angiogram W contrast IA
C1524137|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery+Vertebral artery:Doc:XR.fluor.angio
C1524137|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery+Vertebral artery:Document:XR.fluor.angio
C1525834|Should-L XR Grashey+Ax+ Y
C1525834|Shoulder - left X-ray Grashey and axillary and Y
C1525834|Views Grashey & axillary & Y:Find:Pt:Shoulder.left:Doc:XR
C1525834|Views Grashey & axillary & Y:Finding:Point in time:Shoulder.left:Document:XR
C1525969|Sacrum XR AP+Lat
C1525969|Sacrum X-ray AP and lateral
C1525969|Views AP & lateral:Finding:Point in time:Sacrum:Document:XR
C1525969|Views AP & lateral:Find:Pt:Sacrum:Doc:XR
C1526004|Elbow - right X-ray tomograph
C1526004|Elbow-R XRTomo
C1526004|Multisection:Find:Pt:Elbow.right:Doc:XR.tomo
C1526004|Multisection:Finding:Point in time:Elbow.right:Document:XR.tomo
C1526116|Shoulder - right X-ray tomograph
C1526116|Should-R XRTomo
C1526116|Multisection:Finding:Point in time:Shoulder.right:Document:XR.tomo
C1526116|Multisection:Find:Pt:Shoulder.right:Doc:XR.tomo
C1526128|Toes-R XR stand
C1526128|Toes - right X-ray standing
C1526128|Views^standing:Find:Pt:Toes.right:Doc:XR
C1526128|Views^standing:Finding:Point in time:Toes.right:Document:XR
C1526038|Hip-R XR 3V
C1526038|Hip - right X-ray 3 views
C1526038|Views 3:Find:Pt:Hip.right:Doc:XR
C1526038|Views 3:Finding:Point in time:Hip.right:Document:XR
C1526054|Humerus-R XR
C1526054|Humerus - right X-ray
C1526054|Views:Find:Pt:Humerus.right:Doc:XR
C1526054|Views:Finding:Point in time:Humerus.right:Document:XR
C1526064|Knee-R XR AP+Lat+Obl
C1526064|Knee - right X-ray AP and lateral and oblique
C1526064|Views AP & lateral & oblique:Find:Pt:Knee.right:Doc:XR
C1526064|Views AP & lateral & oblique:Finding:Point in time:Knee.right:Document:XR
C1526095|Scapula - right X-ray Y
C1526095|Scapula-R XR Y
C1526095|View Y:Finding:Point in time:Scapula.right:Document:XR
C1526095|View Y:Find:Pt:Scapula.right:Doc:XR
C1526209|Adrenal a-R XRA W contr IA
C1526209|Adrenal artery - right Fluoroscopic angiogram W contrast IA
C1526209|Views^W contrast Intra-arterial:Finding:Point in time:Adrenal artery.right:Document:XR.fluor.angio
C1526209|Views^W contrast IA:Find:Pt:Adrenal artery.right:Doc:XR.fluor.angio
C1526210|Adrenal v-R XRA W contr IV
C1526210|Adrenal vein - right Fluoroscopic angiogram W contrast IV
C1526210|Views^W contrast Intravenous:Finding:Point in time:Adrenal vein.right:Document:XR.fluor.angio
C1526210|Views^W contrast IV:Find:Pt:Adrenal vein.right:Doc:XR.fluor.angio
C1526224|Renal v-R XRA W contr IV
C1526224|Renal vein - right Fluoroscopic angiogram W contrast IV
C1526224|Views^W contrast Intravenous:Finding:Point in time:Renal vein.right:Document:XR.fluor.angio
C1526224|Views^W contrast IV:Find:Pt:Renal vein.right:Doc:XR.fluor.angio
C1525138|US Guidance for aspiration of cyst of Breast - bilateral
C1525138|Brst-Bl US Cyst Asp guid
C1525138|Guidance for aspiration of cyst:Finding:Point in time:Breast.bilateral:Document:Ultrasound
C1525138|Guidance for aspiration of cyst:Find:Pt:Breast.bilateral:Doc:US
C1526284|Lower extremity - right US
C1526284|LE-R US
C1526284|Multisection:Find:Pt:Lower extremity.right:Doc:US
C1526284|Multisection:Finding:Point in time:Lower extremity.right:Document:Ultrasound
C1525149|Finger.4th-R XR
C1525149|Finger fourth - right X-ray
C1525149|Views:Find:Pt:Finger.fourth.right:Doc:XR
C1525149|Views:Finding:Point in time:Finger.fourth.right:Document:XR
C1526308|Knee XR Merchants 30+45+60 Deg
C1526308|Knee X-ray Merchants 30 and 45 and 60 degrees
C1526308|Views Merchants 30 & 45 & 60 degrees:Find:Pt:Knee:Doc:XR
C1526308|Views Merchants 30 & 45 & 60 degrees:Finding:Point in time:Knee:Document:XR
C1526325|Knee-R XR 2V Obl
C1526325|Knee - right X-ray 2 views Oblique
C1526325|Views 2 oblique:Find:Pt:Knee.right:Doc:XR
C1526325|Views 2 oblique:Finding:Point in time:Knee.right:Document:XR
C1524511|LE-R MRI W contr IV
C1524511|Lower extremity - right MRI W contrast IV
C1524511|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.right:Document:MRI
C1524511|Multisection^W contrast IV:Find:Pt:Lower extremity.right:Doc:MRI
C1524903|Posterior fossa MRI WO contrast
C1524903|Post fossa MRI WO contr
C1524903|Multisection^WO contrast:Find:Pt:Posterior fossa:Doc:MRI
C1524903|Multisection^WO contrast:Finding:Point in time:Posterior fossa:Document:MRI
C1524910|Sternum CT WO contr
C1524910|Sternum CT WO contrast
C1524910|Multisection^WO contrast:Finding:Point in time:Sternum:Document:Computerized Tomography
C1524910|Multisection^WO contrast:Find:Pt:Sternum:Doc:CT
C1524922|Superior vena cava MRI WO contrast
C1524922|SVC MRI WO contr
C1524922|Multisection^WO contrast:Finding:Point in time:Vena cava.superior:Document:MRI
C1524922|Multisection^WO contrast:Find:Pt:Vena cava.superior:Doc:MRI
C1524932|Lower extremity - left X-ray Single view
C1524932|LE-L XR 1V
C1524932|View 1:Finding:Point in time:Lower extremity.left:Document:XR
C1524932|View 1:Find:Pt:Lower extremity.left:Doc:XR
C1524940|Ankle X-ray lateral
C1524940|Ankle XR Lat
C1524940|View lateral:Finding:Point in time:Ankle:Document:XR
C1524940|View lateral:Find:Pt:Ankle:Doc:XR
C1524619|Abdomen X-ray 3 views
C1524619|Abd XR 3V
C1524619|Views 3:Find:Pt:Abdomen:Doc:XR
C1524619|Views 3:Finding:Point in time:Abdomen:Document:XR
C1524951|Hip - left X-ray lateral
C1524951|Hip-L XR Lat
C1524951|View lateral:Finding:Point in time:Hip.left:Document:XR
C1524951|View lateral:Find:Pt:Hip.left:Doc:XR
C1524967|Knee X-ray oblique
C1524967|Knee XR Obl
C1524967|Views oblique:Find:Pt:Knee:Doc:XR
C1524967|Views oblique:Finding:Point in time:Knee:Document:XR
C1524968|Chest X-ray left anterior oblique
C1524968|Chest XR L-Ant Obl
C1524968|View L-anterior oblique:Find:Pt:Chest:Doc:XR
C1524968|View L-anterior oblique:Finding:Point in time:Chest:Document:XR
C1524625|Elbow XR 3V
C1524625|Elbow X-ray 3 views
C1524625|Views 3:Find:Pt:Elbow:Doc:XR
C1524625|Views 3:Finding:Point in time:Elbow:Document:XR
C1524655|Shoulder - bilateral X-ray 4 views
C1524655|Should-Bl XR 4V
C1524655|Views 4:Finding:Point in time:Shoulder.bilateral:Document:XR
C1524655|Views 4:Find:Pt:Shoulder.bilateral:Doc:XR
C1524161|Hip XR 2V
C1524161|Hip X-ray 2 views
C1524161|Views 2:Find:Pt:Hip:Doc:XR
C1524161|Views 2:Finding:Point in time:Hip:Document:XR
C1524365|LE CT
C1524365|Lower extremity CT
C1524365|Multisection:Finding:Point in time:Lower extremity:Document:Computerized Tomography
C1524365|Multisection:Find:Pt:Lower extremity:Doc:CT
C1524377|Upper extremity - right CT
C1524377|UE-R CT
C1524377|Multisection:Find:Pt:Upper extremity.right:Doc:CT
C1524377|Multisection:Finding:Point in time:Upper extremity.right:Document:Computerized Tomography
C1524389|Ft-R CT
C1524389|Foot - right CT
C1524389|Multisection:Find:Pt:Foot.right:Doc:CT
C1524389|Multisection:Finding:Point in time:Foot.right:Document:Computerized Tomography
C1524738|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hand:Document:Computerized Tomography
C1524738|Multisection^WO & W contrast IV:Find:Pt:Hand:Doc:CT
C1524738|Hand CT WO and W contrast IV
C1524738|Hand CT WO+W contr IV
C1524741|Multisection^WO & W contrast IV:Find:Pt:Hand.right:Doc:CT
C1524741|Hand - right CT WO and W contrast IV
C1524741|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hand.right:Document:Computerized Tomography
C1524741|Hand-R CT WO+W contr IV
C1524418|Upper arm-R CT
C1524418|Upper arm - right CT
C1524418|Multisection:Finding:Point in time:Upper arm.right:Document:Computerized Tomography
C1524418|Multisection:Find:Pt:Upper arm.right:Doc:CT
C1524779|Scapula - right MRI WO and W contrast IV
C1524779|Multisection^WO & W contrast Intravenous:Finding:Point in time:Scapula.right:Document:MRI
C1524779|Multisection^WO & W contrast IV:Find:Pt:Scapula.right:Doc:MRI
C1524779|Scapula-R MRI WO+W contr IV
C1524796|Lower leg - right CT WO and W contrast IV
C1524796|Multisection^WO & W contrast IV:Find:Pt:Lower leg.right:Doc:CT
C1524796|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower leg.right:Document:Computerized Tomography
C1524796|Lower leg-R CT WO+W contr IV
C1525068|Ft-Bl XR AP+Lat+Obl
C1525068|Foot - bilateral X-ray AP and lateral and oblique
C1525068|Views AP & lateral & oblique:Find:Pt:Foot.bilateral:Doc:XR
C1525068|Views AP & lateral & oblique:Finding:Point in time:Foot.bilateral:Document:XR
C1525078|Chest XR PA+AP Lat-Decub
C1525078|Chest X-ray PA and AP lateral-decubitus
C1525078|Views PA & AP lateral-decubitus:Find:Pt:Chest:Doc:XR
C1525078|Views PA & AP lateral-decubitus:Finding:Point in time:Chest:Document:XR
C1830180|Hip - right DXA Bone density
C1830180|Bone density:MAric:Pt:Hip.right:Qn:XR.DXA
C1830180|Bone density:Mass Aeric:Point in time:Hip.right:Quantitative:XR.DXA
C1830180|Hip-R DXA BDM
C1830208|LE.R-ves CT.Angio WO+W contr IV
C1830208|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.right>Vessels:Doc:CT.angio
C1830208|Lower extremity - right Vessels CT angiogram WO and W contrast IV
C1830208|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.right>Vessels:Document:Computerized Tomography.angio
C1830216|Maxillofacial CT WO+W red contr vol IV
C1830216|Maxillofacial region CT WO and W reduced contrast volume IV
C1830216|Multisection^WO & W reduced contrast volume Intravenous:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1830216|Multisection^WO & W reduced contrast volume IV:Find:Pt:Head>Maxillofacial region:Doc:CT
C1830260|Superior mesenteric vessels MRI angiogram
C1830260|SM ves MRI.Angio
C1830260|Multisection:Find:Pt:Superior mesenteric vessels:Doc:MRI.angio
C1830260|Multisection:Finding:Point in time:Superior mesenteric vessels:Document:MRI.angio
C1715400|Ac arch MRI.Angio WO contr
C1715400|Aortic arch MRI angiogram WO contrast
C1715400|Multisection^WO contrast:Finding:Point in time:Aortic arch:Document:MRI.angio
C1715400|Multisection^WO contrast:Find:Pt:Aortic arch:Doc:MRI.angio
C1715420|Brain SPECT W Tc99mBicisate IV
C1715420|Brain SPECT W Tc-99m bicisate IV
C1715420|Multisection^W Tc-99m bicisate IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1715420|Multisection^W Tc-99m bicisate Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1715451|Ft XR AP+Lat port
C1715451|Foot X-ray AP and lateral portable
C1715451|Views AP & lateral portable:Find:Pt:Foot:Doc:XR
C1715451|Views AP & lateral portable:Finding:Point in time:Foot:Document:XR
C1715456|Pelvis X-ray GE 3 Portable views
C1715456|Pelvis XR GE 3V Port
C1715456|Views GE 3 portable:Finding:Point in time:Pelvis:Document:XR
C1715456|Views GE 3 portable:Find:Pt:Pelvis:Doc:XR
C1715472|Chest X-ray GE 4 views
C1715472|Chest XR GE 4V
C1715472|Views GE 4:Find:Pt:Chest:Doc:XR
C1715472|Views GE 4:Finding:Point in time:Chest:Document:XR
C1643597|Multisection^W radionuclide Intravenous:Finding:Point in time:Bone:Narrative:Radnuc.SPECT
C1643597|Multisection^W radionuclide IV:Find:Pt:Bone:Nar:Radnuc.SPECT
C1643597|Deprecated Bone SPECT W RNC IV
C1643597|Deprecated Bone SPECT
C1644149|Upper extremity artery US limited
C1644149|UE a US Ltd
C1644149|Multisection limited:Finding:Point in time:Upper extremity artery:Document:Ultrasound
C1644149|Multisection limited:Find:Pt:Upper extremity artery:Doc:US
C1644150|Hip-L XR AP+Lat port
C1644150|Hip - left X-ray AP and lateral portable
C1644150|Views AP & lateral portable:Find:Pt:Hip.left:Doc:XR
C1644150|Views AP & lateral portable:Finding:Point in time:Hip.left:Document:XR
C1706624|Finger fourth - right X-ray GE 3 views
C1706624|Finger.4th-R XR GE 3V
C1706624|Finger fourth - right Narrative X-ray GE 3 views
C1706624|Views GE 3:Finding:Point in time:Finger.fourth.right:Document:XR
C1706624|Views GE 3:Find:Pt:Finger.fourth.right:Doc:XR
C1717247|CT Guidance for percutaneous drainage of abscess of Unspecified body region
C1717247|XXX CT PC Abscess Drain guid
C1717247|Guidance for percutaneous drainage of abscess:Find:Pt:XXX:Doc:CT
C1717247|Guidance for percutaneous drainage of abscess:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1715093|Carotid artery - bilateral US.doppler
C1715093|Carot a-Bl DOP
C1715093|Multisection:Find:Pt:Carotid artery.bilateral:Doc:US.doppler
C1715093|Multisection:Finding:Point in time:Carotid artery.bilateral:Document:Ultrasound.doppler
C1715119|Tibioperoneal arteries Fluoroscopic angiogram Angioplasty W contrast IA
C1715119|Tibioperon aa XRA Angpsty W contr IA
C1715119|Angioplasty^W contrast IA:Find:Pt:Tibioperoneal arteries:Doc:XR.fluor.angio
C1715119|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibioperoneal arteries:Document:XR.fluor.angio
C1636067|Views AP^WO & W R-bending:Find:Pt:Spine.lumbar:Doc:XR
C1636067|Views AP^WO & W R-bending:Finding:Point in time:Spine.lumbar:Document:XR
C1636067|L-spine XR AP WO+W R-bending
C1636067|Lumbar spine X-ray AP W and WO right bending
C1637231|Sinuses X-ray Waters stereo
C1637231|Sinuses XR Waters Stereo
C1637231|View Waters stereo:Find:Pt:Sinuses:Doc:XR
C1637231|View Waters stereo:Finding:Point in time:Sinuses:Document:XR
C1642068|US Guidance for biopsy of Mediastinum
C1642068|Mediastinum US Bx guid
C1642068|Guidance for biopsy:Finding:Point in time:Mediastinum:Document:Ultrasound
C1642068|Guidance for biopsy:Find:Pt:Mediastinum:Doc:US
C1639386|Carotid artery - right US limited
C1639386|Carot a-R US Ltd
C1639386|Multisection limited:Finding:Point in time:Carotid artery.right:Document:Ultrasound
C1639386|Multisection limited:Find:Pt:Carotid artery.right:Doc:US
C1626769|Hrt RI W DBM+RNC IV
C1626769|Heart Scan W dobutamine and W radionuclide IV
C1626769|Views^W dobutamine & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1626769|Views^W dobutamine & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1643243|Pelvis+Hip-R XR AP+Lat Frog Port
C1643243|Pelvis and Hip - right X-ray AP and lateral frog portable
C1643243|Views AP & lateral frog portable:Find:Pt:Pelvis+Hip.right:Doc:XR
C1643243|Views AP & lateral frog portable:Finding:Point in time:Pelvis+Hip.right:Document:XR
C1633447|Multisection^WO & W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:MRI
C1633447|XXX MRI WO+W contr IV
C1633447|Unspecified body region MRI WO and W contrast IV
C1633447|Multisection^WO & W contrast IV:Find:Pt:XXX:Doc:MRI
C1645328|Multisection^WO & W contrast IV:Find:Pt:Clavicle:Doc:MRI
C1645328|Clavicle MRI WO and W contrast IV
C1645328|Multisection^WO & W contrast Intravenous:Finding:Point in time:Clavicle:Document:MRI
C1645328|Clavicle MRI WO+W contr IV
C1632227|Hrt RI Gated+WM W RNC IV
C1632227|Heart Scan gated and wall motion
C1632227|Views gated & wall motion^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1632227|Views gated & wall motion^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1632262|Bladder+Urethra MRI Cine
C1632262|Urinary Bladder and Urethra MRI cine
C1632262|Multisection cine:Find:Pt:Urinary bladder+Urethra:Doc:MRI
C1632262|Multisection cine:Finding:Point in time:Urinary bladder+Urethra:Document:MRI
C1954301|Skull.base MRI WO contr
C1954301|Skull.base MRI WO contrast
C1954301|Multisection^WO contrast:Finding:Point in time:Skull.base:Document:MRI
C1954301|Multisection^WO contrast:Find:Pt:Skull.base:Doc:MRI
C1954312|Submandibular gland - bilateral Fluoroscopy W contrast intra salivary duct
C1954312|Views^W contrast intra salivary duct:Finding:Point in time:Submandibular gland.bilateral:Document:XR.fluor
C1954312|Views^W contrast intra salivary duct:Find:Pt:Submandibular gland.bilateral:Doc:XR.fluor
C1954312|Submandib gland-Bl Flr W contr intra SD
C1953944|Deprecated Multisection^WO contrast:Finding:Point in time:Temporal bones:Narrative:MRI
C1953944|Deprecated Temporal bones MRI W contr IV
C1953944|Multisection^WO contrast:Finding:Point in time:Temporal bone:Narrative:MRI
C1953944|Multisection^WO contrast:Find:Pt:Temporal bone:Nar:MRI
C1953947|Multisection^WO & W contrast Intrathecal:Finding:Point in time:Spine.thoracic:Document:MRI
C1953947|Multisection^WO & W contrast IT:Find:Pt:Spine.thoracic:Doc:MRI
C1953947|T-spine MRI WO+W contr IT
C1953947|Thoracic spine MRI WO and W contrast IT
C1953949|Nasoph CT WO+W contr IV
C1953949|Multisection^WO & W contrast IV:Find:Pt:Nasopharynx:Doc:CT
C1953949|Nasopharynx CT WO and W contrast IV
C1953949|Multisection^WO & W contrast Intravenous:Finding:Point in time:Nasopharynx:Document:Computerized Tomography
C1953968|Knee - left X-ray AP single view
C1953968|Knee-L XR AP 1V
C1953968|View AP:Finding:Point in time:Knee.left:Document:XR
C1953968|View AP:Find:Pt:Knee.left:Doc:XR
C1953982|Hand-Bl XR AP+Lat
C1953982|Hand - bilateral X-ray AP and lateral
C1953982|Views AP & lateral:Finding:Point in time:Hand.bilateral:Document:XR
C1953982|Views AP & lateral:Find:Pt:Hand.bilateral:Doc:XR
C3174372|Sagittal sinus vein - right Fluoroscopic angiogram W contrast IV
C3174372|SS v-R XRA W contr IV
C3174372|Views^W contrast Intravenous:Finding:Point in time:Sagittal sinus vein.right:Document:XR.fluor.angio
C3174372|Views^W contrast IV:Find:Pt:Sagittal sinus vein.right:Doc:XR.fluor.angio
C3533481|Guidance for injection of sclerosing agent:Find:Pt:Extremity veins.right:Doc:US
C3533481|Guidance for injection of sclerosing agent:Finding:Point in time:Extremity veins.right:Document:Ultrasound
C3533481|Extr vv-R US Sclerosing agent inj guid
C3533481|US Guidance for injection of sclerosing agent of Extremity veins - right
C3533797|Multisection^WO contrast:Find:Pt:Facial bones:Doc:CT
C3533797|Face CT WO contr
C3533797|Facial bones CT WO contrast
C3533797|Multisection^WO contrast:Finding:Point in time:Facial bones:Document:Computerized Tomography
C3262984|Ankle - bilateral MRI WO contrast
C3262984|Ankle-Bl MRI WO contr
C3262984|Multisection^WO contrast:Finding:Point in time:Ankle.bilateral:Document:MRI
C3262984|Multisection^WO contrast:Find:Pt:Ankle.bilateral:Doc:MRI
C3263002|Upper arm - bilateral MRI W contrast IV
C3263002|Upper arm-Bl MRI W contr IV
C3263002|Multisection^W contrast Intravenous:Finding:Point in time:Upper arm.bilateral:Document:MRI
C3263002|Multisection^W contrast IV:Find:Pt:Upper arm.bilateral:Doc:MRI
C3263035|VC MRI
C3263035|Vena cava MRI
C3263035|Multisection:Finding:Point in time:Vena cava:Document:MRI
C3263035|Multisection:Find:Pt:Vena cava:Doc:MRI
C3263046|Parotid gland Scan W Tc-99m pertechnetate IV
C3263046|Parotid gland RI W Tc99mP IV
C3263046|Views^W Tc-99m pertechnetate Intravenous:Finding:Point in time:Parotid gland:Document:Radnuc
C3263046|Views^W Tc-99m pertechnetate IV:Find:Pt:Parotid gland:Doc:Radnuc
C3484381|Knee-R XR Sunrise
C3484381|Knee - right X-ray Sunrise
C3484381|View Sunrise:Finding:Point in time:Knee.right:Document:XR
C3484381|View Sunrise:Find:Pt:Knee.right:Doc:XR
C3261715|Bladder US Ltd
C3261715|Multisection limited:Find:Pt:Urinary bladder:Doc:US
C3261715|Urinary bladder US limited
C3261715|Multisection limited:Finding:Point in time:Urinary bladder:Document:Ultrasound
C3263093|Extr a-L US
C3263093|Extremity artery - left US
C3263093|Multisection:Find:Pt:Extremity artery.left:Doc:US
C3263093|Multisection:Finding:Point in time:Extremity artery.left:Document:Ultrasound
C3263094|Renal a US
C3263094|Renal artery US
C3263094|Multisection:Finding:Point in time:Renal artery:Document:Ultrasound
C3263094|Multisection:Find:Pt:Renal artery:Doc:US
C3263105|Zygomatic arch X-ray 2 views
C3263105|Zygomatic arch XR 2V
C3263105|Views 2:Find:Pt:Zygomatic arch:Doc:XR
C3263105|Views 2:Finding:Point in time:Zygomatic arch:Document:XR
C3261473|Ankle - right X-ray Single view
C3261473|Ankle-R XR 1V
C3261473|View 1:Finding:Point in time:Ankle.right:Document:XR
C3261473|View 1:Find:Pt:Ankle.right:Doc:XR
C3262906|Abd CT Bx guid WO contr
C3262906|CT Guidance for biopsy of Abdomen-- WO contrast
C3262906|Guidance for biopsy^WO contrast:Find:Pt:Abdomen:Doc:CT
C3262906|Guidance for biopsy^WO contrast:Finding:Point in time:Abdomen:Document:Computerized Tomography
C0944158|Views:Finding:Point in time:Humerus:Narrative:XR
C0944158|Humerus X-ray
C0944158|Humerus XR
C0944158|Views:Find:Pt:Humerus:Doc:XR
C0944158|Views:Finding:Point in time:Humerus:Document:XR
C0942165|Scapula - left X-ray
C0942165|Scapula-L XR
C0942165|Views:Finding:Point in time:Scapula.left:Document:XR
C0942165|Views:Find:Pt:Scapula.left:Doc:XR
C0942193|Ankle - left MRI WO and W contrast IV
C0942193|Multisection^WO & W contrast Intravenous:Finding:Point in time:Ankle.left:Document:MRI
C0942193|Multisection^WO & W contrast IV:Find:Pt:Ankle.left:Doc:MRI
C0942193|Ankle-L MRI WO+W contr IV
C0942210|Wrist - left MRI WO and W contrast IV
C0942210|Multisection^WO & W contrast Intravenous:Finding:Point in time:Wrist.left:Document:MRI
C0942210|Multisection^WO & W contrast IV:Find:Pt:Wrist.left:Doc:MRI
C0942210|Wrist-L MRI WO+W contr IV
C0942238|Finger - left MRI
C0942238|Finger-L MRI
C0942238|Multisection:Find:Pt:Finger.left:Doc:MRI
C0942238|Multisection:Finding:Point in time:Finger.left:Document:MRI
C0942263|Should-L MRI
C0942263|Shoulder - left MRI
C0942263|Multisection:Finding:Point in time:Shoulder.left:Document:MRI
C0942263|Multisection:Find:Pt:Shoulder.left:Doc:MRI
C0947256|Scrotum+Test-R US
C0947256|Scrotum and Testicle - right US
C0947256|Multisection:Find:Pt:Scrotum+Testicle.right:Doc:US
C0947256|Multisection:Finding:Point in time:Scrotum+Testicle.right:Document:Ultrasound
C0945336|Cent v-Bl XRA LT per cath plac guid
C0945336|Fluoroscopic angiogram Guidance for placement of longterm peripheral catheter in Central vein - bilateral
C0945336|Guidance for placement of longterm peripheral catheter:Find:Pt:Central vein.bilateral:Doc:XR.fluor.angio
C0945336|Guidance for placement of longterm peripheral catheter:Finding:Point in time:Central vein.bilateral:Document:XR.fluor.angio
C0945346|Hand - left X-ray 2 views
C0945346|Hand-L XR 2V
C0945346|Views 2:Finding:Point in time:Hand.left:Document:XR
C0945346|Views 2:Find:Pt:Hand.left:Doc:XR
C0882021|Lung XR W contr IB
C0882021|Lung X-ray W contrast intrabronchial
C0882021|Views^W contrast intrabronchial:Find:Pt:Lung:Doc:XR
C0882021|Views^W contrast intrabronchial:Finding:Point in time:Lung:Document:XR
C0882104|Skull X-ray Waters
C0882104|Skull XR Waters
C0882104|View Waters:Find:Pt:Skull:Doc:XR
C0882104|View Waters:Finding:Point in time:Skull:Document:XR
C0882114|C-spine CT W contr IT
C0882114|Multisection^W contrast IT:Find:Pt:Spine.cervical:Doc:CT
C0882114|Multisection^W contrast Intrathecal:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C0882114|Cervical spine CT W contrast IT
C0882191|Wrist MRI WO+W contr IV
C0882191|Multisection^WO & W contrast Intravenous:Finding:Point in time:Wrist:Document:MRI
C0882191|Multisection^WO & W contrast IV:Find:Pt:Wrist:Doc:MRI
C0882191|Wrist MRI WO and W contrast IV
C0882219|XXX Flr Bx guid
C0882219|Fluoroscopy Guidance for biopsy of Unspecified body region
C0882219|Guidance for biopsy:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C0882219|Guidance for biopsy:Find:Pt:XXX:Doc:XR.fluor
C0942090|Vein-R XRA W contr IV
C0942090|Vein - right Fluoroscopic angiogram W contrast IV
C0942090|Views^W contrast IV:Find:Pt:Vein.right:Doc:XR.fluor.angio
C0942090|Views^W contrast Intravenous:Finding:Point in time:Vein.right:Document:XR.fluor.angio
C0942102|Carot a-R XRA W contr IA
C0942102|Carotid artery - right Fluoroscopic angiogram W contrast IA
C0942102|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.right:Document:XR.fluor.angio
C0942102|Views^W contrast IA:Find:Pt:Carotid artery.right:Doc:XR.fluor.angio
C0942127|Clavicle - right X-ray
C0942127|Clavicle-R XR
C0942127|Views:Finding:Point in time:Clavicle.right:Document:XR
C0942127|Views:Find:Pt:Clavicle.right:Doc:XR
C2607994|Hip - left X-ray
C2607994|Hip-L XR
C2607994|Views:Find:Pt:Hip.left:Doc:XR
C2607994|Views:Finding:Point in time:Hip.left:Document:XR
C0881777|Acetabulum X-ray
C0881777|Acetabulum XR
C0881777|Views:Find:Pt:Acetabulum:Doc:XR
C0881777|Views:Finding:Point in time:Acetabulum:Document:XR
C0881837|Mammogram Guidance for biopsy of Breast
C0881837|Brst Mam Bx guid
C0881837|Guidance for biopsy:Finding:Point in time:Breast:Document:Mam
C0881837|Guidance for biopsy:Find:Pt:Breast:Doc:Mam
C0881860|Chest MRI
C0881860|Multisection:Finding:Point in time:Chest:Narrative:MRI
C0881860|Multisection:Find:Pt:Chest:Doc:MRI
C0881860|Multisection:Finding:Point in time:Chest:Document:MRI
C0881869|Chest XR L-Obl port
C0881869|Chest X-ray left oblique portable
C0881869|View L-oblique portable:Find:Pt:Chest:Doc:XR
C0881869|View L-oblique portable:Finding:Point in time:Chest:Document:XR
C0881882|Chest X-ray tomograph
C0881882|Chest XRTomo
C0881882|Multisection:Find:Pt:Chest:Doc:XR.tomo
C0881882|Multisection:Finding:Point in time:Chest:Document:XR.tomo
C0881917|Face MRI WO+W contr IV
C0881917|Face MRI WO and W contrast IV
C0881917|Multisection^WO & W contrast IV:Find:Pt:Face:Doc:MRI
C0881917|Multisection^WO & W contrast Intravenous:Finding:Point in time:Face:Document:MRI
C0881970|IAC XRTomo
C0881970|Internal auditory canal X-ray tomograph
C0881970|Multisection:Finding:Point in time:Internal auditory canal:Document:XR.tomo
C0881970|Multisection:Find:Pt:Internal auditory canal:Doc:XR.tomo
C0881996|Abd XR AP+AP L-Lat Decub
C0881996|Abdomen X-ray AP and AP left lateral-decubitus
C0881996|Views AP & AP L-lateral-decubitus:Find:Pt:Abdomen:Doc:XR
C0881996|Views AP & AP L-lateral-decubitus:Finding:Point in time:Abdomen:Document:XR
C1114481|Multisection^WO & W contrast IV:Find:Pt:Internal auditory canal:Doc:MRI
C1114481|Multisection^WO & W contrast Intravenous:Finding:Point in time:Internal auditory canal:Document:MRI
C1114481|IAC MRI WO+W contr IV
C1114481|Internal auditory canal MRI WO and W contrast IV
C1114942|T-spine XR Obl 1V
C1114942|View oblique:Find:Pt:Spine.thoracic:Doc:XR
C1114942|View oblique:Finding:Point in time:Spine.thoracic:Document:XR
C1114942|Thoracic spine X-ray oblique single view
C1114642|Adrenal v XRA W contr IV
C1114642|Adrenal vein Fluoroscopic angiogram W contrast IV
C1114642|Views^W contrast IV:Find:Pt:Adrenal vein:Doc:XR.fluor.angio
C1114642|Views^W contrast Intravenous:Finding:Point in time:Adrenal vein:Document:XR.fluor.angio
C1114649|Extr lymph Flr W contr IL
C1114649|Extremity lymphatics Fluoroscopy W contrast intra lymphatic
C1114649|Views^W contrast intra lymphatic:Find:Pt:Extremity lymphatics:Doc:XR.fluor
C1114649|Views^W contrast intra lymphatic:Finding:Point in time:Extremity lymphatics:Document:XR.fluor
C1114651|Periph vv-Bl XRA W contr IV
C1114651|Peripheral veins - bilateral Fluoroscopic angiogram W contrast IV
C1114651|Views^W contrast IV:Find:Pt:Peripheral veins.bilateral:Doc:XR.fluor.angio
C1114651|Views^W contrast Intravenous:Finding:Point in time:Peripheral veins.bilateral:Document:XR.fluor.angio
C1114955|Pelvis ves MRI.Angio
C1114955|Pelvis vessels MRI angiogram
C1114955|Multisection:Finding:Point in time:Pelvis vessels:Document:MRI.angio
C1114955|Multisection:Find:Pt:Pelvis vessels:Doc:MRI.angio
C1114685|Temporomandibular joint - right X-ray
C1114685|TMJ-R XR
C1114685|Views:Finding:Point in time:Temporomandibular joint.right:Document:XR
C1114685|Views:Find:Pt:Temporomandibular joint.right:Doc:XR
C1114455|UE CT WO contr
C1114455|Upper extremity CT WO contrast
C1114455|Multisection^WO contrast:Find:Pt:Upper extremity:Doc:CT
C1114455|Multisection^WO contrast:Finding:Point in time:Upper extremity:Document:Computerized Tomography
C1114928|Fluoroscopy Guidance for placement of tube in Gastrointestine
C1114928|GI Flr Tube plac guid
C1114928|Guidance for placement of tube:Finding:Point in time:Gastrointestine:Document:XR.fluor
C1114928|Guidance for placement of tube:Find:Pt:Gastrointestine:Doc:XR.fluor
C1114465|Vein XRA Angpsty W contr IV
C1114465|Vein Fluoroscopic angiogram Angioplasty W contrast IV
C1114465|Angioplasty^W contrast Intravenous:Finding:Point in time:Vein:Document:XR.fluor.angio
C1114465|Angioplasty^W contrast IV:Find:Pt:Vein:Doc:XR.fluor.angio
C1114929|View:Finding:Point in time:To be specified in another part of the message:Narrative:XR.fluor
C1114929|XXX Flr 1V
C1114929|Unspecified body region Fluoroscopy Single view
C1114929|View 1:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1114929|View 1:Find:Pt:XXX:Doc:XR.fluor
C1114467|US Guidance for placement of catheter in Central vein-- Tunneled
C1114467|Centl v US Cath plac guid Tunneled
C1114467|Guidance for placement of catheter^tunneled:Finding:Point in time:Central vein:Document:Ultrasound
C1114467|Guidance for placement of catheter^tunneled:Find:Pt:Central vein:Doc:US
C1543472|Shoulder - right X-ray 3 views and Y
C1543472|Should-R XR 3V+Y
C1543472|Views 3 & Y:Finding:Point in time:Shoulder.right:Document:XR
C1543472|Views 3 & Y:Find:Pt:Shoulder.right:Doc:XR
C1543796|Prostate RI W Tc99mPMSA IV
C1543796|Prostate Scan W Tc-99m capromab pendatide IV
C1543796|Views^W Tc-99m capromab pendatide IV:Find:Pt:Prostate:Doc:Radnuc
C1543796|Views^W Tc-99m capromab pendatide Intravenous:Finding:Point in time:Prostate:Document:Radnuc
C1543809|Stomach Scan for gastric emptying liquid phase W radionuclide PO
C1543809|Stom RI LPGE W RNC PO
C1543809|Views for gastric emptying liquid phase^W radionuclide Oral:Finding:Point in time:Stomach:Document:Radnuc
C1543809|Views for gastric emptying liquid phase^W radionuclide PO:Find:Pt:Stomach:Doc:Radnuc
C1543812|GI SPECT W RNC IV
C1543812|Gastrointestine SPECT
C1543812|Multisection^W radionuclide IV:Find:Pt:Gastrointestine:Doc:Radnuc.SPECT
C1543812|Multisection^W radionuclide Intravenous:Finding:Point in time:Gastrointestine:Document:Radnuc.SPECT
C1542903|RI W I-131 mIBG IV
C1542903|Scan W I-131 MIBG IV
C1542903|Views^W I-131 MIBG IV:Find:Pt:^Patient:Doc:Radnuc
C1542903|Views^W I-131 MIBG Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543878|Peritoneovenous shunt Scan for patency W In-111 IT
C1543878|PV shunt RI for Pat W In-111 IT
C1543878|Views for shunt patency^W In-111 Intrathecal:Finding:Point in time:Peritoneovenous shunt:Document:Radnuc
C1543878|Views for shunt patency^W In-111 IT:Find:Pt:Peritoneovenous shunt:Doc:Radnuc
C1543893|Hrt RI FP Rest+stress+W RNC IV
C1543893|Heart Scan first pass at rest and W stress and W radionuclide IV
C1543893|Views first pass^at rest & W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543893|Views first pass^at rest & W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1542927|Hrt SPECT WM W RNC IV
C1542927|Heart SPECT wall motion
C1542927|Multisection wall motion^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1542927|Multisection wall motion^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543927|Bone SPECT Mul Areas W RNC IV
C1543927|Bone SPECT multiple areas
C1543927|Multisection multiple areas^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc.SPECT
C1543927|Multisection multiple areas^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc.SPECT
C1543951|Hrt RI Gated+WM W Stress+W RNC IV
C1543951|Heart Scan gated and wall motion W stress and W radionuclide IV
C1543951|Views gated & wall motion^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543951|Views gated & wall motion^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543953|Lung RI Clear W Tc99mDTPA AeroIH
C1543953|Lung Scan Clearance W Tc-99m DTPA aerosol IH
C1543953|Views for clearance^W Tc-99m DTPA aerosol IH:Find:Pt:Lung:Doc:Radnuc
C1543953|Views for clearance^W Tc-99m DTPA aerosol Inhalation:Finding:Point in time:Lung:Document:Radnuc
C1543954|Lung RI PF W Particulate RNC IV
C1543954|Lung Scan perfusion W particulate radionuclide IV
C1543954|Views perfusion^W particulate radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1543954|Views perfusion^W particulate radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1543955|Lung RI VP W RNC IH SB+Particulate IV
C1543955|Views ventilation & perfusion^W radionuclide IH single breath & W particulate radionuclide IV:Find:Pt:Lung:Doc:Radnuc
C1543955|Lung Scan ventilation and perfusion W radionuclide IH single breath and W particulate radionuclide IV
C1543955|Views ventilation & perfusion^W radionuclide Inhalation single breath & W particulate radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc
C1543517|Lower extremity vessels - right US.doppler limited
C1543517|LE ves-R DOP Ltd
C1543517|Multisection limited:Find:Pt:Lower extremity vessels.right:Doc:US.doppler
C1543517|Multisection limited:Finding:Point in time:Lower extremity vessels.right:Document:Ultrasound.doppler
C1543523|Upper extremity artery US.doppler
C1543523|UE a DOP
C1543523|Multisection:Finding:Point in time:Upper extremity artery:Document:Ultrasound.doppler
C1543523|Multisection:Find:Pt:Upper extremity artery:Doc:US.doppler
C1543570|Abd wall US
C1543570|Abdominal wall US
C1543570|Multisection:Finding:Point in time:Abdominal wall:Document:Ultrasound
C1543570|Multisection:Find:Pt:Abdominal wall:Doc:US
C1526353|Bone density:Tscore:Pt:Hip:Qn:XR.DXA
C1526353|Hip DXA [T-score] Bone density
C1526353|Hip DXA T-score BDM
C1526353|Bone density:T Score:Point in time:Hip:Quantitative:XR.DXA
C1543590|Wrist-R XR Lat W FE
C1543590|Wrist - right X-ray lateral W flexion and W extension
C1543590|Views lateral^W flexion & W extension:Finding:Point in time:Wrist.right:Document:XR
C1543590|Views lateral^W flexion & W extension:Find:Pt:Wrist.right:Doc:XR
C1542860|GI+Resp Sys XR for FB
C1542860|Gastrointestinal system and Respiratory system X-ray for foreign body
C1542860|View for foreign body:Find:Pt:Gastrointestinal system+Respiratory system:Doc:XR
C1542860|View for foreign body:Finding:Point in time:Gastrointestinal system+Respiratory system:Document:XR
C1526764|Wrist-R XR Ulnar+Radial Deviation
C1526764|Wrist - right X-ray ulnar deviation and radial deviation
C1526764|Views ulnar deviation & radial deviation:Finding:Point in time:Wrist.right:Document:XR
C1526764|Views ulnar deviation & radial deviation:Find:Pt:Wrist.right:Doc:XR
C1543716|Hrt SPECT for Infarct W Tc99mPyp IV
C1543716|Heart SPECT for infarct W Tc-99m PYP IV
C1543716|Multisection for infarct^W Tc-99m PYP IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543716|Multisection for infarct^W Tc-99m PYP Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1524427|Knee-Bl CT
C1524427|Knee - bilateral CT
C1524427|Multisection:Finding:Point in time:Knee.bilateral:Document:Computerized Tomography
C1524427|Multisection:Find:Pt:Knee.bilateral:Doc:CT
C1524176|Scapula MRI
C1524176|Multisection:Finding:Point in time:Scapula:Document:MRI
C1524176|Multisection:Find:Pt:Scapula:Doc:MRI
C1524824|Breast - right MRI WO contrast
C1524824|Brst-R MRI WO contr
C1524824|Multisection^WO contrast:Find:Pt:Breast.right:Doc:MRI
C1524824|Multisection^WO contrast:Finding:Point in time:Breast.right:Document:MRI
C1524844|UE-R MRI WO contr
C1524844|Upper extremity - right MRI WO contrast
C1524844|Multisection^WO contrast:Find:Pt:Upper extremity.right:Doc:MRI
C1524844|Multisection^WO contrast:Finding:Point in time:Upper extremity.right:Document:MRI
C1525109|Veins MRI angiogram
C1525109|Veins MRI.Angio
C1525109|Multisection:Finding:Point in time:Veins:Document:MRI.angio
C1525109|Multisection:Find:Pt:Veins:Doc:MRI.angio
C1524236|Lower extremity joint - left MRI limited WO contrast
C1524236|LE.joint-L MRI Ltd WO contr
C1524236|Multisection limited^WO contrast:Find:Pt:Lower extremity.joint.left:Doc:MRI
C1524236|Multisection limited^WO contrast:Finding:Point in time:Lower extremity.joint.left:Document:MRI
C1525303|Wrist-L XR Lat W Ext
C1525303|Wrist - left X-ray lateral W extension
C1525303|View lateral^W extension:Find:Pt:Wrist.left:Doc:XR
C1525303|View lateral^W extension:Finding:Point in time:Wrist.left:Document:XR
C1525322|L-spine XR Lat Xtable
C1525322|View lateral crosstable:Find:Pt:Spine.lumbar:Doc:XR
C1525322|View lateral crosstable:Finding:Point in time:Spine.lumbar:Document:XR
C1525322|Lumbar spine X-ray lateral crosstable
C1525249|Head veins MRI angiogram WO contrast
C1525249|Head vv MRI.Angio WO contr
C1525249|Multisection^WO contrast:Find:Pt:Head veins:Doc:MRI.angio
C1525249|Multisection^WO contrast:Finding:Point in time:Head veins:Document:MRI.angio
C1525333|Foot X-ray lateral standing
C1525333|Ft XR Lat stand
C1525333|View lateral^standing:Find:Pt:Foot:Doc:XR
C1525333|View lateral^standing:Finding:Point in time:Foot:Document:XR
C1525338|Breast - bilateral Mammogram MLO
C1525338|Brst-Bl Mam MLO
C1525338|View MLO:Finding:Point in time:Breast.bilateral:Document:Mam
C1525338|View MLO:Find:Pt:Breast.bilateral:Doc:Mam
C1524685|Breast - left Mammogram roll
C1524685|Brst-L Mam Roll
C1524685|Views roll:Finding:Point in time:Breast.left:Document:Mam
C1524685|Views roll:Find:Pt:Breast.left:Doc:Mam
C1525457|Breast - left Mammogram tangential
C1525457|Brst-L Mam Tangential
C1525457|View tangential:Finding:Point in time:Breast.left:Document:Mam
C1525457|View tangential:Find:Pt:Breast.left:Doc:Mam
C1524229|Scapula-L XR Y
C1524229|Scapula - left X-ray Y
C1524229|View Y:Find:Pt:Scapula.left:Doc:XR
C1524229|View Y:Finding:Point in time:Scapula.left:Document:XR
C1524245|Ankle-L XR AP+Lat+Mortise
C1524245|Ankle - left X-ray AP and lateral and Mortise
C1524245|Views AP & lateral & Mortise:Finding:Point in time:Ankle.left:Document:XR
C1524245|Views AP & lateral & Mortise:Find:Pt:Ankle.left:Doc:XR
C1524252|C-spine XR AP+Odont+Lat W FE
C1524252|Views AP & odontoid & lateral^W flexion & W extension:Find:Pt:Spine.cervical:Doc:XR
C1524252|Views AP & odontoid & lateral^W flexion & W extension:Finding:Point in time:Spine.cervical:Document:XR
C1524252|Cervical spine X-ray AP and odontoid and lateral W flexion and W extension
C1525606|CT Guidance for aspiration of cyst of Abdomen
C1525606|Abd CT Cyst Asp guid
C1525606|Guidance for aspiration of cyst:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1525606|Guidance for aspiration of cyst:Find:Pt:Abdomen:Doc:CT
C1527068|Parotid gland CT
C1527068|Multisection:Find:Pt:Parotid gland:Doc:CT
C1527068|Multisection:Finding:Point in time:Parotid gland:Document:Computerized Tomography
C1525628|Mediastinum XRTomo
C1525628|Mediastinum X-ray tomograph
C1525628|Multisection:Find:Pt:Mediastinum:Doc:XR.tomo
C1525628|Multisection:Finding:Point in time:Mediastinum:Document:XR.tomo
C1525634|Parotid gland CT W contr IV
C1525634|Parotid gland CT W contrast IV
C1525634|Multisection^W contrast Intravenous:Finding:Point in time:Parotid gland:Document:Computerized Tomography
C1525634|Multisection^W contrast IV:Find:Pt:Parotid gland:Doc:CT
C1525642|TMJ-R CT W contr IV
C1525642|Temporomandibular joint - right CT W contrast IV
C1525642|Multisection^W contrast IV:Find:Pt:Temporomandibular joint.right:Doc:CT
C1525642|Multisection^W contrast Intravenous:Finding:Point in time:Temporomandibular joint.right:Document:Computerized Tomography
C1525643|TMJ-R MRI W contr IV
C1525643|Temporomandibular joint - right MRI W contrast IV
C1525643|Multisection^W contrast IV:Find:Pt:Temporomandibular joint.right:Doc:MRI
C1525643|Multisection^W contrast Intravenous:Finding:Point in time:Temporomandibular joint.right:Document:MRI
C1525675|Sternoclavicular joint - bilateral X-ray Serendipity
C1525675|SC joint-Bl XR Serendipity
C1525675|View Serendipity:Find:Pt:Sternoclavicular joint.bilateral:Doc:XR
C1525675|View Serendipity:Finding:Point in time:Sternoclavicular joint.bilateral:Document:XR
C1525677|LS-spine junc XR True AP
C1525677|Spine Lumbosacral Junction X-ray true AP
C1525677|View true AP:Finding:Point in time:Spine.lumbosacral junction:Document:XR
C1525677|View true AP:Find:Pt:Spine.lumbosacral junction:Doc:XR
C1525683|Humerus bicipital groove - bilateral X-ray
C1525683|Humerus bicipital groove-Bl XR
C1525683|Views:Find:Pt:Humerus.bicipital groove.bilateral:Doc:XR
C1525683|Views:Finding:Point in time:Humerus.bicipital groove.bilateral:Document:XR
C1525720|Celiac a+SMA+IMA XRA W contr IA
C1525720|Celiac artery and Superior mesenteric artery and Inferior mesenteric artery Fluoroscopic angiogram W contrast IA
C1525720|Views^W contrast Intra-arterial:Finding:Point in time:Celiac artery+Superior mesenteric artery+Inferior mesenteric artery:Document:XR.fluor.angio
C1525720|Views^W contrast IA:Find:Pt:Celiac artery+Superior mesenteric artery+Inferior mesenteric artery:Doc:XR.fluor.angio
C1525741|Intraosseous vv XRA W contr IV
C1525741|Intraosseous veins Fluoroscopic angiogram W contrast IV
C1525741|Views^W contrast IV:Find:Pt:Intraosseous veins:Doc:XR.fluor.angio
C1525741|Views^W contrast Intravenous:Finding:Point in time:Intraosseous veins:Document:XR.fluor.angio
C1525742|Jugular v-L XRA W contr IV
C1525742|Jugular vein - left Fluoroscopic angiogram W contrast IV
C1525742|Views^W contrast Intravenous:Finding:Point in time:Jugular vein.left:Document:XR.fluor.angio
C1525742|Views^W contrast IV:Find:Pt:Jugular vein.left:Doc:XR.fluor.angio
C1524691|Wrist - left MRI W contrast IS
C1524691|Multisection^W contrast Intrasynovial:Finding:Point in time:Wrist.left:Document:MRI
C1524691|Wrist-L MRI W contr IS
C1524691|Multisection^W contrast IS:Find:Pt:Wrist.left:Doc:MRI
C1525878|Acromioclavicular Joint X-ray WO weight
C1525878|AC joint XR WO Wt
C1525878|Views^WO weight:Finding:Point in time:Acromioclavicular joint:Document:XR
C1525878|Views^WO weight:Find:Pt:Acromioclavicular joint:Doc:XR
C1525994|Wrist - right X-ray 2 views tunnel.carpal
C1525994|Wrist-R XR 2V Tunnel
C1525994|Views 2 tunnel.carpal:Find:Pt:Wrist.right:Doc:XR
C1525994|Views 2 tunnel.carpal:Finding:Point in time:Wrist.right:Document:XR
C1526003|Views oblique:Finding:Point in time:Elbow.right:Narrative:XR
C1526003|Elbow-R XR Obl
C1526003|Elbow - right X-ray oblique
C1526003|Views oblique:Find:Pt:Elbow.right:Doc:XR
C1526003|Views oblique:Finding:Point in time:Elbow.right:Document:XR
C1526124|Temporomandibular joint - right X-ray tomograph
C1526124|TMJ-R XRTomo
C1526124|Multisection:Find:Pt:Temporomandibular joint.right:Doc:XR.tomo
C1526124|Multisection:Finding:Point in time:Temporomandibular joint.right:Document:XR.tomo
C1526046|Hip-R XR Lat
C1526046|Hip - right X-ray lateral
C1526046|View lateral:Find:Pt:Hip.right:Doc:XR
C1526046|View lateral:Finding:Point in time:Hip.right:Document:XR
C1526065|Knee-R XR AP+Lat+Sunrise
C1526065|Knee - right X-ray AP and lateral and Sunrise
C1526065|Views AP & lateral & Sunrise:Find:Pt:Knee.right:Doc:XR
C1526065|Views AP & lateral & Sunrise:Finding:Point in time:Knee.right:Document:XR
C1525121|Brst-R Mam True Lat
C1525121|Breast - right Mammogram true lateral
C1525121|View true lateral:Finding:Point in time:Breast.right:Document:Mam
C1525121|View true lateral:Find:Pt:Breast.right:Doc:Mam
C1526156|Sinuses XR Lat+Caldwell+Waters
C1526156|Sinuses X-ray lateral and Caldwell and Waters
C1526156|Views lateral & Caldwell & Waters:Finding:Point in time:Sinuses:Document:XR
C1526156|Views lateral & Caldwell & Waters:Find:Pt:Sinuses:Doc:XR
C1526310|Bladder Flr W Chain+contr IB
C1526310|Urinary bladder Fluoroscopy W chain and contrast intra bladder
C1526310|Views^W chain & contrast intra bladder:Find:Pt:Urinary bladder:Doc:XR.fluor
C1526310|Views^W chain & contrast intra bladder:Finding:Point in time:Urinary bladder:Document:XR.fluor
C1526328|Tib+Fib-R XR 2V Obl
C1526328|Tibia - right and Fibula - right X-ray 2 views Oblique
C1526328|Views 2 oblique:Finding:Point in time:Tibia.right+Fibula.right:Document:XR
C1526328|Views 2 oblique:Find:Pt:Tibia.right+Fibula.right:Doc:XR
C1524469|Knee MRI W contrast IS
C1524469|Multisection^W contrast Intrasynovial:Finding:Point in time:Knee:Document:MRI
C1524469|Multisection^W contrast IS:Find:Pt:Knee:Doc:MRI
C1524469|Knee MRI W contr IS
C1524872|Hip - left CT WO contrast
C1524872|Hip-L CT WO contr
C1524872|Multisection^WO contrast:Finding:Point in time:Hip.left:Document:Computerized Tomography
C1524872|Multisection^WO contrast:Find:Pt:Hip.left:Doc:CT
C1524522|Ft CT W contr IV
C1524522|Foot CT W contrast IV
C1524522|Multisection^W contrast IV:Find:Pt:Foot:Doc:CT
C1524522|Multisection^W contrast Intravenous:Finding:Point in time:Foot:Document:Computerized Tomography
C1524533|Forearm-R CT W contr IV
C1524533|Forearm - right CT W contrast IV
C1524533|Multisection^W contrast Intravenous:Finding:Point in time:Forearm.right:Document:Computerized Tomography
C1524533|Multisection^W contrast IV:Find:Pt:Forearm.right:Doc:CT
C1524540|Hand-R MRI W contr IV
C1524540|Hand - right MRI W contrast IV
C1524540|Multisection^W contrast IV:Find:Pt:Hand.right:Doc:MRI
C1524540|Multisection^W contrast Intravenous:Finding:Point in time:Hand.right:Document:MRI
C1524171|Hip-R CT W contr IV
C1524171|Hip - right CT W contrast IV
C1524171|Multisection^W contrast IV:Find:Pt:Hip.right:Doc:CT
C1524171|Multisection^W contrast Intravenous:Finding:Point in time:Hip.right:Document:Computerized Tomography
C1524906|Spine CT WO contrast
C1524906|Spine CT WO contr
C1524906|Multisection^WO contrast:Find:Pt:Spine:Doc:CT
C1524906|Multisection^WO contrast:Finding:Point in time:Spine:Document:Computerized Tomography
C1524918|Uterus MRI WO contr
C1524918|Uterus MRI WO contrast
C1524918|Multisection^WO contrast:Find:Pt:Uterus:Doc:MRI
C1524918|Multisection^WO contrast:Finding:Point in time:Uterus:Document:MRI
C1524586|Should-L CT W contr IV
C1524586|Shoulder - left CT W contrast IV
C1524586|Multisection^W contrast IV:Find:Pt:Shoulder.left:Doc:CT
C1524586|Multisection^W contrast Intravenous:Finding:Point in time:Shoulder.left:Document:Computerized Tomography
C1524199|Shoulder - left X-ray Single view
C1524199|Should-L XR 1V
C1524199|View 1:Find:Pt:Shoulder.left:Doc:XR
C1524199|View 1:Finding:Point in time:Shoulder.left:Document:XR
C1524308|Chest CT Bx guid W contr IV
C1524308|CT Guidance for biopsy of Chest-- W contrast IV
C1524308|Guidance for biopsy^W contrast IV:Find:Pt:Chest:Doc:CT
C1524308|Guidance for biopsy^W contrast Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C1524130|Multisection^WO & W contrast IV:Find:Pt:Internal auditory canal:Doc:CT
C1524130|IAC CT WO+W contr IV
C1524130|Internal auditory canal CT WO and W contrast IV
C1524130|Multisection^WO & W contrast Intravenous:Finding:Point in time:Internal auditory canal:Document:Computerized Tomography
C1524329|CT Guidance for nerve block of Abdomen
C1524329|Abd CT Nerve Block guid
C1524329|Guidance for nerve block:Find:Pt:Abdomen:Doc:CT
C1524329|Guidance for nerve block:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524340|Ankle-L CT
C1524340|Ankle - left CT
C1524340|Multisection:Finding:Point in time:Ankle.left:Document:Computerized Tomography
C1524340|Multisection:Find:Pt:Ankle.left:Doc:CT
C1524641|Thumb-L XR 3V
C1524641|Thumb - left X-ray 3 views
C1524641|Views 3:Finding:Point in time:Thumb.left:Document:XR
C1524641|Views 3:Find:Pt:Thumb.left:Doc:XR
C1524997|Elbow - bilateral X-ray 2 views
C1524997|Elbow-Bl XR 2V
C1524997|Views 2:Find:Pt:Elbow.bilateral:Doc:XR
C1524997|Views 2:Finding:Point in time:Elbow.bilateral:Document:XR
C1524729|Multisection^WO & W contrast Intravenous:Finding:Point in time:Foot.left:Document:Computerized Tomography
C1524729|Foot - left CT WO and W contrast IV
C1524729|Multisection^WO & W contrast IV:Find:Pt:Foot.left:Doc:CT
C1524729|Ft-L CT WO+W contr IV
C1524737|Multisection^WO & W contrast Intravenous:Finding:Point in time:Forearm.right:Document:MRI
C1524737|Multisection^WO & W contrast IV:Find:Pt:Forearm.right:Doc:MRI
C1524737|Forearm - right MRI WO and W contrast IV
C1524737|Forearm-R MRI WO+W contr IV
C1524739|Multisection^WO & W contrast IV:Find:Pt:Hand.left:Doc:CT
C1524739|Hand - left CT WO and W contrast IV
C1524739|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hand.left:Document:Computerized Tomography
C1524739|Hand-L CT WO+W contr IV
C1524760|Multisection^WO & W contrast IV:Find:Pt:Upper extremity.joint:Doc:MRI
C1524760|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity.joint:Document:MRI
C1524760|UE joint MRI WO+W contr IV
C1524760|Upper extremity.joint MRI WO and W contrast IV
C1525034|Femur-L XR AP+Lat
C1525034|Femur - left X-ray AP and lateral
C1525034|Views AP & lateral:Find:Pt:Femur.left:Doc:XR
C1525034|Views AP & lateral:Finding:Point in time:Femur.left:Document:XR
C1525046|Humerus-Bl XR AP+Lat
C1525046|Humerus - bilateral X-ray AP and lateral
C1525046|Views AP & lateral:Finding:Point in time:Humerus.bilateral:Document:XR
C1525046|Views AP & lateral:Find:Pt:Humerus.bilateral:Doc:XR
C1527047|Hip MRI
C1527047|Multisection:Finding:Point in time:Hip:Narrative:MRI
C1527047|Multisection:Find:Pt:Hip:Doc:MRI
C1527047|Multisection:Finding:Point in time:Hip:Document:MRI
C1524778|Multisection^WO & W contrast Intravenous:Finding:Point in time:Scapula.left:Document:MRI
C1524778|Scapula-L MRI WO+W contr IV
C1524778|Multisection^WO & W contrast IV:Find:Pt:Scapula.left:Doc:MRI
C1524778|Scapula - left MRI WO and W contrast IV
C1524788|Multisection^WO & W contrast IV:Find:Pt:Spine.thoracic:Doc:CT
C1524788|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C1524788|T-spine CT WO+W contr IV
C1524788|Thoracic spine CT WO and W contrast IV
C1830193|XXX CT Drain guid W contr IV
C1830193|CT Guidance for drainage of Unspecified body region-- W contrast IV
C1830193|Guidance for drainage^W contrast IV:Find:Pt:XXX:Doc:CT
C1830193|Guidance for drainage^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1830209|LE.L vels CT.Angio WO+W contr IV
C1830209|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.left>Vessels:Document:Computerized Tomography.angio
C1830209|Lower extremity - left Vessels CT angiogram WO and W contrast IV
C1830209|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.left>Vessels:Doc:CT.angio
C1830241|Spine Lumbosacral Junction X-ray
C1830241|LS-spine junc XR
C1830241|Views:Find:Pt:Spine.lumbosacral junction:Doc:XR
C1830241|Views:Finding:Point in time:Spine.lumbosacral junction:Document:XR
C1830245|Elbow - left X-ray GE 3 views
C1830245|Elbow-L XR GE 3V
C1830245|Views GE 3:Finding:Point in time:Elbow.left:Document:XR
C1830245|Views GE 3:Find:Pt:Elbow.left:Doc:XR
C1830254|Deprecated Chest XR PA+Lat+Obl
C1830254|Deprecated Chest X-ray PA & lateral & oblique
C1830254|Views PA & lateral & oblique:Find:Pt:Chest:Nar:XR
C1830254|Views PA & lateral & oblique:Finding:Point in time:Chest:Narrative:XR
C1715416|Brain RI Flow W Tc99mBicisate IV
C1715416|Brain Scan flow W Tc-99m bicisate IV
C1715416|Views flow^W Tc-99m bicisate Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1715416|Views flow^W Tc-99m bicisate IV:Find:Pt:Brain:Doc:Radnuc
C1715436|Chest Pleura US Bx needle guid
C1715436|US Guidance for needle biopsy of Chest Pleura
C1715436|Guidance for biopsy.needle:Finding:Point in time:Chest>Pleura:Document:Ultrasound
C1715436|Guidance for biopsy.needle:Find:Pt:Chest>Pleura:Doc:US
C1715437|US Guidance for drainage of Pancreas
C1715437|Pancreas US Drain guid
C1715437|Guidance for drainage:Find:Pt:Pancreas:Doc:US
C1715437|Guidance for drainage:Finding:Point in time:Pancreas:Document:Ultrasound
C1715484|XXX Flr Tube plac guid
C1715484|Fluoroscopy Guidance for placement of tube in Unspecified body region
C1715484|Guidance for placement of tube:Find:Pt:XXX:Doc:XR.fluor
C1715484|Guidance for placement of tube:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1714915|Thigh ves-L MRI.Angio WO contr
C1714915|Thigh vessels - left MRI angiogram WO contrast
C1714915|Multisection^WO contrast:Finding:Point in time:Thigh vessels.left:Document:MRI.angio
C1714915|Multisection^WO contrast:Find:Pt:Thigh vessels.left:Doc:MRI.angio
C1714933|Views 4:Finding:Point in time:Mandible.right:Document:XR
C1714933|Deprecated Mandible-R XR 4V
C1714933|Deprecated Mandible - right X-ray 4 views
C1714933|Views 4:Find:Pt:Mandible.right:Doc:XR
C1714935|C-spine XRVideo
C1714935|Views:Find:Pt:Spine.cervical:Doc:XR.fluor.video
C1714935|Views:Finding:Point in time:Spine.cervical:Document:XR.fluor.video
C1714935|Cervical spine Fluoroscopy video
C1706621|Deprecated Finger.5th-R XR GE 3V
C1706621|Views GE 3:Find:Pt:Finger.fifth.right:Nar:XR
C1706621|Deprecated Finger fifth Right X-ray GE 3 views
C1706621|Views GE 3:Finding:Point in time:Finger.fifth.right:Narrative:XR
C1714955|Bone CT
C1714955|Guidance for deep biopsy.needle:Finding:Point in time:Bone:Document:Computerized Tomography
C1714955|CT Guidance for deep biopsy.needle of Bone
C1714955|Guidance for deep biopsy.needle:Find:Pt:Bone:Doc:CT
C1717221|Brst-L US Localization guid
C1717221|US Guidance for localization of Breast - left
C1717221|Guidance for localization:Find:Pt:Breast.left:Doc:US
C1717221|Guidance for localization:Finding:Point in time:Breast.left:Document:Ultrasound
C1715101|Kidney - bilateral US
C1715101|Multisection:Find:Pt:Kidney.bilateral:Doc:US
C1715101|Multisection:Finding:Point in time:Kidney.bilateral:Document:Ultrasound
C1715101|Kdny-Bl US
C1715109|Renal v XRA W contr IV+Renin Samp
C1715109|Renal vein Fluoroscopic angiogram W contrast IV and W renin sampling
C1715109|Views^W contrast Intravenous & W renin sampling:Finding:Point in time:Renal vein:Document:XR.fluor.angio
C1715109|Views^W contrast IV & W renin sampling:Find:Pt:Renal vein:Doc:XR.fluor.angio
C1636059|L-spine XR AP W+WO R+L-bending
C1636059|Views AP^W R-bending & W L-bending & WO bending:Find:Pt:Spine.lumbar:Doc:XR
C1636059|Views AP^W R-bending & W L-bending & WO bending:Finding:Point in time:Spine.lumbar:Document:XR
C1636059|Lumbar spine X-ray AP W right bending and W left bending and WO bending
C1636062|Chest XR R-Obl+L-Obl W nipple markers
C1636062|Chest X-ray right oblique and left oblique W nipple markers
C1636062|Views R-oblique & L-oblique^W nipple markers:Find:Pt:Chest:Doc:XR
C1636062|Views R-oblique & L-oblique^W nipple markers:Finding:Point in time:Chest:Document:XR
C1636070|US Guidance for aspiration of cyst of Thyroid
C1636070|Thyroid US Cyst Asp guid
C1636070|Guidance for aspiration of cyst:Finding:Point in time:Thyroid:Document:Ultrasound
C1636070|Guidance for aspiration of cyst:Find:Pt:Thyroid:Doc:US
C1636078|Surgical specimen US
C1636078|Surg Spec US
C1636078|Multisection:Find:Pt:Surgical specimen:Doc:US
C1636078|Multisection:Finding:Point in time:Surgical specimen:Document:Ultrasound
C1643245|Ankle - right X-ray portable
C1643245|Ankle-R XR port
C1643245|Views portable:Find:Pt:Ankle.right:Doc:XR
C1643245|Views portable:Finding:Point in time:Ankle.right:Document:XR
C1631785|Extremity CT WO contrast
C1631785|Extr CT WO contr
C1631785|Multisection^WO contrast:Find:Pt:Extremity:Doc:CT
C1631785|Multisection^WO contrast:Finding:Point in time:Extremity:Document:Computerized Tomography
C1978441|Portal+Hepatic v XRA TIPS plac guid
C1978441|Fluoroscopic angiogram Guidance for placement of transjugular intrahepatic portosystemic shunt in Portal vein and Hepatic vein
C1978441|Guidance for placement of transjugular intrahepatic portosystemic shunt:Find:Pt:Portal vein+Hepatic vein:Doc:XR.fluor.angio
C1978441|Guidance for placement of transjugular intrahepatic portosystemic shunt:Finding:Point in time:Portal vein+Hepatic vein:Document:XR.fluor.angio
C1977321|Thoracic Spine vessels MRI angiogram
C1977321|T-spine ves MRI.Angio
C1977321|Multisection:Finding:Point in time:Spine.thoracic vessels:Document:MRI.angio
C1977321|Multisection:Find:Pt:Spine.thoracic vessels:Doc:MRI.angio
C1953948|Spine CT WO+W contr IT
C1953948|Spine CT WO and W contrast IT
C1953948|Multisection^WO & W contrast IT:Find:Pt:Spine:Doc:CT
C1953948|Multisection^WO & W contrast Intrathecal:Finding:Point in time:Spine:Document:Computerized Tomography
C1953957|Orbit CT WO and W contrast IV
C1953957|Orbit CT WO+W contr IV
C1953957|Multisection^WO & W contrast IV:Find:Pt:Head>Orbit:Doc:CT
C1953957|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head>Orbit:Document:Computerized Tomography
C1953981|L-spine+Sacrum XR 4V
C1953981|Spine Lumbar and Sacrum X-ray 4 views
C1953981|Views 4:Finding:Point in time:Spine.lumbar+Sacrum:Document:XR
C1953981|Views 4:Find:Pt:Spine.lumbar+Sacrum:Doc:XR
C1953988|Ankle-Bl XR GE 3V
C1953988|Ankle - bilateral X-ray GE 3 views
C1953988|Views GE 3:Find:Pt:Ankle.bilateral:Doc:XR
C1953988|Views GE 3:Finding:Point in time:Ankle.bilateral:Document:XR
C2734944|Esoph PET
C2734944|Esophagus PET
C2734944|Multisection:Find:Pt:Esophagus:Doc:Radnuc.PET
C2734944|Multisection:Finding:Point in time:Esophagus:Document:Radnuc.PET
C3174148|US Guidance for placement of needle in Unspecified body region
C3174148|XXX US Needle plac guid
C3174148|Guidance for placement of needle:Find:Pt:XXX:Doc:US
C3174148|Guidance for placement of needle:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C3174369|SS v+Jugular v-L XRA W contr IV
C3174369|Sagittal sinus and Jugular veins - left Fluoroscopic angiogram W contrast IV
C3174369|Views^W contrast Intravenous:Finding:Point in time:Sagittal sinus vein.left+Jugular vein.left:Document:XR.fluor.angio
C3174369|Views^W contrast IV:Find:Pt:Sagittal sinus vein.left+Jugular vein.left:Doc:XR.fluor.angio
C3533573|Multisection:Find:Pt:Axilla.left:Doc:US
C3533573|Axilla-L US
C3533573|Axilla - left US
C3533573|Multisection:Finding:Point in time:Axilla.left:Document:Ultrasound
C3533549|Guidance for kyphoplasty:Find:Pt:Spine.thoracic:Doc:XR.fluor
C3533549|T-spine Flr Kyphoplasty guid
C3533549|Guidance for kyphoplasty:Finding:Point in time:Spine.thoracic:Document:XR.fluor
C3533549|Fluoroscopy Guidance for kyphoplasty of Thoracic spine
C3533903|Brst-Bl FFDM-DBT Screening
C3533903|Breast - bilateral FFD mammogram-tomosynthesis screening
C3533903|Multisection screening:Find:Pt:Breast.bilateral:Doc:Mam.FFD.tomosynthesis
C3533903|Multisection screening:Finding:Point in time:Breast.bilateral:Document:Mam.FFD.tomosynthesis
C3533794|Multisection^WO & W contrast IV:Find:Pt:Chest+Abdomen+Pelvis:Doc:CT
C3533794|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest+Abdomen+Pelvis:Document:Computerized Tomography
C3533794|Chest+Abd+Pelvis CT WO+W contr IV
C3533794|Chest and Abdomen and Pelvis CT WO and W contrast IV
C3533792|Chest+Abd+Pelvis CT W contr IV
C3533792|Multisection^W contrast IV:Find:Pt:Chest+Abdomen+Pelvis:Doc:CT
C3533792|Multisection^W contrast Intravenous:Finding:Point in time:Chest+Abdomen+Pelvis:Document:Computerized Tomography
C3533792|Chest and Abdomen and Pelvis CT W contrast IV
C3262931|Multisection^WO & W contrast:Finding:Point in time:Pulmonary vessels:Document:Computerized Tomography.angio
C3262931|Deprecated Pulmonary vessels CT angiogram WO and W contrast
C3262931|Multisection^WO & W contrast:Find:Pt:Pulmonary vessels:Doc:CT.angio
C3262931|Deprecated Pulm ves CT.Angio WO+W contr
C3262968|Knee - left X-ray Sunrise and (views standing)
C3262968|Knee-L XR Sunrise+(views Stand)
C3262968|View Sunrise & (views^standing):Find:Pt:Knee.left:Doc:XR
C3262968|View Sunrise & (views^standing):Finding:Point in time:Knee.left:Document:XR
C3262972|Shoulder - left X-ray AP and Grashey and axillary
C3262972|Should-L XR AP+Grashey+Ax
C3262972|Views AP & Grashey & axillary:Finding:Point in time:Shoulder.left:Document:XR
C3262972|Views AP & Grashey & axillary:Find:Pt:Shoulder.left:Doc:XR
C3482448|T-spine Flr W contr ID
C3482448|Views^W contrast intradisc:Find:Pt:Spine.thoracic:Doc:XR.fluor
C3482448|Views^W contrast intradisc:Finding:Point in time:Spine.thoracic:Document:XR.fluor
C3482448|Thoracic spine Fluoroscopy W contrast intradisc
C3263019|MRI Guidance for needle biopsy of Pancreas
C3263019|Pancreas MRI Bx needle guid
C3263019|Guidance for biopsy.needle:Find:Pt:Pancreas:Doc:MRI
C3263019|Guidance for biopsy.needle:Finding:Point in time:Pancreas:Document:MRI
C3262467|Salivary gland MRI Bx needle guid
C3262467|MRI Guidance for needle biopsy of Salivary gland
C3262467|Guidance for biopsy.needle:Find:Pt:Salivary gland:Doc:MRI
C3262467|Guidance for biopsy.needle:Finding:Point in time:Salivary gland:Document:MRI
C3263042|Liver SPECT W Tc99mSC IV
C3263042|Liver SPECT W Tc-99m SC IV
C3263042|Multisection^W Tc-99m Subcutaneous Intravenous:Finding:Point in time:Liver:Document:Radnuc.SPECT
C3263042|Multisection^W Tc-99m SC IV:Find:Pt:Liver:Doc:Radnuc.SPECT
C3263051|Urinary Bladder and Urethra SPECT W contrast intra bladder during voiding
C3263051|Bladder+Urethra SPECT W contr IB void
C3263051|Multisection^W contrast intra bladder during voiding:Find:Pt:Urinary bladder+Urethra:Doc:Radnuc.SPECT
C3263051|Multisection^W contrast intra bladder during voiding:Finding:Point in time:Urinary bladder+Urethra:Document:Radnuc.SPECT
C3263065|Pulmonary artery Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C3263065|PA XRA PTA of ves W contr IA
C3263065|Percutaneous transluminal angioplasty of vessel^W contrast Intra-arterial:Finding:Point in time:Pulmonary artery:Document:XR.fluor.angio
C3263065|Percutaneous transluminal angioplasty of vessel^W contrast IA:Find:Pt:Pulmonary artery:Doc:XR.fluor.angio
C3263099|Scrotum and Testicle US limited
C3263099|Scrotum+Test US Ltd
C3263099|Multisection limited:Find:Pt:Scrotum+Testicle:Doc:US
C3263099|Multisection limited:Finding:Point in time:Scrotum+Testicle:Document:Ultrasound
C3263107|Ankle-L XR 1V
C3263107|Ankle - left X-ray Single view
C3263107|View 1:Find:Pt:Ankle.left:Doc:XR
C3263107|View 1:Finding:Point in time:Ankle.left:Document:XR
C3262900|Brachiocephalic artery Fluoroscopic angiogram W contrast IA
C3262900|BrachCeph a XRA W contr IA
C3262900|Views^W contrast Intra-arterial:Finding:Point in time:Brachiocephalic artery:Document:XR.fluor.angio
C3262900|Views^W contrast IA:Find:Pt:Brachiocephalic artery:Doc:XR.fluor.angio
C3262921|Muscle CT Bx needle guid
C3262921|CT Guidance for needle biopsy of Muscle
C3262921|Guidance for biopsy.needle:Find:Pt:Muscle:Doc:CT
C3262921|Guidance for biopsy.needle:Finding:Point in time:Muscle:Document:Computerized Tomography
C3262924|Thyroid CT Bx needle guid
C3262924|CT Guidance for needle biopsy of Thyroid
C3262924|Guidance for biopsy.needle:Finding:Point in time:Thyroid:Document:Computerized Tomography
C3262924|Guidance for biopsy.needle:Find:Pt:Thyroid:Doc:CT
C2607996|Views:Finding:Point in time:Spine:Narrative:XR
C2607996|Spine X-ray
C2607996|Spine XR
C2607996|Views:Find:Pt:Spine:Doc:XR
C2607996|Views:Finding:Point in time:Spine:Document:XR
C0942170|Thumb - bilateral X-ray
C0942170|Thumb-Bl XR
C0942170|Views:Finding:Point in time:Thumb.bilateral:Document:XR
C0942170|Views:Find:Pt:Thumb.bilateral:Doc:XR
C0942225|Extremity - bilateral US
C0942225|Extr-Bl US
C0942225|Multisection:Find:Pt:Extremity.bilateral:Doc:US
C0942225|Multisection:Finding:Point in time:Extremity.bilateral:Document:Ultrasound
C0945325|Upper extremity - bilateral MRI
C0945325|UE-Bl MRI
C0945325|Multisection:Find:Pt:Upper extremity.bilateral:Doc:MRI
C0945325|Multisection:Finding:Point in time:Upper extremity.bilateral:Document:MRI
C0942257|Popliteal space-Bl US
C0942257|Popliteal space - bilateral US
C0942257|Multisection:Find:Pt:Popliteal space.bilateral:Doc:US
C0942257|Multisection:Finding:Point in time:Popliteal space.bilateral:Document:Ultrasound
C0942266|Scrotum+Test-Bl US
C0942266|Scrotum and Testicle - bilateral US
C0942266|Multisection:Finding:Point in time:Scrotum+Testicle.bilateral:Document:Ultrasound
C0942266|Multisection:Find:Pt:Scrotum+Testicle.bilateral:Doc:US
C0942286|Brst-R Mam Bx Str Guid
C0942286|Guidance for stereotactic biopsy:Find:Pt:Breast.right:Doc:Mam
C0942286|Mammogram Guidance for stereotactic biopsy of Breast - right
C0942286|Guidance for stereotactic biopsy:Finding:Point in time:Breast.right:Document:Mam
C0942296|Guidance for placement of large bore catheter into vessel in Central vein - left
C0942296|Cent v-L LB Cath plac guid into ves
C0942296|Guidance for placement of large bore catheter into vessel:Find:Pt:Central vein.left:Doc
C0942296|Guidance for placement of large bore catheter into vessel:Finding:Point in time:Central vein.left:Document
C0942324|Brst-R Mam Bx guid
C0942324|Mammogram Guidance for biopsy of Breast - right
C0942324|Guidance for biopsy:Find:Pt:Breast.right:Doc:Mam
C0942324|Guidance for biopsy:Finding:Point in time:Breast.right:Document:Mam
C0942328|Mammogram Guidance for aspiration of cyst of Breast - left
C0942328|Brst-L Mam Cyst Asp guid
C0942328|Guidance for aspiration of cyst:Finding:Point in time:Breast.left:Document:Mam
C0942328|Guidance for aspiration of cyst:Find:Pt:Breast.left:Doc:Mam
C0882018|Lower leg MRI
C0882018|Multisection:Finding:Point in time:Lower leg:Document:MRI
C0882018|Multisection:Find:Pt:Lower leg:Doc:MRI
C0882043|Orbit-Bl CT W contr IV
C0882043|Orbit - bilateral CT W contrast IV
C0882043|Multisection^W contrast Intravenous:Finding:Point in time:Head>Orbit.bilateral:Document:Computerized Tomography
C0882043|Multisection^W contrast IV:Find:Pt:Head>Orbit.bilateral:Doc:CT
C0882045|Orbit-Bl MRI W contr IV
C0882045|Orbit - bilateral MRI W contrast IV
C0882045|Multisection^W contrast Intravenous:Finding:Point in time:Orbit.bilateral:Document:MRI
C0882045|Multisection^W contrast IV:Find:Pt:Orbit.bilateral:Doc:MRI
C0882071|US Guidance for biopsy of Prostate
C0882071|Prostate US Bx guid
C0882071|Guidance for biopsy:Finding:Point in time:Prostate:Document:Ultrasound
C0882071|Guidance for biopsy:Find:Pt:Prostate:Doc:US
C0882075|Pulm RI VP W 133Xe IH+Tc99mMAA IV
C0882075|Views ventilation & perfusion^W Xe-133 Inhalation & W Tc-99m MAA Intravenous:Finding:Point in time:Pulmonary system:Document:Radnuc
C0882075|Views ventilation & perfusion^W Xe-133 IH & W Tc-99m MAA IV:Find:Pt:Pulmonary system:Doc:Radnuc
C0882075|Pulmonary system Scan ventilation and perfusion W Xe-133 IH and W Tc-99m MAA IV
C0882086|Views:Finding:Point in time:Scapula:Narrative:XR
C0882086|Scapula XR
C0882086|Scapula X-ray
C0882086|Views:Find:Pt:Scapula:Doc:XR
C0882086|Views:Finding:Point in time:Scapula:Document:XR
C0882090|Should US
C0882090|Shoulder US
C0882090|Multisection:Find:Pt:Shoulder:Doc:US
C0882090|Multisection:Finding:Point in time:Shoulder:Document:Ultrasound
C0882564|XXX MRI.Angio W contr IV
C0882564|Unspecified body region MRI angiogram W contrast IV
C0882564|Multisection^W contrast IV:Find:Pt:XXX:Doc:MRI.angio
C0882564|Multisection^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:MRI.angio
C0882566|XXX Infusion port plac guide
C0882566|Guidance for placement of infusion port in Unspecified body region
C0882566|Guidance for placement of infusion port:Find:Pt:XXX:Doc
C0882566|Guidance for placement of infusion port:Finding:Point in time:To be specified in another part of the message:Document
C0942095|Views^W contrast IS:Find:Pt:Hip.right:Doc:XR.fluor
C0942095|Hip - right Fluoroscopy W contrast IS
C0942095|Hip-R Flr W contr IS
C0942095|Views^W contrast Intrasynovial:Finding:Point in time:Hip.right:Document:XR.fluor
C0942113|Scrotum+Test-R RI W Tc99mP IV
C0942113|Scrotum and Testicle - right Scan W Tc-99m pertechnetate IV
C0942113|Views^W Tc-99m pertechnetate Intravenous:Finding:Point in time:Scrotum+Testicle.right:Document:Radnuc
C0942113|Views^W Tc-99m pertechnetate IV:Find:Pt:Scrotum+Testicle.right:Doc:Radnuc
C0881798|US Guidance for drainage of Abdomen
C0881798|Abd US Drain guid
C0881798|Guidance for drainage:Find:Pt:Abdomen:Doc:US
C0881798|Guidance for drainage:Finding:Point in time:Abdomen:Document:Ultrasound
C0881821|TO ves MRI.Angio W contr IV
C0881821|Thoracic outlet vessels MRI angiogram W contrast IV
C0881821|Multisection^W contrast Intravenous:Finding:Point in time:Thoracic outlet vessels:Document:MRI.angio
C0881821|Multisection^W contrast IV:Find:Pt:Thoracic outlet vessels:Doc:MRI.angio
C0881895|US Guidance for biopsy of cyst of Unspecified body region
C0881895|XXX US Cyst Bx guid
C0881895|Guidance for biopsy of cyst:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C0881895|Guidance for biopsy of cyst:Find:Pt:XXX:Doc:US
C0881937|Liver Flr TJ Bx guid W contr IV
C0881937|Fluoroscopy Guidance for transjugular biopsy of Liver-- W contrast IV
C0881937|Guidance for biopsy.transjugular ^W contrast IV:Find:Pt:Liver:Doc:XR.fluor
C0881937|Guidance for biopsy.transjugular^W contrast Intravenous:Finding:Point in time:Liver:Document:XR.fluor
C0881952|Head.cistern CT W contr IT
C0881952|Multisection^W contrast Intrathecal:Finding:Point in time:Head>Cerebral cisterns:Document:Computerized Tomography
C0881952|Multisection^W contrast IT:Find:Pt:Head>Cerebral cisterns:Doc:CT
C0881952|Head Cerebral cist CT W contr IT
C0881952|Cerebral cisterns CT W contrast IT
C0882537|Joint RI W In-111 Intrajoint
C0882537|Joint Scan W In-111 intrajoint
C0882537|Views^W In-111 intrajoint:Find:Pt:Joint:Doc:Radnuc
C0882537|Views^W In-111 intrajoint:Finding:Point in time:Joint:Document:Radnuc
C0882538|Views^W radionuclide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C0882538|Kidney - bilateral Scan
C0882538|Views^W radionuclide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C0882538|Kdny-Bl RI W RNC IV
C1114516|Guidance for drainage:Finding:Point in time:To be specified in another part of the message:Narrative:ULTRASOUND
C1114516|US Guidance for drainage of Unspecified body region
C1114516|XXX US Drain guid
C1114516|Guidance for drainage:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1114516|Guidance for drainage:Find:Pt:XXX:Doc:US
C1114517|US Guidance for needle biopsy of Unspecified body region
C1114517|XXX US Bx needle guid
C1114517|Guidance for biopsy.needle:Find:Pt:XXX:Doc:US
C1114517|Guidance for biopsy.needle:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1114521|Uterus+FT US
C1114521|Uterus and Fallopian tubes US
C1114521|Multisection:Find:Pt:Uterus+Fallopian tubes:Doc:US
C1114521|Multisection:Finding:Point in time:Uterus+Fallopian tubes:Document:Ultrasound
C1114939|Zygomatic arch XR port
C1114939|Zygomatic arch X-ray portable
C1114939|Views portable:Find:Pt:Zygomatic arch:Doc:XR
C1114939|Views portable:Finding:Point in time:Zygomatic arch:Document:XR
C1114555|Chest XR PA+Lat+R-Obl+L-Obl
C1114555|Chest X-ray PA and lateral and right oblique and left oblique
C1114555|Views PA & lateral & R-oblique & L-oblique:Find:Pt:Chest:Doc:XR
C1114555|Views PA & lateral & R-oblique & L-oblique:Finding:Point in time:Chest:Document:XR
C1114570|Views^W contrast retrograde via urethra:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C1114570|Kidney - bilateral Fluoroscopy W contrast retrograde via urethra
C1114570|Views^W contrast retrograde via urethra:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C1114570|VIEWS^RETROGRADE VIA URETHRA:FINDING:POINT IN TIME:KIDNEYS AND COLLECTING SYSTEM:NARRATIVE:XR.FLUOR
C1114570|Kdny-Bl Flr W contr RU
C1114608|Abd ves CT.Angio WO+W contr IV
C1114608|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Vessels:Document:Computerized Tomography.angio
C1114608|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Vessels:Doc:CT.angio
C1114608|Abdominal vessels CT angiogram WO and W contrast IV
C1114621|Carot a.ext XRA W contr IA
C1114621|Carotid artery.external Fluoroscopic angiogram W contrast IA
C1114621|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.external:Document:XR.fluor.angio
C1114621|Views^W contrast IA:Find:Pt:Carotid artery.external:Doc:XR.fluor.angio
C1114629|IMA XRA W contr IA
C1114629|Internal mammary artery Fluoroscopic angiogram W contrast IA
C1114629|Views^W contrast IA:Find:Pt:Mammary artery.internal:Doc:XR.fluor.angio
C1114629|Views^W contrast Intra-arterial:Finding:Point in time:Mammary artery.internal:Document:XR.fluor.angio
C1114952|Adrenal artery - bilateral Fluoroscopic angiogram W contrast IA
C1114952|Adrenal a-Bl XRA W contr IA
C1114952|Views^W contrast Intra-arterial:Finding:Point in time:Adrenal artery.bilateral:Document:XR.fluor.angio
C1114952|Views^W contrast IA:Find:Pt:Adrenal artery.bilateral:Doc:XR.fluor.angio
C1114650|Extr lymph-Bl Flr W contr IL
C1114650|Extremity lymphatics - bilateral Fluoroscopy W contrast intra lymphatic
C1114650|Views^W contrast intra lymphatic:Finding:Point in time:Extremity lymphatics.bilateral:Document:XR.fluor
C1114650|Views^W contrast intra lymphatic:Find:Pt:Extremity lymphatics.bilateral:Doc:XR.fluor
C1114418|Orbit - bilateral CT WO contrast
C1114418|Orbit-Bl CT WO contr
C1114418|Multisection^WO contrast:Finding:Point in time:Head>Orbit.bilateral:Document:Computerized Tomography
C1114418|Multisection^WO contrast:Find:Pt:Head>Orbit.bilateral:Doc:CT
C1543423|Should-L XR AP(w IR+ER)+Ax+Y
C1543423|Shoulder - left X-ray AP (W internal rotation and W external rotation) and axillary and Y
C1543423|Views AP (W internal rotation & W external rotation) & axillary & Y:Find:Pt:Shoulder.left:Doc:XR
C1543423|Views AP (W internal rotation & W external rotation) & axillary & Y:Finding:Point in time:Shoulder.left:Document:XR
C1543492|Genitourinary system US
C1543492|GU US
C1543492|Multisection:Find:Pt:Genitourinary system:Doc:US
C1543492|Multisection:Finding:Point in time:Genitourinary system:Document:Ultrasound
C1543810|Stom RI GE W Tc99mSC PO
C1543810|Stomach Scan for gastric emptying W Tc-99m SC PO
C1543810|Views for gastric emptying ^W Tc-99m SC PO:Find:Pt:Stomach:Doc:Radnuc
C1543810|Views for gastric emptying^W Tc-99m Subcutaneous Oral:Finding:Point in time:Stomach:Document:Radnuc
C1543856|Bone Scan static limited
C1543856|Bone RI Static Ltd W RNC IV
C1543856|Views static limited ^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543856|Views static limited^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543860|Bone Scan whole body
C1543860|Bone RI WB W RNC IV
C1543860|Views whole body^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543860|Views whole body^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543865|Bone marrow SPECT
C1543865|BM SPECT W RNC IV
C1543865|Multisection^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc.SPECT
C1543865|Multisection^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc.SPECT
C1542902|RI Delayed W I-131 mIBG IV
C1542902|Scan delayed W I-131 MIBG IV
C1542902|Views delayed^W I-131 MIBG Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542902|Views delayed^W I-131 MIBG IV:Find:Pt:^Patient:Doc:Radnuc
C1543922|Salivary gland RI Static W RNC IV
C1543922|Salivary gland Scan static
C1543922|Views static^W radionuclide Intravenous:Finding:Point in time:Salivary gland:Document:Radnuc
C1543922|Views static^W radionuclide IV:Find:Pt:Salivary gland:Doc:Radnuc
C1543945|Hrt RI Gated+EF Rest+W RNC IV
C1543945|Heart Scan gated and ejection fraction at rest and W radionuclide IV
C1543945|Views gated & ejection fraction^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543945|Views gated & ejection fraction^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542857|Joint Scan limited
C1542857|Joint RI Ltd W RNC IV
C1542857|Views limited^W radionuclide Intravenous:Finding:Point in time:Joint:Document:Radnuc
C1542857|Views limited^W radionuclide IV:Find:Pt:Joint:Doc:Radnuc
C1543963|Prostate RI Mul Areas W Tc99mPMSA IV
C1543963|Prostate Scan multiple areas W Tc-99m capromab pendatide IV
C1543963|Views multiple areas^W Tc-99m capromab pendatide IV:Find:Pt:Prostate:Doc:Radnuc
C1543963|Views multiple areas^W Tc-99m capromab pendatide Intravenous:Finding:Point in time:Prostate:Document:Radnuc
C1543518|LE ves-R DOP
C1543518|Lower extremity vessels - right US.doppler
C1543518|Multisection:Find:Pt:Lower extremity vessels.right:Doc:US.doppler
C1543518|Multisection:Finding:Point in time:Lower extremity vessels.right:Document:Ultrasound.doppler
C1543158|UE MRI W contr IV
C1543158|Upper extremity MRI W contrast IV
C1543158|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity:Document:MRI
C1543158|Multisection^W contrast IV:Find:Pt:Upper extremity:Doc:MRI
C1543165|Head vessels US.doppler limited
C1543165|Head ves DOP Ltd
C1543165|Multisection limited:Finding:Point in time:Head vessels:Document:Ultrasound.doppler
C1543165|Multisection limited:Find:Pt:Head vessels:Doc:US.doppler
C1543177|Unspecified body region X-ray W manual stress
C1543177|XXX XR W Stress
C1543177|Views^W manual stress:Find:Pt:XXX:Doc:XR
C1543177|Views^W manual stress:Finding:Point in time:To be specified in another part of the message:Document:XR
C1543585|Pancreas transplant US
C1543585|Multisection:Finding:Point in time:Pancreas transplant:Document:Ultrasound
C1543585|Multisection:Find:Pt:Pancreas transplant:Doc:US
C1543597|US Guidance for biopsy of Lymph node
C1543597|LN US Bx guid
C1543597|Guidance for biopsy:Finding:Point in time:Lymph node:Document:Ultrasound
C1543597|Guidance for biopsy:Find:Pt:Lymph node:Doc:US
C1524265|Patella-R XR PA+Lat+Sunrise
C1524265|Patella - right X-ray PA and lateral and Sunrise
C1524265|Views PA & lateral & Sunrise:Find:Pt:Patella.right:Doc:XR
C1524265|Views PA & lateral & Sunrise:Finding:Point in time:Patella.right:Document:XR
C1524266|Should-R XR Grashey+Outlet
C1524266|Shoulder - right X-ray Grashey and outlet
C1524266|Views Grashey & outlet:Finding:Point in time:Shoulder.right:Document:XR
C1524266|Views Grashey & outlet:Find:Pt:Shoulder.right:Doc:XR
C1526765|Views^W contrast IA:Find:Pt:Upper extremity arteries.right:Nar:XR.fluor.angio
C1526765|Deprecated Upper extremity arteries Right X-ray fluoroscopy angio W contrast IA
C1526765|Deprecated UE aa-R XRA W contr IA
C1526765|Views^W contrast Intra-arterial:Finding:Point in time:Upper extremity arteries.right:Narrative:XR.fluor.angio
C1526767|Lymph Abd+Pelvic-R Flr W contr IL
C1526767|Lymphatics abdominal and Lymphatics pelvic - right Fluoroscopy W contrast intra lymphatic
C1526767|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.abdominal+Lymphatics.pelvic.right:Doc:XR.fluor
C1526767|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.abdominal+Lymphatics.pelvic.right:Document:XR.fluor
C1543730|Hrt SPECT W Stress+W RNC IV
C1543730|Heart SPECT W stress and W radionuclide IV
C1543730|Multisection^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543730|Multisection^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1542965|Lacrimal duct RI W RNC intra LD
C1542965|Lacrimal duct Scan W radionuclide intra lacrimal duct
C1542965|Views^W radionuclide intra lacrimal duct:Find:Pt:Lacrimal duct:Doc:Radnuc
C1542965|Views^W radionuclide intra lacrimal duct:Finding:Point in time:Lacrimal duct:Document:Radnuc
C1542968|Esophagus Scan for reflux W radionuclide PO
C1542968|Esoph RI for Reflux W RNC PO
C1542968|Views for reflux^W radionuclide PO:Find:Pt:Esophagus:Doc:Radnuc
C1542968|Views for reflux^W radionuclide Oral:Finding:Point in time:Esophagus:Document:Radnuc
C1526788|Upper extremity - left MRI WO contrast
C1526788|UE-L MRI WO contr
C1526788|Multisection^WO contrast:Find:Pt:Upper extremity.left:Doc:MRI
C1526788|Multisection^WO contrast:Finding:Point in time:Upper extremity.left:Document:MRI
C1526811|Brst-L Mam True Lat
C1526811|Breast - left Mammogram true lateral
C1526811|View true lateral:Find:Pt:Breast.left:Doc:Mam
C1526811|View true lateral:Finding:Point in time:Breast.left:Document:Mam
C1524186|Lower leg CT
C1524186|Multisection:Finding:Point in time:Lower leg:Document:Computerized Tomography
C1524186|Multisection:Find:Pt:Lower leg:Doc:CT
C1524816|Multisection^WO contrast:Finding:Point in time:Abdomen>Aorta.abdominal:Document:Computerized Tomography
C1524816|Multisection^WO contrast:Find:Pt:Abdomen>Aorta.abdominal:Doc:CT
C1524816|Abd Aorta CT WO contr
C1524816|Abdominal Aorta CT WO contrast
C1524817|Ab Ao MRI.Angio WO contr
C1524817|Aorta abdominal MRI angiogram WO contrast
C1524817|Multisection^WO contrast:Find:Pt:Aorta.abdominal:Doc:MRI.angio
C1524817|Multisection^WO contrast:Finding:Point in time:Aorta.abdominal:Document:MRI.angio
C1524831|Elbow-L MRI WO contr
C1524831|Elbow - left MRI WO contrast
C1524831|Multisection^WO contrast:Finding:Point in time:Elbow.left:Document:MRI
C1524831|Multisection^WO contrast:Find:Pt:Elbow.left:Doc:MRI
C1525179|Pulm ves MRI.Angio
C1525179|Pulmonary vessels MRI angiogram
C1525179|Multisection:Find:Pt:Pulmonary vessels:Doc:MRI.angio
C1525179|Multisection:Finding:Point in time:Pulmonary vessels:Document:MRI.angio
C1524465|Hip - left MRI W contrast IS
C1524465|Hip-L MRI W contr IS
C1524465|Multisection^W contrast IS:Find:Pt:Hip.left:Doc:MRI
C1524465|Multisection^W contrast Intrasynovial:Finding:Point in time:Hip.left:Document:MRI
C1525300|Wrist - bilateral X-ray W clenched fist
C1525300|Wrist-Bl XR W clenched fist
C1525300|View^W clenched fist:Find:Pt:Wrist.bilateral:Doc:XR
C1525300|View^W clenched fist:Finding:Point in time:Wrist.bilateral:Document:XR
C1525308|Foot X-ray Harris
C1525308|Ft XR Harris
C1525308|View Harris:Find:Pt:Foot:Doc:XR
C1525308|View Harris:Finding:Point in time:Foot:Document:XR
C1524232|Acromioclavicular joint - left X-ray Zanca
C1524232|AC joint-L XR Zanca
C1524232|View Zanca:Finding:Point in time:Acromioclavicular joint.left:Document:XR
C1524232|View Zanca:Find:Pt:Acromioclavicular joint.left:Doc:XR
C1525480|Ft-L XR 2V stand
C1525480|Foot - left X-ray 2 views standing
C1525480|Views 2^standing:Finding:Point in time:Foot.left:Document:XR
C1525480|Views 2^standing:Find:Pt:Foot.left:Doc:XR
C1525487|Abd XR AP(sup+Lat Decub) Port
C1525487|Abdomen X-ray AP (supine and lateral-decubitus) portable
C1525487|Views AP (supine & lateral-decubitus) portable:Finding:Point in time:Abdomen:Document:XR
C1525487|Views AP (supine & lateral-decubitus) portable:Find:Pt:Abdomen:Doc:XR
C1525501|Knee XR AP+Lat Xtable
C1525501|Knee X-ray AP and lateral crosstable
C1525501|Views AP & lateral crosstable:Finding:Point in time:Knee:Document:XR
C1525501|Views AP & lateral crosstable:Find:Pt:Knee:Doc:XR
C1525526|Should-Bl XR AP+Ax+Y
C1525526|Shoulder - bilateral X-ray AP and axillary and Y
C1525526|Views AP & axillary & Y:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525526|Views AP & axillary & Y:Find:Pt:Shoulder.bilateral:Doc:XR
C1525558|Foot - left X-ray tarsal
C1525558|Ft-L XR Tarsal
C1525558|Views tarsal:Finding:Point in time:Foot.left:Document:XR
C1525558|Views tarsal:Find:Pt:Foot.left:Doc:XR
C1525560|Should-Bl XR Grashey+Ax+Outlet+Zanca
C1525560|Shoulder - bilateral X-ray Grashey and axillary and outlet and Zanca
C1525560|Views Grashey & axillary & outlet & Zanca:Find:Pt:Shoulder.bilateral:Doc:XR
C1525560|Views Grashey & axillary & outlet & Zanca:Finding:Point in time:Shoulder.bilateral:Document:XR
C1525617|XXX CT for fistula
C1525617|Multisection for fistula:Find:Pt:XXX:Doc:CT
C1525617|Unspecified body region CT for fistula
C1525617|Multisection for fistula:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1525627|LS-spine junc CT
C1525627|Spine Lumbosacral Junction CT
C1525627|Multisection:Find:Pt:Spine.lumbosacral junction:Doc:CT
C1525627|Multisection:Finding:Point in time:Spine.lumbosacral junction:Document:Computerized Tomography
C1525633|Brain+IAC MRI W contr IV
C1525633|Brain and Internal auditory canal MRI W contrast IV
C1525633|Multisection^W contrast IV:Find:Pt:Brain+Internal auditory canal:Doc:MRI
C1525633|Multisection^W contrast Intravenous:Finding:Point in time:Brain+Internal auditory canal:Document:MRI
C1525651|Parotid gland MRI WO and W contrast IV
C1525651|Multisection^WO & W contrast IV:Find:Pt:Parotid gland:Doc:MRI
C1525651|Parotid gland MRI WO+W contr IV
C1525651|Multisection^WO & W contrast Intravenous:Finding:Point in time:Parotid gland:Document:MRI
C1525662|Parotid gland CT WO contrast
C1525662|Parotid gland CT WO contr
C1525662|Multisection^WO contrast:Finding:Point in time:Parotid gland:Document:Computerized Tomography
C1525662|Multisection^WO contrast:Find:Pt:Parotid gland:Doc:CT
C1525663|Parotid gland MRI WO contrast
C1525663|Parotid gland MRI WO contr
C1525663|Multisection^WO contrast:Finding:Point in time:Parotid gland:Document:MRI
C1525663|Multisection^WO contrast:Find:Pt:Parotid gland:Doc:MRI
C1525739|UE vv-Bl XRA W contr IV
C1525739|Upper extremity veins - bilateral Fluoroscopic angiogram W contrast IV
C1525739|Views^W contrast IV:Find:Pt:Upper extremity veins.bilateral:Doc:XR.fluor.angio
C1525739|Views^W contrast Intravenous:Finding:Point in time:Upper extremity veins.bilateral:Document:XR.fluor.angio
C1525791|Lower extremity arteries Fluoroscopic angiogram W contrast IA
C1525791|LE aa XRA W contr IA
C1525791|Views^W contrast IA:Find:Pt:Lower extremity arteries:Doc:XR.fluor.angio
C1525791|Views^W contrast Intra-arterial:Finding:Point in time:Lower extremity arteries:Document:XR.fluor.angio
C1525874|Acromioclavicular joint - bilateral X-ray W weight
C1525874|AC joint-Bl XR W Wt
C1525874|Views^W weight:Find:Pt:Acromioclavicular joint.bilateral:Doc:XR
C1525874|Views^W weight:Finding:Point in time:Acromioclavicular joint.bilateral:Document:XR
C1524134|Ac arch+Carot a.ext-Bl XRA W contr IA
C1524134|Aortic arch and Carotid artery.external - bilateral Fluoroscopic angiogram W contrast IA
C1524134|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery.external.bilateral:Document:XR.fluor.angio
C1524134|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery.external.bilateral:Doc:XR.fluor.angio
C1525888|Nasal bones X-ray 3 views
C1525888|Nasal bones XR 3V
C1525888|Views 3:Find:Pt:Nasal bones:Doc:XR
C1525888|Views 3:Finding:Point in time:Nasal bones:Document:XR
C1525934|View 1:Finding:Point in time:Pelvis:Narrative:XR
C1525934|Pelvis X-ray Single view
C1525934|Pelvis XR 1V
C1525934|View 1:Finding:Point in time:Pelvis:Document:XR
C1525934|View 1:Find:Pt:Pelvis:Doc:XR
C1525940|Pelvis X-ray AP single view
C1525940|Pelvis XR AP 1V
C1525940|View AP:Find:Pt:Pelvis:Doc:XR
C1525940|View AP:Finding:Point in time:Pelvis:Document:XR
C1525821|Finger.5th-L XR
C1525821|Finger fifth - left X-ray
C1525821|Views:Find:Pt:Finger.fifth.left:Doc:XR
C1525821|Views:Finding:Point in time:Finger.fifth.left:Document:XR
C1525952|Pelvis X-ray AP 20 degree cephalic angle
C1525952|Pelvis XR AP 20 Deg Ceph Angle
C1525952|View AP 20 degree cephalic angle:Find:Pt:Pelvis:Doc:XR
C1525952|View AP 20 degree cephalic angle:Finding:Point in time:Pelvis:Document:XR
C1525959|Wrist-R XR Ltd
C1525959|Wrist - right X-ray limited
C1525959|Views limited:Finding:Point in time:Wrist.right:Document:XR
C1525959|Views limited:Find:Pt:Wrist.right:Doc:XR
C1526006|Femur-R XR 2V
C1526006|Femur - right X-ray 2 views
C1526006|Views 2:Find:Pt:Femur.right:Doc:XR
C1526006|Views 2:Finding:Point in time:Femur.right:Document:XR
C1526015|Ft-R XR 3V
C1526015|Foot - right X-ray 3 views
C1526015|Views 3:Finding:Point in time:Foot.right:Document:XR
C1526015|Views 3:Find:Pt:Foot.right:Doc:XR
C1526020|Foot - right X-ray oblique single view
C1526020|Ft-R XR Obl 1V
C1526020|View oblique:Find:Pt:Foot.right:Doc:XR
C1526020|View oblique:Finding:Point in time:Foot.right:Document:XR
C1526022|Ft-R XRTomo
C1526022|Foot - right X-ray tomograph
C1526022|Multisection:Find:Pt:Foot.right:Doc:XR.tomo
C1526022|Multisection:Finding:Point in time:Foot.right:Document:XR.tomo
C1526026|Hand-R XR AP+Lat
C1526026|Hand - right X-ray AP and lateral
C1526026|Views AP & lateral:Find:Pt:Hand.right:Doc:XR
C1526026|Views AP & lateral:Finding:Point in time:Hand.right:Document:XR
C1526106|Shoulder - right X-ray Garth
C1526106|Should-R XR Garth
C1526106|View Garth:Find:Pt:Shoulder.right:Doc:XR
C1526106|View Garth:Finding:Point in time:Shoulder.right:Document:XR
C1526132|Shoulder X-ray 2 views
C1526132|Should XR 2V
C1526132|Views 2:Find:Pt:Shoulder:Doc:XR
C1526132|Views 2:Finding:Point in time:Shoulder:Document:XR
C1526087|Ribs-R XR Ant+Lat
C1526087|Ribs - right X-ray anterior and lateral
C1526087|Views anterior & lateral:Finding:Point in time:Ribs.right:Document:XR
C1526087|Views anterior & lateral:Find:Pt:Ribs.right:Doc:XR
C1526096|Should-R XR Stryker Notch
C1526096|Shoulder - right X-ray Stryker Notch
C1526096|View Stryker Notch:Finding:Point in time:Shoulder.right:Document:XR
C1526096|View Stryker Notch:Find:Pt:Shoulder.right:Doc:XR
C1526159|Skull XR 2V
C1526159|Skull X-ray 2 views
C1526159|Views 2:Find:Pt:Skull:Doc:XR
C1526159|Views 2:Finding:Point in time:Skull:Document:XR
C1526162|Skull XR Towne
C1526162|Skull X-ray Towne
C1526162|View Towne:Find:Pt:Skull:Doc:XR
C1526162|View Towne:Finding:Point in time:Skull:Document:XR
C1525917|Scrotum+Test US Bx guid
C1525917|US Guidance for biopsy of Scrotum and Testicle
C1525917|Guidance for biopsy:Finding:Point in time:Scrotum+Testicle:Document:Ultrasound
C1525917|Guidance for biopsy:Find:Pt:Scrotum+Testicle:Doc:US
C1525148|Finger third - right X-ray
C1525148|Finger.3rd-R XR
C1525148|Views:Find:Pt:Finger.third.right:Doc:XR
C1525148|Views:Finding:Point in time:Finger.third.right:Document:XR
C1526327|Kidney-R Flr W contr RU
C1526327|Kidney - right Fluoroscopy W contrast retrograde via urethra
C1526327|Views^W contrast retrograde via urethra:Finding:Point in time:Kidney.right:Document:XR.fluor
C1526327|Views^W contrast retrograde via urethra:Find:Pt:Kidney.right:Doc:XR.fluor
C1524470|Knee-L MRI W contr IS
C1524470|Multisection^W contrast Intrasynovial:Finding:Point in time:Knee.left:Document:MRI
C1524470|Multisection^W contrast IS:Find:Pt:Knee.left:Doc:MRI
C1524470|Knee - left MRI W contrast IS
C1524479|Ankle CT W contr IV
C1524479|Ankle CT W contrast IV
C1524479|Multisection^W contrast Intravenous:Finding:Point in time:Ankle:Document:Computerized Tomography
C1524479|Multisection^W contrast IV:Find:Pt:Ankle:Doc:CT
C1524493|Brst MRI W contr IV
C1524493|Breast MRI W contrast IV
C1524493|Multisection^W contrast Intravenous:Finding:Point in time:Breast:Document:MRI
C1524493|Multisection^W contrast IV:Find:Pt:Breast:Doc:MRI
C1524869|Hip CT WO contrast
C1524869|Hip CT WO contr
C1524869|Multisection^WO contrast:Finding:Point in time:Hip:Document:Computerized Tomography
C1524869|Multisection^WO contrast:Find:Pt:Hip:Doc:CT
C1524536|Hand MRI W contr IV
C1524536|Hand MRI W contrast IV
C1524536|Multisection^W contrast IV:Find:Pt:Hand:Doc:MRI
C1524536|Multisection^W contrast Intravenous:Finding:Point in time:Hand:Document:MRI
C1524167|Hip-Bl CT W contr IV
C1524167|Hip - bilateral CT W contrast IV
C1524167|Multisection^W contrast Intravenous:Finding:Point in time:Hip.bilateral:Document:Computerized Tomography
C1524167|Multisection^W contrast IV:Find:Pt:Hip.bilateral:Doc:CT
C1524169|Hip-L CT W contr IV
C1524169|Hip - left CT W contrast IV
C1524169|Multisection^W contrast Intravenous:Finding:Point in time:Hip.left:Document:Computerized Tomography
C1524169|Multisection^W contrast IV:Find:Pt:Hip.left:Doc:CT
C1524590|Spine MRI W contr IV
C1524590|Spine MRI W contrast IV
C1524590|Multisection^W contrast Intravenous:Finding:Point in time:Spine:Document:MRI
C1524590|Multisection^W contrast IV:Find:Pt:Spine:Doc:MRI
C1524613|Elbow - right CT WO and W contrast IV
C1524613|Multisection^WO & W contrast IV:Find:Pt:Elbow.right:Doc:CT
C1524613|Multisection^WO & W contrast Intravenous:Finding:Point in time:Elbow.right:Document:Computerized Tomography
C1524613|Elbow-R CT WO+W contr IV
C1524617|Lower extremity - left MRI WO and W contrast IV
C1524617|Multisection^WO & W contrast IV:Find:Pt:Lower extremity.left:Doc:MRI
C1524617|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity.left:Document:MRI
C1524617|LE-L MRI WO+W contr IV
C1524948|Hand - bilateral X-ray lateral
C1524948|Hand-Bl XR Lat
C1524948|View lateral:Find:Pt:Hand.bilateral:Doc:XR
C1524948|View lateral:Finding:Point in time:Hand.bilateral:Document:XR
C1524953|Knee-Bl XR Lat
C1524953|Knee - bilateral X-ray lateral
C1524953|View lateral:Finding:Point in time:Knee.bilateral:Document:XR
C1524953|View lateral:Find:Pt:Knee.bilateral:Doc:XR
C1524312|Abd CT Drain guid
C1524312|CT Guidance for drainage of Abdomen
C1524312|Guidance for drainage:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524312|Guidance for drainage:Find:Pt:Abdomen:Doc:CT
C1525001|Femur - bilateral X-ray 2 views
C1525001|Femur-Bl XR 2V
C1525001|Views 2:Finding:Point in time:Femur.bilateral:Document:XR
C1525001|Views 2:Find:Pt:Femur.bilateral:Doc:XR
C1525023|Ankle-Bl XR AP+Lat
C1525023|Ankle - bilateral X-ray AP and lateral
C1525023|Views AP & lateral:Find:Pt:Ankle.bilateral:Doc:XR
C1525023|Views AP & lateral:Finding:Point in time:Ankle.bilateral:Document:XR
C1524756|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper arm.right:Document:MRI
C1524756|Upper arm-R MRI WO+W contr IV
C1524756|Multisection^WO & W contrast IV:Find:Pt:Upper arm.right:Doc:MRI
C1524756|Upper arm - right MRI WO and W contrast IV
C1525029|Elbow-Bl XR AP+Lat
C1525029|Elbow - bilateral X-ray AP and lateral
C1525029|Views AP & lateral:Find:Pt:Elbow.bilateral:Doc:XR
C1525029|Views AP & lateral:Finding:Point in time:Elbow.bilateral:Document:XR
C1525038|Radius+Ulna-Bl XR AP+Lat
C1525038|Radius - bilateral and Ulna - bilateral X-ray AP and lateral
C1525038|Views AP & lateral:Finding:Point in time:Radius.bilateral+Ulna.bilateral:Document:XR
C1525038|Views AP & lateral:Find:Pt:Radius.bilateral+Ulna.bilateral:Doc:XR
C1525050|Mandible XR AP+Lat
C1525050|Mandible X-ray AP and lateral
C1525050|Views AP & lateral:Finding:Point in time:Mandible:Document:XR
C1525050|Views AP & lateral:Find:Pt:Mandible:Doc:XR
C1525053|Scapula-Bl XR AP+Lat
C1525053|Scapula - bilateral X-ray AP and lateral
C1525053|Views AP & lateral:Finding:Point in time:Scapula.bilateral:Document:XR
C1525053|Views AP & lateral:Find:Pt:Scapula.bilateral:Doc:XR
C1524399|Wrist+Hand MRI
C1524399|Wrist and Hand MRI
C1524399|Multisection:Finding:Point in time:Wrist+Hand:Document:MRI
C1524399|Multisection:Find:Pt:Wrist+Hand:Doc:MRI
C1524413|Humerus X-ray tomograph
C1524413|Humerus XRTomo
C1524413|Multisection:Finding:Point in time:Humerus:Document:XR.tomo
C1524413|Multisection:Find:Pt:Humerus:Doc:XR.tomo
C1524785|Spine MRI WO and W contrast IV
C1524785|Spine MRI WO+W contr IV
C1524785|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine:Document:MRI
C1524785|Multisection^WO & W contrast IV:Find:Pt:Spine:Doc:MRI
C1524797|Multisection^WO & W contrast IV:Find:Pt:Lower leg.right:Doc:MRI
C1524797|Lower leg - right MRI WO and W contrast IV
C1524797|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower leg.right:Document:MRI
C1524797|Lower leg-R MRI WO+W contr IV
C1525089|BDs Flr Balloon dilatation W contr
C1525089|Biliary ducts Fluoroscopy Balloon dilatation W contrast
C1525089|Balloon dilatation^W contrast:Find:Pt:Biliary ducts:Doc:XR.fluor
C1525089|Balloon dilatation^W contrast:Finding:Point in time:Biliary ducts:Document:XR.fluor
C1830190|Guidance for biopsy^WO & W contrast IV:Find:Pt:XXX:Doc:CT
C1830190|CT Guidance for biopsy of Unspecified body region-- WO and W contrast IV
C1830190|XXX CT Bx guid WO+W contr IV
C1830190|Guidance for biopsy^WO & W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1830233|Orbit+Face+Neck MRI WO contr
C1830233|Orbit and Face and Neck MRI WO contrast
C1830233|Multisection^WO contrast:Find:Pt:Orbit+Face+Neck:Doc:MRI
C1830233|Multisection^WO contrast:Finding:Point in time:Orbit+Face+Neck:Document:MRI
C1830243|Breast FFD mammogram
C1830243|Brst FFDM
C1830243|Views:Find:Pt:Breast:Doc:Mam.FFD
C1830243|Views:Finding:Point in time:Breast:Document:Mam.FFD
C1830265|Lower extremity vein - bilateral US
C1830265|LE v-Bl US
C1830265|Multisection:Find:Pt:Lower extremity vein.bilateral:Doc:US
C1830265|Multisection:Finding:Point in time:Lower extremity vein.bilateral:Document:Ultrasound
C1830280|Should XR port
C1830280|Shoulder X-ray portable
C1830280|Views portable:Finding:Point in time:Shoulder:Document:XR
C1830280|Views portable:Find:Pt:Shoulder:Doc:XR
C1830284|Hrt SPECT Gated+EF Rest+stress+W RNC IV
C1830284|Heart SPECT gated and ejection fraction at rest and W stress and W radionuclide IV
C1830284|Multisection gated & ejection fraction^at rest & W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1830284|Multisection gated & ejection fraction^at rest & W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1715381|Muscle CT Guidance for deep biopsy
C1715381|CT Guidance for deep biopsy of Muscle
C1715381|Guidance for deep biopsy:Find:Pt:Muscle:Doc:CT
C1715381|Guidance for deep biopsy:Finding:Point in time:Muscle:Document:Computerized Tomography
C1632803|Views frontal stereo:Finding:Point in time:Chest:Narrative:XR
C1632803|Chest X-ray frontal stereo
C1632803|Chest XR Frontal Stereo
C1632803|Views frontal stereo:Find:Pt:Chest:Doc:XR
C1632803|Views frontal stereo:Finding:Point in time:Chest:Document:XR
C1714530|Thumb-L XR GE 3V
C1714530|Thumb - left X-ray GE 3 views
C1714530|Views GE 3:Find:Pt:Thumb.left:Doc:XR
C1714530|Views GE 3:Finding:Point in time:Thumb.left:Document:XR
C1714899|Knee-L XR GE 3V
C1714899|Knee - left X-ray GE 3 views
C1714899|Views GE 3:Find:Pt:Knee.left:Doc:XR
C1714899|Views GE 3:Finding:Point in time:Knee.left:Document:XR
C1714905|Axilla-L MRI W contr IV
C1714905|Axilla - left MRI W contrast IV
C1714905|Multisection^W contrast IV:Find:Pt:Axilla.left:Doc:MRI
C1714905|Multisection^W contrast Intravenous:Finding:Point in time:Axilla.left:Document:MRI
C1717257|Thigh ves-R MRI.Angio WO contr
C1717257|Thigh vessels - right MRI angiogram WO contrast
C1717257|Multisection^WO contrast:Find:Pt:Thigh vessels.right:Doc:MRI.angio
C1717257|Multisection^WO contrast:Finding:Point in time:Thigh vessels.right:Document:MRI.angio
C1715037|Thyroid SPECT flow
C1715037|Thyroid SPECT Flow W RNC IV
C1715037|Multisection flow^W radionuclide IV:Find:Pt:Thyroid:Doc:Radnuc.SPECT
C1715037|Multisection flow^W radionuclide Intravenous:Finding:Point in time:Thyroid:Document:Radnuc.SPECT
C1637282|Brst-R Mam Bx CN Str Guid
C1637282|Guidance for stereotactic biopsy.core needle:Find:Pt:Breast.right:Doc:Mam
C1637282|Guidance for stereotactic biopsy.core needle:Finding:Point in time:Breast.right:Document:Mam
C1637282|Mammogram Guidance for stereotactic core needle biopsy of Breast - right
C1636074|Pelvis US transabdominal and transvaginal
C1636074|Pelvis US Transabdom+Transvag
C1636074|Multisection transabdominal & transvaginal:Find:Pt:Pelvis:Doc:US
C1636074|Multisection transabdominal & transvaginal:Finding:Point in time:Pelvis:Document:Ultrasound
C1642564|Pelvis vessels US.doppler limited
C1642564|Pelvis ves DOP Ltd
C1642564|Multisection limited:Finding:Point in time:Pelvis vessels:Document:Ultrasound.doppler
C1642564|Multisection limited:Find:Pt:Pelvis vessels:Doc:US.doppler
C1642087|Femur-R XR port
C1642087|Femur - right X-ray portable
C1642087|Views portable:Finding:Point in time:Femur.right:Document:XR
C1642087|Views portable:Find:Pt:Femur.right:Doc:XR
C1632986|Chest CT Abscess drain guid
C1632986|Guidance for drainage of abscess:Find:Pt:Chest:Doc:CT
C1632986|Guidance for drainage of abscess:Finding:Point in time:Chest:Document:Computerized Tomography
C1632986|CT Guidance for drainage of abscess of Chest
C1954375|Sacroiliac joint - bilateral X-ray GE 3 views
C1954375|SIJ-Bl XR GE 3V
C1954375|Views GE 3:Finding:Point in time:Sacroiliac joint.bilateral:Document:XR
C1954375|Views GE 3:Find:Pt:Sacroiliac joint.bilateral:Doc:XR
C1953325|Views:Finding:Point in time:Pelvis+Spine.lumbar:Narrative:XR
C1953325|Pelvis+L-spine XR
C1953325|Pelvis and Spine Lumbar X-ray
C1953325|Views:Find:Pt:Pelvis+Spine.lumbar:Doc:XR
C1953325|Views:Finding:Point in time:Pelvis+Spine.lumbar:Document:XR
C1953978|Mastoid - right X-ray 3 views
C1953978|Mastoid-R XR 3V
C1953978|Views 3:Find:Pt:Mastoid.right:Doc:XR
C1953978|Views 3:Finding:Point in time:Mastoid.right:Document:XR
C1953993|Ribs - bilateral and Chest X-ray GE 3 and PA Chest views
C1953993|Views GE 3 & PA chest:Finding:Point in time:Ribs.bilateral+Chest:Document:XR
C1953993|Views GE 3 & PA chest:Find:Pt:Ribs.bilateral+Chest:Doc:XR
C1953993|Ribs-Bl+Chest XR GE 3V+PA Chst
C1952656|TMJ-R XR Open+Closed Mouth
C1952656|Temporomandibular joint - right X-ray open and closed mouth
C1952656|Views open & closed mouth:Find:Pt:Temporomandibular joint.right:Doc:XR
C1952656|Views open & closed mouth:Finding:Point in time:Temporomandibular joint.right:Document:XR
C2925706|Head+Neck PET
C2925706|Head and Neck PET
C2925706|Multisection:Finding:Point in time:Head+Neck:Document:Radnuc.PET
C2925706|Multisection:Find:Pt:Head+Neck:Doc:Radnuc.PET
C3174152|Lung - left X-ray W contrast intrabronchial
C3174152|Lung-L XR W contr IB
C3174152|Views^W contrast intrabronchial:Finding:Point in time:Lung.left:Document:XR
C3174152|Views^W contrast intrabronchial:Find:Pt:Lung.left:Doc:XR
C3174366|Kidney - bilateral Fluoroscopy View for cyst examination
C3174366|View for cyst examination:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C3174366|View for cyst examination:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C3174366|Kdny-Bl Flr View for cyst exam
C3169530|Extr-R US Ltd
C3169530|Extremity - right US limited
C3169530|Multisection limited:Find:Pt:Extremity.right:Doc:US
C3169530|Multisection limited:Finding:Point in time:Extremity.right:Document:Ultrasound
C3533565|Extr v-Bl US Sclerosing agent inj guid
C3533565|US Guidance for injection of sclerosing agent of Extremity vein - bilateral
C3533565|Guidance for injection of sclerosing agent:Find:Pt:Extremity vein.bilateral:Doc:US
C3533565|Guidance for injection of sclerosing agent:Finding:Point in time:Extremity vein.bilateral:Document:Ultrasound
C3533791|Multisection^W contrast Intravenous:Finding:Point in time:Aorta+Femoral artery.bilateral:Document:Computerized Tomography.angio
C3533791|Deprecated Aorta and Femoral artery - bilateral CT angiogram W contrast IV
C3533791|Multisection^W contrast IV:Find:Pt:Aorta+Femoral artery.bilateral:Doc:CT.angio
C3533791|Deprecated Aorta+Fem a-Bl CT.Angio W con
C3262961|Hip - left X-ray Danelius Miller
C3262961|Hip-L XR Danelius Miller
C3262961|View Danelius Miller:Find:Pt:Hip.left:Doc:XR
C3262961|View Danelius Miller:Finding:Point in time:Hip.left:Document:XR
C3262981|Circle of Willis MRI angiogram WO and W contrast IV
C3262981|Circle of Willis MRI.Angio WO+W contr IV
C3262981|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head+Neck>Circle of Willis:Document:MRI.angio
C3262981|Multisection^WO & W contrast IV:Find:Pt:Head+Neck>Circle of Willis:Doc:MRI.angio
C3482444|Deprecated Spine Cervical CT stereotactic
C3482444|Multisection stereotactic:Find:Pt:Spine.cervical:Doc:CT
C3482444|Deprecated C-spine CT Stereo
C3482444|Multisection stereotactic:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C3263089|US Guidance for needle biopsy of Pancreas
C3263089|Pancreas US Bx needle guid
C3263089|Guidance for biopsy.needle:Finding:Point in time:Pancreas:Document:Ultrasound
C3263089|Guidance for biopsy.needle:Find:Pt:Pancreas:Doc:US
C3261472|Tib+Fib-L XR 1V
C3261472|Tibia - left and Fibula - left X-ray Single view
C3261472|View 1:Finding:Point in time:Tibia.left+Fibula.left:Document:XR
C3261472|View 1:Find:Pt:Tibia.left+Fibula.left:Doc:XR
C3261474|Elbow - right X-ray Single view
C3261474|Elbow-R XR 1V
C3261474|View 1:Finding:Point in time:Elbow.right:Document:XR
C3261474|View 1:Find:Pt:Elbow.right:Doc:XR
C3262883|Knee-Bl XR 2V+Sunrise
C3262883|Knee - bilateral X-ray 2 views and Sunrise
C3262883|Views 2 & Sunrise:Find:Pt:Knee.bilateral:Doc:XR
C3262883|Views 2 & Sunrise:Finding:Point in time:Knee.bilateral:Document:XR
C3262886|Knee - bilateral X-ray 4 views and Sunrise and tunnel
C3262886|Knee-Bl XR 4V+Sunrise+Tunnel
C3262886|Views 4 & Sunrise & tunnel:Find:Pt:Knee.bilateral:Doc:XR
C3262886|Views 4 & Sunrise & tunnel:Finding:Point in time:Knee.bilateral:Document:XR
C3262899|Fluoroscopy Guidance for biopsy of Bone
C3262899|Bone Flr Bx guid
C3262899|Guidance for biopsy:Finding:Point in time:Bone:Document:XR.fluor
C3262899|Guidance for biopsy:Find:Pt:Bone:Doc:XR.fluor
C0942167|Should-Bl XR
C0942167|Shoulder - bilateral X-ray
C0942167|Views:Finding:Point in time:Shoulder.bilateral:Document:XR
C0942167|Views:Find:Pt:Shoulder.bilateral:Doc:XR
C0945322|Breast - right US
C0945322|Brst-R US
C0945322|Multisection:Find:Pt:Breast.right:Doc:US
C0945322|Multisection:Finding:Point in time:Breast.right:Document:Ultrasound
C0945326|Finger-Bl MRI
C0945326|Finger - bilateral MRI
C0945326|Multisection:Find:Pt:Finger.bilateral:Doc:MRI
C0945326|Multisection:Finding:Point in time:Finger.bilateral:Document:MRI
C0942264|Shoulder - right US
C0942264|Should-R US
C0942264|Multisection:Finding:Point in time:Shoulder.right:Document:Ultrasound
C0942264|Multisection:Find:Pt:Shoulder.right:Doc:US
C0942280|Breast - bilateral US limited
C0942280|Brst-Bl US Ltd
C0942280|Multisection limited:Finding:Point in time:Breast.bilateral:Document:Ultrasound
C0942280|Multisection limited:Find:Pt:Breast.bilateral:Doc:US
C0942308|CT Guidance for injection of Sacroiliac joint - right
C0942308|SIJ-R CT Inj guid
C0942308|Guidance for injection:Find:Pt:Sacroiliac joint.right:Doc:CT
C0942308|Guidance for injection:Finding:Point in time:Sacroiliac joint.right:Document:Computerized Tomography
C0942338|Hand-L XR Arthritis
C0942338|Hand - left X-ray arthritis
C0942338|View arthritis:Find:Pt:Hand.left:Doc:XR
C0942338|View arthritis:Finding:Point in time:Hand.left:Document:XR
C0882023|Lymphatics Fluoroscopy W contrast intra lymphatic
C0882023|Lymph Flr W contr IL
C0882023|Views^W contrast intra lymphatic:Find:Pt:Lymphatics:Doc:XR.fluor
C0882023|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics:Document:XR.fluor
C0882542|Mesenteric artery Fluoroscopic angiogram Angioplasty W contrast IA
C0882542|Mesenteric a XRA Angpsty W contr IA
C0882542|Angioplasty^W contrast IA:Find:Pt:Mesenteric artery:Doc:XR.fluor.angio
C0882542|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Mesenteric artery:Document:XR.fluor.angio
C0882057|Pelvis CT
C0882057|Multisection:Finding:Point in time:Pelvis:Narrative:Computerized Tomography
C0882057|Multisection:Find:Pt:Pelvis:Doc:CT
C0882057|Multisection:Finding:Point in time:Pelvis:Document:Computerized Tomography
C0882060|Pelvis US
C0882060|Multisection:Find:Pt:Pelvis:Doc:US
C0882060|Multisection:Finding:Point in time:Pelvis:Document:Ultrasound
C0882079|Rectum Flr p contr PR during def
C0882079|Rectum Fluoroscopy post contrast PR during defecation
C0882079|View^post contrast PR during defecation:Find:Pt:Rectum:Doc:XR.fluor
C0882079|View^post contrast Rectal during defecation:Finding:Point in time:Rectum:Document:XR.fluor
C0882112|Spine facet joint Flr Inj guid
C0882112|Fluoroscopy Guidance for injection of Spine facet joint
C0882112|Guidance for injection:Finding:Point in time:Spine facet joint:Document:XR.fluor
C0882112|Guidance for injection:Find:Pt:Spine facet joint:Doc:XR.fluor
C0882133|L-spine XR W FE
C0882133|Views^W flexion & W extension:Find:Pt:Spine.lumbar:Doc:XR
C0882133|Views^W flexion & W extension:Finding:Point in time:Spine.lumbar:Document:XR
C0882133|Lumbar spine X-ray W flexion and W extension
C0882137|L-spine+SIJ-Bl XR
C0882137|Spine.lumbar and Sacroiliac joint - bilateral X-ray
C0882137|Views:Finding:Point in time:Spine.lumbar+Sacroiliac joint.bilateral:Document:XR
C0882137|Views:Find:Pt:Spine.lumbar+Sacroiliac joint.bilateral:Doc:XR
C0882143|T-spine XR
C0882143|Views:Find:Pt:Spine.thoracic:Doc:XR
C0882143|Views:Finding:Point in time:Spine.thoracic:Document:XR
C0882143|Thoracic spine X-ray
C0882158|Placement check of gastrostomy tube W contrast via GI tube
C0882158|Flr GT plac Ck W contr via GI tb
C0882158|Placement check of gastrostomy tube^W contrast via GI tube:Find:Pt:Stomach:Doc:XR.fluor
C0882158|Placement check of gastrostomy tube^W contrast via GI tube:Finding:Point in time:Stomach:Document:XR.fluor
C2718102|Deprecated Thigh MRI Multisection
C2718102|Deprecated Thigh MRI
C2718102|Multisection:Find:Pt:Thigh:Nar:MRI
C2718102|Multisection:Finding:Point in time:Thigh:Narrative:MRI
C0882207|XXX CT Radiosurg guid
C0882207|CT Guidance for radiosurgery of Unspecified body region
C0882207|Guidance for radiosurgery:Find:Pt:XXX:Doc:CT
C0882207|Guidance for radiosurgery:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0942126|Clavicle-Bl XR
C0942126|Clavicle - bilateral X-ray
C0942126|Views:Find:Pt:Clavicle.bilateral:Doc:XR
C0942126|Views:Finding:Point in time:Clavicle.bilateral:Document:XR
C0881872|Chest XR PA+Lat Upr port
C0881872|Chest X-ray PA and lateral upright portable
C0881872|Views PA & lateral upright portable:Finding:Point in time:Chest:Document:XR
C0881872|Views PA & lateral upright portable:Find:Pt:Chest:Doc:XR
C0881945|Head CT W contr IV
C0881945|Head CT W contrast IV
C0881945|Multisection^W contrast Intravenous:Finding:Point in time:Head:Document:Computerized Tomography
C0881945|Multisection^W contrast IV:Find:Pt:Head:Doc:CT
C0881954|Multisection^WO & W contrast Intravenous:Finding:Point in time:Internal auditory canal+Posterior fossa:Document:MRI
C0881954|Internal auditory canal and Posterior fossa MRI WO and W contrast IV
C0881954|Multisection^WO & W contrast IV:Find:Pt:Internal auditory canal+Posterior fossa:Doc:MRI
C0881954|IAC+Post fossa MRI WO+W contr IV
C0881994|Abd XR AP+Lat
C0881994|Abdomen X-ray AP and lateral
C0881994|Views AP & lateral:Find:Pt:Abdomen:Doc:XR
C0881994|Views AP & lateral:Finding:Point in time:Abdomen:Document:XR
C1114488|Pituitary+ST MRI WO contr
C1114488|Pituitary and Sella turcica MRI WO contrast
C1114488|Multisection^WO contrast:Finding:Point in time:Pituitary+Sella turcica:Document:MRI
C1114488|Multisection^WO contrast:Find:Pt:Pituitary+Sella turcica:Doc:MRI
C1114934|Hip MRI WO and W contrast IV
C1114934|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip:Document:MRI
C1114934|Hip MRI WO+W contr IV
C1114934|Multisection^WO & W contrast IV:Find:Pt:Hip:Doc:MRI
C1116466|Unspecified body region US during surgery
C1116466|XXX US in Surg
C1116466|Multisection^during surgery:Find:Pt:XXX:Doc:US
C1116466|Multisection^during surgery:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C1114531|T+L-spine XR Scoli stand
C1114531|Spine Thoracic and Lumbar X-ray scoliosis standing
C1114531|Views scoliosis^standing:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1114531|Views scoliosis^standing:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1114545|R & L-oblique views:Find:Pt:Chest:Nar:XR
C1114545|Deprecated Chest XR R & L-oblique
C1114545|Deprecated Chest X-ray R-oblique & L-oblique upright
C1114545|R & L-oblique views:Finding:Point in time:Chest:Narrative:XR
C1114585|Finger second X-ray
C1114585|Finger.2nd XR
C1114585|Views:Find:Pt:Finger.second:Doc:XR
C1114585|Views:Finding:Point in time:Finger.second:Document:XR
C1114586|Finger.3rd XR
C1114586|Finger third X-ray
C1114586|Views:Find:Pt:Finger.third:Doc:XR
C1114586|Views:Finding:Point in time:Finger.third:Document:XR
C1114592|Joint X-ray Single view
C1114592|Joint XR 1V
C1114592|View 1:Finding:Point in time:Joint:Document:XR
C1114592|View 1:Find:Pt:Joint:Doc:XR
C1114601|Elbow MRI WO contr
C1114601|Elbow MRI WO contrast
C1114601|Multisection^WO contrast:Finding:Point in time:Elbow:Document:MRI
C1114601|Multisection^WO contrast:Find:Pt:Elbow:Doc:MRI
C1114947|Head CT WO contrast
C1114947|Head CT WO contr
C1114947|Multisection^WO contrast:Finding:Point in time:Head:Document:Computerized Tomography
C1114947|Multisection^WO contrast:Find:Pt:Head:Doc:CT
C1114612|Lacrimal duct Fluoroscopy W contrast intra lacrimal duct
C1114612|Lacrimal duct Flr W contr intra LD
C1114612|Views^W contrast intra lacrimal duct:Find:Pt:Lacrimal duct:Doc:XR.fluor
C1114612|Views^W contrast intra lacrimal duct:Finding:Point in time:Lacrimal duct:Document:XR.fluor
C1114654|Multisection^WO & W contrast IV:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:MRI
C1114654|Spine Cervical and Thoracic and Lumbar MRI WO and W contrast IV
C1114654|C+T+L-spine MRI WO+W contr IV
C1114654|Multisection^WO & W contrast Intravenous:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:MRI
C1114671|Extremity veins MRI angiogram
C1114671|Extr vv MRI.Angio
C1114671|Multisection:Find:Pt:Extremity veins:Doc:MRI.angio
C1114671|Multisection:Finding:Point in time:Extremity veins:Document:MRI.angio
C1114458|Chest Fluoroscopy
C1114458|Chest Flr
C1114458|Views:Find:Pt:Chest:Doc:XR.fluor
C1114458|Views:Finding:Point in time:Chest:Document:XR.fluor
C1543434|Views^W contrast retrograde:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C1543434|Kidney - bilateral Fluoroscopy W contrast retrograde
C1543434|Views^W contrast retrograde:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C1543434|Kdny-Bl Flr W contr retro
C1543736|RI WB W Ga-67 IV
C1543736|Views whole body^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543736|Views whole body^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543736|Scan whole body W Ga-67 IV
C1543738|RI for Abscess W Ga-67 IV
C1543738|Views for abscess^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543738|Views for abscess^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543738|Scan for abscess W Ga-67 IV
C1543783|Hrt RI PF W ADE+Tc99mMIBI IV
C1543783|Heart Scan perfusion W adenosine and W Tc-99m Sestamibi IV
C1543783|Views perfusion^W adenosine & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc
C1543783|Views perfusion^W adenosine & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542976|Spleen RI W RNC Heat Damaged RBC IV
C1542976|Spleen Scan W radionuclide tagged heat damaged RBC IV
C1542976|Views^W radionuclide tagged heat damaged RBC IV:Find:Pt:Spleen:Doc:Radnuc
C1542976|Views^W radionuclide tagged heat damaged RBC Intravenous:Finding:Point in time:Spleen:Document:Radnuc
C1543863|BM SPECT Ltd W RNC IV
C1543863|Bone marrow SPECT limited
C1543863|Multisection limited^W radionuclide IV:Find:Pt:Bone marrow:Doc:Radnuc.SPECT
C1543863|Multisection limited^W radionuclide Intravenous:Finding:Point in time:Bone marrow:Document:Radnuc.SPECT
C1543877|Parotid gland RI Flow W RNC IV
C1543877|Parotid gland Scan flow
C1543877|Views flow^W radionuclide Intravenous:Finding:Point in time:Parotid gland:Document:Radnuc
C1543877|Views flow^W radionuclide IV:Find:Pt:Parotid gland:Doc:Radnuc
C1543889|Brain RI Delayed Static W RNC IV
C1543889|Brain Scan delayed static
C1543889|Views delayed static^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc
C1543889|Views delayed static^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1542852|Hrt RI Gated+WM+EF W RNC IV
C1542852|Heart Scan gated and wall motion and ejection fraction
C1542852|Views gated & wall motion & ejection fraction^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1542852|Views gated & wall motion & ejection fraction^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1542856|RI Mul Areas W Ga-67 IV
C1542856|Views multiple areas^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1542856|Views multiple areas^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1542856|Scan multiple areas W Ga-67 IV
C1543519|Lower extremity vein - right US.doppler
C1543519|LE v-R DOP
C1543519|Multisection:Finding:Point in time:Lower extremity vein.right:Document:Ultrasound.doppler
C1543519|Multisection:Find:Pt:Lower extremity vein.right:Doc:US.doppler
C1543175|Brst.duct Mam W contr intra Dct
C1543175|Breast duct Mammogram W contrast intra duct
C1543175|Views^W contrast intra duct:Find:Pt:Breast.duct:Doc:Mam
C1543175|Views^W contrast intra duct:Finding:Point in time:Breast.duct:Document:Mam
C1543219|Carotid artery.cervical - bilateral Fluoroscopic angiogram W contrast IA
C1543219|Carot a.cervical-Bl XRA W contr IA
C1543219|Views^W contrast IA:Find:Pt:Carotid artery.cervical.bilateral:Doc:XR.fluor.angio
C1543219|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.cervical.bilateral:Document:XR.fluor.angio
C1525162|Kidney Transplant US Bx guid
C1525162|US Guidance for biopsy of Kidney transplant
C1525162|Guidance for biopsy:Find:Pt:Kidney transplant:Doc:US
C1525162|Guidance for biopsy:Finding:Point in time:Kidney transplant:Document:Ultrasound
C1543268|Brst.duct-R Mam W contr intra Dcts
C1543268|Breast duct - right Mammogram W contrast intra multiple ducts
C1543268|Views^W contrast intra multiple ducts:Finding:Point in time:Breast.duct.right:Document:Mam
C1543268|Views^W contrast intra multiple ducts:Find:Pt:Breast.duct.right:Doc:Mam
C1543723|Hrt RI Rest+W DBM+RNC IV
C1543723|Heart Scan at rest and W dobutamine and W radionuclide IV
C1543723|Views^at rest & W dobutamine & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543723|Views^at rest & W dobutamine & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1526796|Ankle - left X-ray 2 views W manual stress
C1526796|Ankle-L XR 2V W Stress
C1526796|Views 2^W manual stress:Finding:Point in time:Ankle.left:Document:XR
C1526796|Views 2^W manual stress:Find:Pt:Ankle.left:Doc:XR
C1524851|Foot CT WO contrast
C1524851|Ft CT WO contr
C1524851|Multisection^WO contrast:Find:Pt:Foot:Doc:CT
C1524851|Multisection^WO contrast:Finding:Point in time:Foot:Document:Computerized Tomography
C1525173|Upper extremity vessels - left MRI angiogram
C1525173|UE ves-L MRI.Angio
C1525173|Multisection:Finding:Point in time:Upper extremity vessels.left:Document:MRI.angio
C1525173|Multisection:Find:Pt:Upper extremity vessels.left:Doc:MRI.angio
C1524439|Upper extremity vessels MRI angiogram
C1524439|UE ves MRI.Angio
C1524439|Multisection:Finding:Point in time:Upper extremity vessels:Document:MRI.angio
C1524439|Multisection:Find:Pt:Upper extremity vessels:Doc:MRI.angio
C1524442|Head CT limited
C1524442|Head CT Ltd
C1524442|Multisection limited:Finding:Point in time:Head:Document:Computerized Tomography
C1524442|Multisection limited:Find:Pt:Head:Doc:CT
C3853707|Orbit MRI WO+W contr IV
C3853707|Multisection^WO & W contrast IV:Find:Pt:Orbit:Doc:MRI
C3853707|Orbit MRI WO and W contrast IV
C3853707|Multisection^WO & W contrast Intravenous:Finding:Point in time:Orbit:Document:MRI
C1525227|Neck vv MRI.Angio WO+W contr IV
C1525227|Neck veins MRI angiogram WO and W contrast IV
C1525227|Multisection^WO & W contrast Intravenous:Finding:Point in time:Neck veins:Document:MRI.angio
C1525227|Multisection^WO & W contrast IV:Find:Pt:Neck veins:Doc:MRI.angio
C1525339|Ankle XR Mortise
C1525339|Ankle X-ray Mortise
C1525339|View Mortise:Find:Pt:Ankle:Doc:XR
C1525339|View Mortise:Finding:Point in time:Ankle:Document:XR
C1524681|Should-L XR Outlet
C1524681|Shoulder - left X-ray outlet
C1524681|View outlet:Find:Pt:Shoulder.left:Doc:XR
C1524681|View outlet:Finding:Point in time:Shoulder.left:Document:XR
C1525347|Should-L XR Stryker Notch
C1525347|Shoulder - left X-ray Stryker Notch
C1525347|View Stryker Notch:Finding:Point in time:Shoulder.left:Document:XR
C1525347|View Stryker Notch:Find:Pt:Shoulder.left:Doc:XR
C1525514|Knee-L XR AP+Lat+Tunnel
C1525514|Knee - left X-ray AP and lateral and tunnel
C1525514|Views AP & lateral & tunnel:Find:Pt:Knee.left:Doc:XR
C1525514|Views AP & lateral & tunnel:Finding:Point in time:Knee.left:Document:XR
C1525515|Knee XR AP+Lat+Obl+Tunnel
C1525515|Knee X-ray AP and lateral and oblique and tunnel
C1525515|Views AP & lateral & oblique & tunnel:Find:Pt:Knee:Doc:XR
C1525515|Views AP & lateral & oblique & tunnel:Finding:Point in time:Knee:Document:XR
C1525533|Ankle-Bl XR Lat+Mortise
C1525533|Ankle - bilateral X-ray lateral and Mortise
C1525533|Views lateral & Mortise:Finding:Point in time:Ankle.bilateral:Document:XR
C1525533|Views lateral & Mortise:Find:Pt:Ankle.bilateral:Doc:XR
C1525583|Elbow Flr W contr IS
C1525583|Elbow Fluoroscopy W contrast IS
C1525583|Views^W contrast IS:Find:Pt:Elbow:Doc:XR.fluor
C1525583|Views^W contrast Intrasynovial:Finding:Point in time:Elbow:Document:XR.fluor
C1525591|Cerebral v XRA W contr IV
C1525591|Cerebral vein Fluoroscopic angiogram W contrast IV
C1525591|Views^W contrast Intravenous:Finding:Point in time:Cerebral vein:Document:XR.fluor.angio
C1525591|Views^W contrast IV:Find:Pt:Cerebral vein:Doc:XR.fluor.angio
C1525604|L-spine XR stand
C1525604|Views^standing:Find:Pt:Spine.lumbar:Doc:XR
C1525604|Views^standing:Finding:Point in time:Spine.lumbar:Document:XR
C1525604|Lumbar spine X-ray standing
C1525611|Brain+Larynx MRI W contr IV
C1525611|Brain and Larynx MRI W contrast IV
C1525611|Multisection^W contrast IV:Find:Pt:Brain+Larynx:Doc:MRI
C1525611|Multisection^W contrast Intravenous:Finding:Point in time:Brain+Larynx:Document:MRI
C1525623|TMJ-Bl MRI
C1525623|Temporomandibular joint - bilateral MRI
C1525623|Multisection:Finding:Point in time:Temporomandibular joint.bilateral:Document:MRI
C1525623|Multisection:Find:Pt:Temporomandibular joint.bilateral:Doc:MRI
C1525656|TMJ-L MRI WO+W contr IV
C1525656|Multisection^WO & W contrast IV:Find:Pt:Temporomandibular joint.left:Doc:MRI
C1525656|Temporomandibular joint - left MRI WO and W contrast IV
C1525656|Multisection^WO & W contrast Intravenous:Finding:Point in time:Temporomandibular joint.left:Document:MRI
C1525711|Ac arch+VA-L XRA W contr IA
C1525711|Aortic arch and Vertebral artery - left Fluoroscopic angiogram W contrast IA
C1525711|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Vertebral artery.left:Document:XR.fluor.angio
C1525711|Views^W contrast IA:Find:Pt:Aortic arch+Vertebral artery.left:Doc:XR.fluor.angio
C1525724|Gastric artery - left Fluoroscopic angiogram W contrast IA
C1525724|Gastric a-L XRA W contr IA
C1525724|Views^W contrast IA:Find:Pt:Gastric artery.left:Doc:XR.fluor.angio
C1525724|Views^W contrast Intra-arterial:Finding:Point in time:Gastric artery.left:Document:XR.fluor.angio
C1525729|Pudendal artery.internal Fluoroscopic angiogram W contrast IA
C1525729|IPA XRA W contr IA
C1525729|Views^W contrast IA:Find:Pt:Pudendal artery.internal:Doc:XR.fluor.angio
C1525729|Views^W contrast Intra-arterial:Finding:Point in time:Pudendal artery.internal:Document:XR.fluor.angio
C1525850|Brst-Bl Mam Mag+Spot
C1525850|Breast - bilateral Mammogram magnification and spot
C1525850|Views magnification & spot:Find:Pt:Breast.bilateral:Doc:Mam
C1525850|Views magnification & spot:Finding:Point in time:Breast.bilateral:Document:Mam
C1525859|Thumb-Bl XR W Stress
C1525859|Thumb - bilateral X-ray W manual stress
C1525859|Views^W manual stress:Finding:Point in time:Thumb.bilateral:Document:XR
C1525859|Views^W manual stress:Find:Pt:Thumb.bilateral:Doc:XR
C1524135|Ac arch+Carot a.ext-L XRA W contr IA
C1524135|Aortic arch and Carotid artery.external - left Fluoroscopic angiogram W contrast IA
C1524135|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery.external.left:Document:XR.fluor.angio
C1524135|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery.external.left:Doc:XR.fluor.angio
C1525886|Adrenal v-L XRA W contr IV
C1525886|Views^W contrast IV:Find:Pt:Adrenal vein.left:Doc:XR.fluor.angio
C1525886|Adrenal vein - left Fluoroscopic angiogram W contrast IV
C1525886|Views^W contrast Intravenous:Finding:Point in time:Adrenal vein.left:Document:XR.fluor.angio
C1525814|Cervical Spine vessels MRI angiogram WO contrast
C1525814|C-spine ves MRI.Angio WO contr
C1525814|Multisection^WO contrast:Find:Pt:Spine.cervical vessels:Doc:MRI.angio
C1525814|Multisection^WO contrast:Finding:Point in time:Spine.cervical vessels:Document:MRI.angio
C1526109|Should-R XR Outlet+Y
C1526109|Shoulder - right X-ray outlet and Y
C1526109|Views outlet & Y:Finding:Point in time:Shoulder.right:Document:XR
C1526109|Views outlet & Y:Find:Pt:Shoulder.right:Doc:XR
C1526119|Thumb - right X-ray W manual stress
C1526119|Thumb-R XR W Stress
C1526119|Views^W manual stress:Find:Pt:Thumb.right:Doc:XR
C1526119|Views^W manual stress:Finding:Point in time:Thumb.right:Document:XR
C1526135|Should XR Garth
C1526135|Shoulder X-ray Garth
C1526135|View Garth:Finding:Point in time:Shoulder:Document:XR
C1526135|View Garth:Find:Pt:Shoulder:Doc:XR
C1526165|View 1 limited:Find:Pt:Skull:Nar:XR
C1526165|Deprecated Skull X-ray View
C1526165|Deprecated Skull XR 1V Ltd
C1526165|View 1 limited:Finding:Point in time:Skull:Narrative:XR
C1526206|Periph ves XRA W contr
C1526206|Peripheral vessels Fluoroscopic angiogram W contrast
C1526206|Views^W contrast:Find:Pt:Peripheral vessels:Doc:XR.fluor.angio
C1526206|Views^W contrast:Finding:Point in time:Peripheral vessels:Document:XR.fluor.angio
C1524474|Multisection^W contrast Intrasynovial:Finding:Point in time:Shoulder.left:Document:MRI
C1524474|Multisection^W contrast IS:Find:Pt:Shoulder.left:Doc:MRI
C1524474|Shoulder - left MRI W contrast IS
C1524474|Should-L MRI W contr IS
C1524487|Multisection^W contrast IV:Find:Pt:Abdomen>Aorta.abdominal:Doc:CT
C1524487|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen>Aorta.abdominal:Document:Computerized Tomography
C1524487|Abdominal Aorta CT W contrast IV
C1524487|Abd Aorta CT W contr IV
C1524871|Hip - bilateral MRI WO contrast
C1524871|Hip-Bl MRI WO contr
C1524871|Multisection^WO contrast:Find:Pt:Hip.bilateral:Doc:MRI
C1524871|Multisection^WO contrast:Finding:Point in time:Hip.bilateral:Document:MRI
C1524877|Upper arm - left CT WO contrast
C1524877|Upper arm-L CT WO contr
C1524877|Multisection^WO contrast:Find:Pt:Upper arm.left:Doc:CT
C1524877|Multisection^WO contrast:Finding:Point in time:Upper arm.left:Document:Computerized Tomography
C1524531|Forearm-L CT W contr IV
C1524531|Forearm - left CT W contrast IV
C1524531|Multisection^W contrast Intravenous:Finding:Point in time:Forearm.left:Document:Computerized Tomography
C1524531|Multisection^W contrast IV:Find:Pt:Forearm.left:Doc:CT
C1524895|Knee-R MRI WO contr
C1524895|Knee - right MRI WO contrast
C1524895|Multisection^WO contrast:Finding:Point in time:Knee.right:Document:MRI
C1524895|Multisection^WO contrast:Find:Pt:Knee.right:Doc:MRI
C1524929|Clavicle X-ray Single view
C1524929|Clavicle XR 1V
C1524929|View 1:Find:Pt:Clavicle:Doc:XR
C1524929|View 1:Finding:Point in time:Clavicle:Document:XR
C1524945|Finger.3rd XR Lat
C1524945|Finger third X-ray lateral
C1524945|View lateral:Finding:Point in time:Finger.third:Document:XR
C1524945|View lateral:Find:Pt:Finger.third:Doc:XR
C1524947|Hand XR Lat
C1524947|Hand X-ray lateral
C1524947|View lateral:Finding:Point in time:Hand:Document:XR
C1524947|View lateral:Find:Pt:Hand:Doc:XR
C1524293|Fluoroscopy Guidance for biopsy of Chest
C1524293|Chest Flr Bx guid
C1524293|Guidance for biopsy:Find:Pt:Chest:Doc:XR.fluor
C1524293|Guidance for biopsy:Finding:Point in time:Chest:Document:XR.fluor
C1524294|Chest CT Bx guid
C1524294|CT Guidance for biopsy of Chest
C1524294|Guidance for biopsy:Finding:Point in time:Chest:Document:Computerized Tomography
C1524294|Guidance for biopsy:Find:Pt:Chest:Doc:CT
C1524305|T-spine CT Bx guid
C1524305|Guidance for biopsy:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C1524305|Guidance for biopsy:Find:Pt:Spine.thoracic:Doc:CT
C1524305|CT Guidance for biopsy of Thoracic spine
C1524954|Knee - left X-ray lateral
C1524954|Knee-L XR Lat
C1524954|View lateral:Find:Pt:Knee.left:Doc:XR
C1524954|View lateral:Finding:Point in time:Knee.left:Document:XR
C1524973|Brst Mam
C1524973|Breast Mammogram
C1524973|Views:Find:Pt:Breast:Doc:Mam
C1524973|Views:Finding:Point in time:Breast:Document:Mam
C1524348|Face MRI
C1524348|Multisection:Find:Pt:Face:Doc:MRI
C1524348|Multisection:Finding:Point in time:Face:Document:MRI
C1525005|Scapula - left X-ray 2 views
C1525005|Scapula-L XR 2V
C1525005|Views 2:Finding:Point in time:Scapula.left:Document:XR
C1525005|Views 2:Find:Pt:Scapula.left:Doc:XR
C1525008|C-spine XR 2V
C1525008|Views 2:Find:Pt:Spine.cervical:Doc:XR
C1525008|Views 2:Finding:Point in time:Spine.cervical:Document:XR
C1525008|Cervical spine X-ray 2 views
C1524668|Ft-Bl MRI WO+W contr IV
C1524668|Multisection^WO & W contrast Intravenous:Finding:Point in time:Foot.bilateral:Document:MRI
C1524668|Multisection^WO & W contrast IV:Find:Pt:Foot.bilateral:Doc:MRI
C1524668|Foot - bilateral MRI WO and W contrast IV
C1524750|Multisection^WO & W contrast IV:Find:Pt:Hip.right:Doc:CT
C1524750|Hip-R CT WO+W contr IV
C1524750|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip.right:Document:Computerized Tomography
C1524750|Hip - right CT WO and W contrast IV
C1525037|Radius+Ulna XR AP+Lat
C1525037|Radius and Ulna X-ray AP and lateral
C1525037|Views AP & lateral:Finding:Point in time:Radius+Ulna:Document:XR
C1525037|Views AP & lateral:Find:Pt:Radius+Ulna:Doc:XR
C1524412|Upper arm CT
C1524412|Multisection:Find:Pt:Upper arm:Doc:CT
C1524412|Multisection:Finding:Point in time:Upper arm:Document:Computerized Tomography
C1524781|Should-L CT WO+W contr IV
C1524781|Multisection^WO & W contrast Intravenous:Finding:Point in time:Shoulder.left:Document:Computerized Tomography
C1524781|Shoulder - left CT WO and W contrast IV
C1524781|Multisection^WO & W contrast IV:Find:Pt:Shoulder.left:Doc:CT
C1524791|Multisection^WO & W contrast IV:Find:Pt:Scrotum+Testicle:Doc:MRI
C1524791|Multisection^WO & W contrast Intravenous:Finding:Point in time:Scrotum+Testicle:Document:MRI
C1524791|Scrotum and Testicle MRI WO and W contrast IV
C1524791|Scrotum+Test MRI WO+W contr IV
C1525066|Finger-L XR AP+Lat+Obl
C1525066|Finger - left X-ray AP and lateral and oblique
C1525066|Views AP & lateral & oblique:Finding:Point in time:Finger.left:Document:XR
C1525066|Views AP & lateral & oblique:Find:Pt:Finger.left:Doc:XR
C1525071|Radius+Ulna-L XR Obl
C1525071|Radius - left and Ulna.left X-ray oblique
C1525071|Views oblique:Finding:Point in time:Radius.left+Ulna.left:Document:XR
C1525071|Views oblique:Find:Pt:Radius.left+Ulna.left:Doc:XR
C1525095|CT Guidance for biopsy of Adrenal gland
C1525095|Adrenal CT Bx guid
C1525095|Guidance for biopsy:Finding:Point in time:Abdomen>Adrenal gland:Document:Computerized Tomography
C1525095|Guidance for biopsy:Find:Pt:Abdomen>Adrenal gland:Doc:CT
C1525096|CT Guidance for biopsy of Muscle
C1525096|Muscle CT Bx guid
C1525096|Guidance for biopsy:Find:Pt:Muscle:Doc:CT
C1525096|Guidance for biopsy:Finding:Point in time:Muscle:Document:Computerized Tomography
C1830182|XXX CT Asp or Inj of Cyst guid
C1830182|CT Guidance for aspiration or injection of cyst of Unspecified body region
C1830182|Guidance for aspiration or injection of cyst:Find:Pt:XXX:Doc:CT
C1830182|Guidance for aspiration or injection of cyst:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1830238|Brst-R Mam 1V
C1830238|Breast - right Mammogram Single view
C1830238|View 1:Find:Pt:Breast.right:Doc:Mam
C1830238|View 1:Finding:Point in time:Breast.right:Document:Mam
C1831073|Knee - right X-ray 1 or 2 views
C1831073|Knee-R XR 1V or 2V
C1831073|Views 1 or 2:Find:Pt:Knee.right:Doc:XR
C1831073|Views 1 or 2:Finding:Point in time:Knee.right:Document:XR
C1715403|Renal ves MRI.Angio WO contr
C1715403|Renal vessels MRI angiogram WO contrast
C1715403|Multisection^WO contrast:Find:Pt:Renal vessels:Doc:MRI.angio
C1715403|Multisection^WO contrast:Finding:Point in time:Renal vessels:Document:MRI.angio
C1715412|Hrt RI W Tc99mRBC IV
C1715412|Heart Scan W Tc-99m tagged RBC IV
C1715412|Views^W Tc-99m tagged RBC IV:Find:Pt:Heart:Doc:Radnuc
C1715412|Views^W Tc-99m tagged RBC Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1715421|Kidney SPECT W Tc99mGHA IV
C1715421|Kidney SPECT W Tc-99m glucoheptonate IV
C1715421|Multisection^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Kidney:Document:Radnuc.SPECT
C1715421|Multisection^W Tc-99m glucoheptonate IV:Find:Pt:Kidney:Doc:Radnuc.SPECT
C1715423|Liver US Ablation guid
C1715423|US Guidance for ablation of tissue of Liver
C1715423|Guidance for ablation of tissue:Find:Pt:Liver:Doc:US
C1715423|Guidance for ablation of tissue:Finding:Point in time:Liver:Document:Ultrasound
C1715427|US Guidance for fine needle aspiration of Kidney
C1715427|Kidney US FNA Asp
C1715427|Guidance for aspiration.fine needle:Finding:Point in time:Kidney:Document:Ultrasound
C1715427|Guidance for aspiration.fine needle:Find:Pt:Kidney:Doc:US
C1715428|Brst US FNA Asp
C1715428|US Guidance for fine needle aspiration of Breast
C1715428|Guidance for aspiration.fine needle:Find:Pt:Breast:Doc:US
C1715428|Guidance for aspiration.fine needle:Finding:Point in time:Breast:Document:Ultrasound
C1715430|Head+Neck US
C1715430|Head and Neck US
C1715430|Multisection:Find:Pt:Head+Neck:Doc:US
C1715430|Multisection:Finding:Point in time:Head+Neck:Document:Ultrasound
C1715442|LE-Bl XR AP 1V stand
C1715442|Lower extremity - bilateral X-ray AP single view standing
C1715442|View AP^standing:Find:Pt:Lower extremity.bilateral:Doc:XR
C1715442|View AP^standing:Finding:Point in time:Lower extremity.bilateral:Document:XR
C1715450|Femur XR AP+Lat port
C1715450|Femur X-ray AP and lateral portable
C1715450|Views AP & lateral portable:Find:Pt:Femur:Doc:XR
C1715450|Views AP & lateral portable:Finding:Point in time:Femur:Document:XR
C1648948|Deprecated Views portable:Finding:Point in time:Tibia.left:Narrative:XR
C1648948|Deprecated Tib-L XR port
C1648948|Views portable:Find:Pt:Tibia.left:Nar:XR
C1648948|Views portable:Finding:Point in time:Tibia.left:Narrative:XR
C1648948|Deprecated Tibia Left X-ray Portable
C1626801|Wrist-R XR Scaphoid 1V
C1626801|Wrist - right X-ray scaphoid single view
C1626801|View scaphoid:Find:Pt:Wrist.right:Doc:XR
C1626801|View scaphoid:Finding:Point in time:Wrist.right:Document:XR
C1714789|Elbow-R MRI Dyn W contr IV
C1714789|Elbow - right MRI dynamic W contrast IV
C1714789|Multisection dynamic^W contrast IV:Find:Pt:Elbow.right:Doc:MRI
C1714789|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Elbow.right:Document:MRI
C1714793|Oropharynx MRI
C1714793|Multisection:Find:Pt:Oropharynx:Doc:MRI
C1714793|Multisection:Finding:Point in time:Oropharynx:Document:MRI
C1714799|Brst-L US Bx needle guid
C1714799|US Guidance for needle biopsy of Breast - left
C1714799|Guidance for biopsy.needle:Finding:Point in time:Breast.left:Document:Ultrasound
C1714799|Guidance for biopsy.needle:Find:Pt:Breast.left:Doc:US
C1705866|Finger third - right X-ray GE 3 views
C1705866|Finger.3rd-R XR GE 3V
C1705866|Finger third - right Narrative X-ray GE 3 views
C1705866|Views GE 3:Finding:Point in time:Finger.third.right:Document:XR
C1705866|Views GE 3:Find:Pt:Finger.third.right:Doc:XR
C1715031|Hrt RI PF Ql Rest+W RNC IV
C1715031|Heart Scan perfusion qualitative at rest and W radionuclide IV
C1715031|Views perfusion qualitative^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1715031|Views perfusion qualitative^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1714506|US Guidance for aspiration of Breast
C1714506|Brst US Asp guid
C1714506|Guidance for aspiration:Find:Pt:Breast:Doc:US
C1714506|Guidance for aspiration:Finding:Point in time:Breast:Document:Ultrasound
C1644169|Neck XR AP+Lat
C1644169|Neck X-ray AP and lateral
C1644169|Views AP & lateral:Finding:Point in time:Neck:Document:XR
C1644169|Views AP & lateral:Find:Pt:Neck:Doc:XR
C1630751|CT Guidance for needle biopsy of Abdomen
C1630751|Abd CT Bx needle guid
C1630751|Guidance for biopsy.needle:Find:Pt:Abdomen:Doc:CT
C1630751|Guidance for biopsy.needle:Finding:Point in time:Abdomen:Document:Computerized Tomography
C3484379|Thyroid MRI
C3484379|Multisection:Find:Pt:Thyroid:Doc:MRI
C3484379|Multisection:Finding:Point in time:Thyroid:Document:MRI
C1953939|Deprecated Heel-Bl XR 2V
C1953939|Views 2:Finding:Point in time:Calcaneus.bilateral:Document:XR
C1953939|Deprecated Calcaneus - bilateral X-ray 2 views
C1953939|Views 2:Find:Pt:Calcaneus.bilateral:Doc:XR
C1953954|Upper extremity artery US
C1953954|UE a US
C1953954|Multisection:Find:Pt:Upper extremity artery:Doc:US
C1953954|Multisection:Finding:Point in time:Upper extremity artery:Document:Ultrasound
C1953961|Multisection^WO & W contrast IV:Find:Pt:Clavicle.left:Doc:MRI
C1953961|Clavicle - left MRI WO and W contrast IV
C1953961|Multisection^WO & W contrast Intravenous:Finding:Point in time:Clavicle.left:Document:MRI
C1953961|Clavicle-L MRI WO+W contr IV
C1953964|Clavicle - right MRI WO contrast
C1953964|Clavicle-R MRI WO contr
C1953964|Multisection^WO contrast:Finding:Point in time:Clavicle.right:Document:MRI
C1953964|Multisection^WO contrast:Find:Pt:Clavicle.right:Doc:MRI
C2926621|Hrt CT
C2926621|Heart CT
C2926621|Multisection:Finding:Point in time:Chest>Heart:Document:Computerized Tomography
C2926621|Multisection:Find:Pt:Chest>Heart:Doc:CT
C2925709|AVF XRA W contr IV
C2925709|AV fistula Fluoroscopic angiogram W contrast IV
C2925709|Views^W contrast Intravenous:Finding:Point in time:AV fistula:Document:XR.fluor.angio
C2925709|Views^W contrast IV:Find:Pt:AV fistula:Doc:XR.fluor.angio
C3173522|Breast lymphatics - right Scan W radionuclide intra lymphatic
C3173522|Brst lymphr-R RI W RNC Intra Lymph
C3173522|Views^W radionuclide intra lymphatic:Finding:Point in time:Breast lymphatics.right:Document:Radnuc
C3173522|Views^W radionuclide intra lymphatic:Find:Pt:Breast lymphatics.right:Doc:Radnuc
C3533561|C-spine Flr FJ DN guid
C3533561|Guidance for facet joint denervation:Finding:Point in time:Spine.cervical:Document:XR.fluor
C3533561|Guidance for facet joint denervation:Find:Pt:Spine.cervical:Doc:XR.fluor
C3533561|Fluoroscopy Guidance for facet joint denervation of Cervical spine
C3533553|Guidance for removal of catheter^tunneled:Finding:Point in time:Central vein:Document:XR.fluor
C3533553|Fluoroscopy Guidance for removal of catheter from Central vein-- Tunneled
C3533553|Centl v Flr cath rem guid Tunneled
C3533553|Guidance for removal of catheter^tunneled:Find:Pt:Central vein:Doc:XR.fluor
C3533908|Multisection diagnostic:Find:Pt:Breast.right:Doc:Mam.FFD.tomosynthesis
C3533908|Breast - right FFD mammogram-tomosynthesis diagnostic
C3533908|Multisection diagnostic:Finding:Point in time:Breast.right:Document:Mam.FFD.tomosynthesis
C3533908|Brst-R FFDM-DBT Dx
C3533907|Brst-L FFDM-DBT Dx
C3533907|Breast - left FFD mammogram-tomosynthesis diagnostic
C3533907|Multisection diagnostic:Find:Pt:Breast.left:Doc:Mam.FFD.tomosynthesis
C3533907|Multisection diagnostic:Finding:Point in time:Breast.left:Document:Mam.FFD.tomosynthesis
C3262933|Multisection^W contrast Intrasynovial:Finding:Point in time:Elbow.right:Document:Computerized Tomography
C3262933|Elbow - right CT W contrast IS
C3262933|Elbow-R CT W contr IS
C3262933|Multisection^W contrast IS:Find:Pt:Elbow.right:Doc:CT
C3262945|Guidance for drainage of abscess:Finding:Point in time:Pancreas:Document:XR.fluor
C3262945|Guidance for drainage of abscess:Find:Pt:Pancreas:Doc:XR.fluor
C3262945|Fluoroscopy Guidance for drainage of abscess of Pancreas
C3262945|Pancreas Flr Abscess drain guid
C3262963|Knee - left X-ray 2 views and tunnel standing
C3262963|Knee-L XR 2V+Tunnel stand
C3262963|Views 2 & tunnel^standing:Finding:Point in time:Knee.left:Document:XR
C3262963|Views 2 & tunnel^standing:Find:Pt:Knee.left:Doc:XR
C3262994|Multisection^WO & W contrast Intravenous:Finding:Point in time:Forearm.bilateral:Document:MRI
C3262994|Forearm - bilateral MRI WO and W contrast IV
C3262994|Multisection^WO & W contrast IV:Find:Pt:Forearm.bilateral:Doc:MRI
C3262994|Forearm-Bl MRI WO+W contr IV
C3263001|Multisection^WO & W contrast IV:Find:Pt:Upper arm.bilateral:Doc:MRI
C3263001|Upper arm-Bl MRI WO+W contr IV
C3263001|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper arm.bilateral:Document:MRI
C3263001|Upper arm - bilateral MRI WO and W contrast IV
C3482447|T-spine XR 1V port
C3482447|View 1 portable:Find:Pt:Spine.thoracic:Doc:XR
C3482447|View 1 portable:Finding:Point in time:Spine.thoracic:Document:XR
C3482447|Thoracic spine X-ray Single view portable
C3263023|Lower Extremity Joint MRI W contrast IS
C3263023|Multisection^W contrast Intrasynovial:Finding:Point in time:Lower extremity.joint:Document:MRI
C3263023|LE.joint MRI W contr IS
C3263023|Multisection^W contrast IS:Find:Pt:Lower extremity.joint:Doc:MRI
C3263067|Ankle - right X-ray 3 views standing
C3263067|Ankle-R XR 3V stand
C3263067|Views 3^standing:Finding:Point in time:Ankle.right:Document:XR
C3263067|Views 3^standing:Find:Pt:Ankle.right:Doc:XR
C3263108|Elbow - left X-ray Single view
C3263108|Elbow-L XR 1V
C3263108|View 1:Find:Pt:Elbow.left:Doc:XR
C3263108|View 1:Finding:Point in time:Elbow.left:Document:XR
C3263213|Spinal cord US Bx guid
C3263213|US Guidance for biopsy of Spinal cord
C3263213|Guidance for biopsy:Finding:Point in time:Spinal cord:Document:Ultrasound
C3263213|Guidance for biopsy:Find:Pt:Spinal cord:Doc:US
C3262904|C-spine XR 5V+Swimmers
C3262904|Views 5 & Swimmers:Find:Pt:Spine.cervical:Doc:XR
C3262904|Views 5 & Swimmers:Finding:Point in time:Spine.cervical:Document:XR
C3262904|Cervical spine X-ray 5 views and Swimmers
C3262916|Pelvis CT Bx guid W contr IV
C3262916|CT Guidance for biopsy of Pelvis-- W contrast IV
C3262916|Guidance for biopsy^W contrast Intravenous:Finding:Point in time:Pelvis:Document:Computerized Tomography
C3262916|Guidance for biopsy^W contrast IV:Find:Pt:Pelvis:Doc:CT
C0945315|Deprecated DEXA
C0945315|Views:Find:Pt:Radius+Ulna.bilateral:Nar:XR.DEXA
C0945315|Views:Finding:Point in time:Radius+Ulna.bilateral:Narrative:XR.DEXA
C0945315|Deprecated Radius & Ulna bilateral DEXA Bone density
C0942203|Knee-Bl MRI WO+W contr IV
C0942203|Multisection^WO & W contrast IV:Find:Pt:Knee.bilateral:Doc:MRI
C0942203|Knee - bilateral MRI WO and W contrast IV
C0942203|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee.bilateral:Document:MRI
C0942231|Extremity - right US
C0942231|Extr-R US
C0942231|Multisection:Find:Pt:Extremity.right:Doc:US
C0942231|Multisection:Finding:Point in time:Extremity.right:Document:Ultrasound
C0942240|Foot - bilateral MRI
C0942240|Ft-Bl MRI
C0942240|Multisection:Find:Pt:Foot.bilateral:Doc:MRI
C0942240|Multisection:Finding:Point in time:Foot.bilateral:Document:MRI
C0942250|IAC-R XRTomo
C0942250|Internal auditory canal - right X-ray tomograph
C0942250|Multisection:Find:Pt:Internal auditory canal.right:Doc:XR.tomo
C0942250|Multisection:Finding:Point in time:Internal auditory canal.right:Document:XR.tomo
C0942256|Pelvis+Hip-R MRI
C0942256|Pelvis and Hip - right MRI
C0942256|Multisection:Find:Pt:Pelvis+Hip.right:Doc:MRI
C0942256|Multisection:Finding:Point in time:Pelvis+Hip.right:Document:MRI
C0942289|Vein-L XRA Atherect guid W contr IV
C0942289|Fluoroscopic angiogram Guidance for atherectomy of Vein - left-- W contrast IV
C0942289|Guidance for atherectomy^W contrast IV:Find:Pt:Vein.left:Doc:XR.fluor.angio
C0942289|Guidance for atherectomy^W contrast Intravenous:Finding:Point in time:Vein.left:Document:XR.fluor.angio
C0942331|Brst-L Mam Dx
C0942331|Breast - left Mammogram diagnostic
C0942331|Views diagnostic:Find:Pt:Breast.left:Doc:Mam
C0942331|Views diagnostic:Finding:Point in time:Breast.left:Document:Mam
C0942337|Hand-Bl XR Arthritis
C0942337|Hand - bilateral X-ray arthritis
C0942337|View arthritis:Finding:Point in time:Hand.bilateral:Document:XR
C0942337|View arthritis:Find:Pt:Hand.bilateral:Doc:XR
C0942351|Iliac a-L XRA Angpsty W contr IA
C0942351|Iliac artery - left Fluoroscopic angiogram Angioplasty W contrast IA
C0942351|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Iliac artery.left:Document:XR.fluor.angio
C0942351|Angioplasty^W contrast IA:Find:Pt:Iliac artery.left:Doc:XR.fluor.angio
C0942354|Tibl a-L XRA Angpsty W contr IA
C0942354|Tibial artery - left Fluoroscopic angiogram Angioplasty W contrast IA
C0942354|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibial artery.left:Document:XR.fluor.angio
C0942354|Angioplasty^W contrast IA:Find:Pt:Tibial artery.left:Doc:XR.fluor.angio
C0942356|Administration of vasodilator into catheter of Vein - left
C0942356|Vein-L VD admin into cath
C0942356|Administration of vasodilator into catheter:Find:Pt:Vein.left:Doc
C0942356|Administration of vasodilator into catheter:Finding:Point in time:Vein.left:Document
C0942368|Hand-R XR 2V
C0942368|Hand - right X-ray 2 views
C0942368|Views 2:Find:Pt:Hand.right:Doc:XR
C0942368|Views 2:Finding:Point in time:Hand.right:Document:XR
C0882038|Neck ves MRI.Angio W contr IV
C0882038|Neck vessels MRI angiogram W contrast IV
C0882038|Multisection^W contrast IV:Find:Pt:Neck vessels:Doc:MRI.angio
C0882038|Multisection^W contrast Intravenous:Finding:Point in time:Neck vessels:Document:MRI.angio
C0882054|Iliac artery Internal Fluoroscopic angiogram W contrast IA
C0882054|Iliac a.Int XRA W contr IA
C0882054|Views^W contrast IA:Find:Pt:Iliac artery.internal:Doc:XR.fluor.angio
C0882054|Views^W contrast Intra-arterial:Finding:Point in time:Iliac artery.internal:Document:XR.fluor.angio
C0882055|Pelvis CT Asp guid
C0882055|CT Guidance for aspiration of Pelvis
C0882055|Guidance for aspiration:Finding:Point in time:Pelvis:Document:Computerized Tomography
C0882055|Guidance for aspiration:Find:Pt:Pelvis:Doc:CT
C0882056|CT Guidance for biopsy of Pelvis
C0882056|Pelvis CT Bx guid
C0882056|Guidance for biopsy:Find:Pt:Pelvis:Doc:CT
C0882056|Guidance for biopsy:Finding:Point in time:Pelvis:Document:Computerized Tomography
C0882174|Urinary bladder Scan
C0882174|Bladder RI W RNC IV
C0882174|Views^W radionuclide Intravenous:Finding:Point in time:Urinary bladder:Document:Radnuc
C0882174|Views^W radionuclide IV:Find:Pt:Urinary bladder:Doc:Radnuc
C0882175|Urinary bladder US
C0882175|Bladder US
C0882175|Multisection:Find:Pt:Urinary bladder:Doc:US
C0882175|Multisection:Finding:Point in time:Urinary bladder:Document:Ultrasound
C0882200|CT Guidance for biopsy of Unspecified body region
C0882200|XXX CT Bx guid
C0882200|Guidance for biopsy:Find:Pt:XXX:Doc:CT
C0882200|Guidance for biopsy:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C0884113|Vessel Fluoroscopic angiogram Single view W contrast IA
C0884113|View 1^W contrast IA:Find:Pt:Vessel:Doc:XR.fluor.angio
C0884113|View 1^W contrast Intra-arterial:Finding:Point in time:Vessel:Document:XR.fluor.angio
C0884113|Vesl XRA 1V W contr IA
C0882224|Hepatic artery Fluoroscopic angiogram W contrast IA
C0882224|Hep a XRA W contr IA
C0882224|Views^W contrast Intra-arterial:Finding:Point in time:Hepatic artery:Document:XR.fluor.angio
C0882224|Views^W contrast IA:Find:Pt:Hepatic artery:Doc:XR.fluor.angio
C0942088|Vein-Bl XRA W contr IV
C0942088|Vein - bilateral Fluoroscopic angiogram W contrast IV
C0942088|Views^W contrast IV:Find:Pt:Vein.bilateral:Doc:XR.fluor.angio
C0942088|Views^W contrast Intravenous:Finding:Point in time:Vein.bilateral:Document:XR.fluor.angio
C0945306|Knee-Bl Flr W contr IS
C0945306|Views^W contrast IS:Find:Pt:Knee.bilateral:Doc:XR.fluor
C0945306|Views^W contrast Intrasynovial:Finding:Point in time:Knee.bilateral:Document:XR.fluor
C0945306|Knee - bilateral Fluoroscopy W contrast IS
C0942125|Views:Find:Pt:Carpal bones.right:Nar:XR
C0942125|Views:Finding:Point in time:Carpal bones.right:Narrative:XR
C0942125|Deprecated Carpal bones-R XR
C0942125|Deprecated Carpal bones - right X-ray
C0881784|TA CT
C0881784|Multisection:Find:Pt:Chest>Aorta.thoracic:Doc:CT
C0881784|Multisection:Finding:Point in time:Chest>Aorta.thoracic:Document:Computerized Tomography
C0881784|Thoracic Aorta CT
C0881853|XXX Flr PC drain guid
C0881853|Fluoroscopy Guidance for percutaneous drainage of Unspecified body region
C0881853|Guidance for percutaneous drainage:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C0881853|Guidance for percutaneous drainage:Find:Pt:XXX:Doc:XR.fluor
C0881854|Celiac a XRA W contr IA
C0881854|Celiac artery Fluoroscopic angiogram W contrast IA
C0881854|Views^W contrast IA:Find:Pt:Celiac artery:Doc:XR.fluor.angio
C0881854|Views^W contrast Intra-arterial:Finding:Point in time:Celiac artery:Document:XR.fluor.angio
C0881861|Chest US
C0881861|Multisection:Finding:Point in time:Chest:Document:Ultrasound
C0881861|Multisection:Find:Pt:Chest:Doc:US
C0881995|Abd XR AP (supine+Upr) port
C0881995|Abdomen X-ray AP (supine and upright) portable
C0881995|Views AP (supine & upright) portable:Finding:Point in time:Abdomen:Document:XR
C0881995|Views AP (supine & upright) portable:Find:Pt:Abdomen:Doc:XR
C1114494|Multisection^WO & W contrast IV:Find:Pt:Pelvis+Hip:Doc:MRI
C1114494|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pelvis+Hip:Document:MRI
C1114494|Pelvis+Hip MRI WO+W contr IV
C1114494|Pelvis and Hip MRI WO and W contrast IV
C1114515|Pulm RI VP W RNC IH+IV
C1114515|Pulmonary system Scan ventilation and perfusion W radionuclide IH and W radionuclide IV
C1114515|Views ventilation & perfusion^W radionuclide IH & W radionuclide IV:Find:Pt:Pulmonary system:Doc:Radnuc
C1114515|Views ventilation & perfusion^W radionuclide Inhalation & W radionuclide Intravenous:Finding:Point in time:Pulmonary system:Document:Radnuc
C1114605|Maxillofacial CT W contr IV
C1114605|Maxillofacial region CT W contrast IV
C1114605|Multisection^W contrast IV:Find:Pt:Head>Maxillofacial region:Doc:CT
C1114605|Multisection^W contrast Intravenous:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1114617|Peritoneum Fluoroscopic angiogram W contrast percutaneous
C1114617|Peritoneum XRA W contr PC
C1114617|Views^W contrast percutaneous:Find:Pt:Peritoneum:Doc:XR.fluor.angio
C1114617|Views^W contrast percutaneous:Finding:Point in time:Peritoneum:Document:XR.fluor.angio
C1114954|Chest vessels MRI angiogram
C1114954|Chest ves MRI.Angio
C1114954|Multisection:Find:Pt:Chest vessels:Doc:MRI.angio
C1114954|Multisection:Finding:Point in time:Chest vessels:Document:MRI.angio
C1114669|LE ves MRI.Angio
C1114669|Lower extremity vessels MRI angiogram
C1114669|Multisection:Finding:Point in time:Lower extremity vessels:Document:MRI.angio
C1114669|Multisection:Find:Pt:Lower extremity vessels:Doc:MRI.angio
C1114677|Upper extremity vein US.doppler
C1114677|UE v DOP
C1114677|Multisection:Find:Pt:Upper extremity vein:Doc:US.doppler
C1114677|Multisection:Finding:Point in time:Upper extremity vein:Document:Ultrasound.doppler
C1114420|Pituitary and Sella turcica CT W contrast IV
C1114420|Multisection^W contrast IV:Find:Pt:Head>Pituitary+Sella turcica:Doc:CT
C1114420|Multisection^W contrast Intravenous:Finding:Point in time:Head>Pituitary+Sella turcica:Document:Computerized Tomography
C1114420|Head Pit+Slla turc CT W contr IV
C1114426|T-spine CT WO contr
C1114426|Multisection^WO contrast:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C1114426|Multisection^WO contrast:Find:Pt:Spine.thoracic:Doc:CT
C1114426|Thoracic spine CT WO contrast
C1114434|CT Guidance for fine needle aspiration of Pelvis
C1114434|Pelvis CT FNA Asp
C1114434|Guidance for aspiration.fine needle:Find:Pt:Pelvis:Doc:CT
C1114434|Guidance for aspiration.fine needle:Finding:Point in time:Pelvis:Document:Computerized Tomography
C1526819|Carot a.cervical-L XRA W contr IA
C1526819|Carotid artery.cervical - left Fluoroscopic angiogram W contrast IA
C1526819|Views^W contrast IA:Find:Pt:Carotid artery.cervical.left:Doc:XR.fluor.angio
C1526819|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.cervical.left:Document:XR.fluor.angio
C1543785|Hrt RI PF W DBM+ Tl-201 IV
C1543785|Heart Scan perfusion W dobutamine and W Tl-201 IV
C1543785|Views perfusion^W dobutamine & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1543785|Views perfusion^W dobutamine & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543786|Hrt SPECT PF W Stress+W RNC IV
C1543786|Heart SPECT perfusion W stress and W radionuclide IV
C1543786|Multisection perfusion^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543786|Multisection perfusion^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1542900|Lung SPECT VP W RNC IH+IV
C1542900|Multisection ventilation & perfusion^W radionuclide IH & W radionuclide IV:Find:Pt:Lung:Doc:Radnuc.SPECT
C1542900|Multisection ventilation & perfusion^W radionuclide Inhalation & W radionuclide Intravenous:Finding:Point in time:Lung:Document:Radnuc.SPECT
C1542900|Lung SPECT ventilation and perfusion W radionuclide IH and W radionuclide IV
C1543882|Multisection^W radionuclide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc.SPECT
C1543882|Kidney - bilateral SPECT
C1543882|Multisection^W radionuclide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc.SPECT
C1543882|Kdny-Bl SPECT W RNC IV
C1543522|Testicle ves DOP
C1543522|Testicle vessels US.doppler
C1543522|Multisection:Find:Pt:Testicle vessels:Doc:US.doppler
C1543522|Multisection:Finding:Point in time:Testicle vessels:Document:Ultrasound.doppler
C1543162|Deprecated Uterus+FT US W contr IU
C1543162|Multisection^W contrast intrauterine:Find:Pt:Uterus+Fallopian tubes:Nar:US
C1543162|Deprecated Uterus & Fallopian tubes US W contrast intrauterine
C1543162|Multisection^W contrast intrauterine:Finding:Point in time:Uterus+Fallopian tubes:Narrative:Ultrasound
C1543572|Upper extremity vein - bilateral US.doppler
C1543572|UE v-Bl DOP
C1543572|Multisection:Find:Pt:Upper extremity vein.bilateral:Doc:US.doppler
C1543572|Multisection:Finding:Point in time:Upper extremity vein.bilateral:Document:Ultrasound.doppler
C1543576|Upper extremity artery - left US.doppler
C1543576|UE a-L DOP
C1543576|Multisection:Find:Pt:Upper extremity artery.left:Doc:US.doppler
C1543576|Multisection:Finding:Point in time:Upper extremity artery.left:Document:Ultrasound.doppler
C1543601|Extremity US limited
C1543601|Extr US Ltd
C1543601|Multisection limited:Find:Pt:Extremity:Doc:US
C1543601|Multisection limited:Finding:Point in time:Extremity:Document:Ultrasound
C1543214|Hep vs XRA W contr IV
C1543214|Hepatic veins Fluoroscopic angiogram W contrast IV
C1543214|Views^W contrast IV:Find:Pt:Hepatic veins:Doc:XR.fluor.angio
C1543214|Views^W contrast Intravenous:Finding:Point in time:Hepatic veins:Document:XR.fluor.angio
C1543218|Carot a-Bl+Cerebral a-Bl XRA W contr IA
C1543218|Carotid artery - bilateral and Cerebral artery - bilateral Fluoroscopic angiogram W contrast IA
C1543218|Views^W contrast IA:Find:Pt:Carotid artery.bilateral+Cerebral artery.bilateral:Doc:XR.fluor.angio
C1543218|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.bilateral+Cerebral artery.bilateral:Document:XR.fluor.angio
C1524263|Should-R XR AP+Y
C1524263|Shoulder - right X-ray AP and Y
C1524263|Views AP & Y:Find:Pt:Shoulder.right:Doc:XR
C1524263|Views AP & Y:Finding:Point in time:Shoulder.right:Document:XR
C1526762|Tibia - right X-ray 10 degree caudal angle
C1526762|Tib-R XR 10 Deg Cau Angle
C1526762|View 10 degree caudal angle:Finding:Point in time:Tibia.right:Document:XR
C1526762|View 10 degree caudal angle:Find:Pt:Tibia.right:Doc:XR
C1543715|Heart Scan for infarct
C1543715|Hrt RI for Infarct W RNC IV
C1543715|Views for infarct^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543715|Views for infarct^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543724|Hrt SPECT Rest+stress+W Tc99mMIBI IV
C1543724|Heart SPECT at rest and W stress and W Tc-99m Sestamibi IV
C1543724|Multisection^at rest & W stress & W Tc-99m Sestamibi Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1543724|Multisection^at rest & W stress & W Tc-99m Sestamibi IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543731|RI WB W Tc99mCEA IV
C1543731|Scan whole body W Tc-99m Arcitumomab IV
C1543731|Views whole body^W Tc-99m Arcitumomab Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543731|Views whole body^W Tc-99m Arcitumomab IV:Find:Pt:^Patient:Doc:Radnuc
C1524189|Portal v MRI.Angio
C1524189|Portal vein MRI angiogram
C1524189|Multisection:Find:Pt:Portal vein:Doc:MRI.angio
C1524189|Multisection:Finding:Point in time:Portal vein:Document:MRI.angio
C1524836|LE-Bl MRI WO contr
C1524836|Lower extremity - bilateral MRI WO contrast
C1524836|Multisection^WO contrast:Find:Pt:Lower extremity.bilateral:Doc:MRI
C1524836|Multisection^WO contrast:Finding:Point in time:Lower extremity.bilateral:Document:MRI
C1527064|Orbit MRI
C1527064|Multisection:Finding:Point in time:Orbit:Narrative:MRI
C1527064|Multisection:Find:Pt:Orbit:Doc:MRI
C1527064|Multisection:Finding:Point in time:Orbit:Document:MRI
C1525180|Renal ves-Bl MRI.Angio
C1525180|Renal vessels - bilateral MRI angiogram
C1525180|Multisection:Find:Pt:Renal vessels.bilateral:Doc:MRI.angio
C1525180|Multisection:Finding:Point in time:Renal vessels.bilateral:Document:MRI.angio
C1524443|Internal auditory canal MRI limited
C1524443|IAC MRI Ltd
C1524443|Multisection limited:Find:Pt:Internal auditory canal:Doc:MRI
C1524443|Multisection limited:Finding:Point in time:Internal auditory canal:Document:MRI
C1524234|Brain MRI Ltd WO contr
C1524234|Brain MRI limited WO contrast
C1524234|Multisection limited^WO contrast:Finding:Point in time:Brain:Document:MRI
C1524234|Multisection limited^WO contrast:Find:Pt:Brain:Doc:MRI
C1525287|Thyroid CT WO contr
C1525287|Thyroid CT WO contrast
C1525287|Multisection^WO contrast:Find:Pt:Thyroid:Doc:CT
C1525287|Multisection^WO contrast:Finding:Point in time:Thyroid:Document:Computerized Tomography
C1525302|View decubitus portable:Find:Pt:Abdomen:Nar:XR
C1525302|Deprecated View decubitus portable
C1525302|Deprecated Abd XR Decub Port
C1525302|View decubitus portable:Finding:Point in time:Abdomen:Narrative:XR
C1525321|C-spine XR Lat Xtable
C1525321|View lateral crosstable:Finding:Point in time:Spine.cervical:Document:XR
C1525321|View lateral crosstable:Find:Pt:Spine.cervical:Doc:XR
C1525321|Cervical spine X-ray lateral crosstable
C3853708|Orbit MRI W contr IV
C3853708|Orbit MRI W contrast IV
C3853708|Multisection^W contrast IV:Find:Pt:Orbit:Doc:MRI
C3853708|Multisection^W contrast Intravenous:Finding:Point in time:Orbit:Document:MRI
C1525223|Lower extremity veins - left MRI angiogram WO and W contrast IV
C1525223|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower extremity veins.left:Document:MRI.angio
C1525223|LE vv-L MRI.Angio WO+W contr IV
C1525223|Multisection^WO & W contrast IV:Find:Pt:Lower extremity veins.left:Doc:MRI.angio
C1525276|Multisection^WO & W contrast IV:Find:Pt:Biliary ducts+Pancreatic duct:Doc:MRI
C1525276|Biliary ducts and Pancreatic duct MRI WO and W contrast IV
C1525276|Multisection^WO & W contrast Intravenous:Finding:Point in time:Biliary ducts+Pancreatic duct:Document:MRI
C1525276|BD+PDs MRI WO+W contr IV
C1525329|C-spine XR Lat W Ext
C1525329|View lateral^W extension:Find:Pt:Spine.cervical:Doc:XR
C1525329|View lateral^W extension:Finding:Point in time:Spine.cervical:Document:XR
C1525329|Cervical spine X-ray lateral W extension
C1525467|Knee - bilateral X-ray tunnel
C1525467|Knee-Bl XR V1 Tunnel
C1525467|View tunnel:Find:Pt:Knee.bilateral:Doc:XR
C1525467|View tunnel:Finding:Point in time:Knee.bilateral:Document:XR
C1525518|Knee-Bl XR AP+Lat+Obl+Sunrise+Tunnel
C1525518|Knee - bilateral X-ray AP and lateral and oblique and Sunrise and tunnel
C1525518|Views AP & lateral & oblique & Sunrise & tunnel:Find:Pt:Knee.bilateral:Doc:XR
C1525518|Views AP & lateral & oblique & Sunrise & tunnel:Finding:Point in time:Knee.bilateral:Document:XR
C1525544|Chest XR PA+Lat+AP R-Lat-Decub
C1525544|Chest X-ray PA and lateral and AP right lateral-decubitus
C1525544|Views PA & lateral & AP R-lateral-decubitus:Find:Pt:Chest:Doc:XR
C1525544|Views PA & lateral & AP R-lateral-decubitus:Finding:Point in time:Chest:Document:XR
C1525546|Chest XR PA+Lat+R-Obl
C1525546|Chest X-ray PA and lateral and right oblique
C1525546|Views PA & lateral & R-oblique:Find:Pt:Chest:Doc:XR
C1525546|Views PA & lateral & R-oblique:Finding:Point in time:Chest:Document:XR
C1525579|PA-L XRA W contr IA
C1525579|Views^W contrast Intra-arterial:Finding:Point in time:Pulmonary artery.left:Document:XR.fluor.angio
C1525579|Views^W contrast IA:Find:Pt:Pulmonary artery.left:Doc:XR.fluor.angio
C1525579|Left pulmonary artery Fluoroscopic angiogram W contrast IA
C1525661|Brain+Larynx MRI WO contr
C1525661|Brain and Larynx MRI WO contrast
C1525661|Multisection^WO contrast:Find:Pt:Brain+Larynx:Doc:MRI
C1525661|Multisection^WO contrast:Finding:Point in time:Brain+Larynx:Document:MRI
C1525670|Spine Lumbosacral Junction CT WO contrast
C1525670|LS-spine junc CT WO contr
C1525670|Multisection^WO contrast:Finding:Point in time:Spine.lumbosacral junction:Document:Computerized Tomography
C1525670|Multisection^WO contrast:Find:Pt:Spine.lumbosacral junction:Doc:CT
C1525716|Carotid artery.external - left Fluoroscopic angiogram W contrast IA
C1525716|Carot a.ext-L XRA W contr IA
C1525716|Views^W contrast IA:Find:Pt:Carotid artery.external.left:Doc:XR.fluor.angio
C1525716|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.external.left:Document:XR.fluor.angio
C1525725|Gastroduodenal artery Fluoroscopic angiogram W contrast IA
C1525725|Gastroduodenal a XRA W contr IA
C1525725|Views^W contrast IA:Find:Pt:Gastroduodenal artery:Doc:XR.fluor.angio
C1525725|Views^W contrast Intra-arterial:Finding:Point in time:Gastroduodenal artery:Document:XR.fluor.angio
C1525732|Vertebral artery - bilateral Fluoroscopic angiogram W contrast IA
C1525732|VA-Bl XRA W contr IA
C1525732|Views^W contrast IA:Find:Pt:Vertebral artery.bilateral:Doc:XR.fluor.angio
C1525732|Views^W contrast Intra-arterial:Finding:Point in time:Vertebral artery.bilateral:Document:XR.fluor.angio
C1525848|Brst-Bl Mam Spot
C1525848|Breast - bilateral Mammogram spot
C1525848|Views spot:Finding:Point in time:Breast.bilateral:Document:Mam
C1525848|Views spot:Find:Pt:Breast.bilateral:Doc:Mam
C1524143|Lymphatics - left Fluoroscopy W contrast intra lymphatic
C1524143|Lymph-L Flr W contr IL
C1524143|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.left:Doc:XR.fluor
C1524143|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.left:Document:XR.fluor
C1525938|Pelvis XR AP+Lat
C1525938|Pelvis X-ray AP and lateral
C1525938|Views AP & lateral:Finding:Point in time:Pelvis:Document:XR
C1525938|Views AP & lateral:Find:Pt:Pelvis:Doc:XR
C1525946|Pelvis X-ray inlet
C1525946|Pelvis XR Inlet
C1525946|View inlet:Find:Pt:Pelvis:Doc:XR
C1525946|View inlet:Finding:Point in time:Pelvis:Document:XR
C1525977|AC joint-R XR 2V
C1525977|Acromioclavicular joint - right X-ray 2 views
C1525977|Views 2:Find:Pt:Acromioclavicular joint.right:Doc:XR
C1525977|Views 2:Finding:Point in time:Acromioclavicular joint.right:Document:XR
C1525982|Ankle-R XR AP+Lat+Mortise
C1525982|Ankle - right X-ray AP and lateral and Mortise
C1525982|Views AP & lateral & Mortise:Finding:Point in time:Ankle.right:Document:XR
C1525982|Views AP & lateral & Mortise:Find:Pt:Ankle.right:Doc:XR
C1525897|Wrist-R XR 3V
C1525897|Wrist - right X-ray 3 views
C1525897|Views 3:Find:Pt:Wrist.right:Doc:XR
C1525897|Views 3:Finding:Point in time:Wrist.right:Document:XR
C1525897|VIEWS 3:FINDING:POINT IN TIME:WRIST.RIGHT:NARRATIVE:XR
C1525901|Wrist-R XR 8V
C1525901|Wrist - right X-ray 8 views
C1525901|Views 8:Find:Pt:Wrist.right:Doc:XR
C1525901|Views 8:Finding:Point in time:Wrist.right:Document:XR
C1526044|Hip - right X-ray oblique crosstable
C1526044|Hip-R XR Obl Xtable
C1526044|View oblique crosstable:Find:Pt:Hip.right:Doc:XR
C1526044|View oblique crosstable:Finding:Point in time:Hip.right:Document:XR
C1526047|Hip - right X-ray standing
C1526047|Hip-R XR stand
C1526047|View^standing:Find:Pt:Hip.right:Doc:XR
C1526047|View^standing:Finding:Point in time:Hip.right:Document:XR
C1526083|LE vv-R XRA W contr IV
C1526083|Lower extremity veins - right Fluoroscopic angiogram W contrast IV
C1526083|Views^W contrast IV:Find:Pt:Lower extremity veins.right:Doc:XR.fluor.angio
C1526083|Views^W contrast Intravenous:Finding:Point in time:Lower extremity veins.right:Document:XR.fluor.angio
C1525122|Brst-R Mam XCCL
C1525122|Breast - right Mammogram XCCL
C1525122|View XCCL:Find:Pt:Breast.right:Doc:Mam
C1525122|View XCCL:Finding:Point in time:Breast.right:Document:Mam
C1525123|Breast - right Mammogram magnification
C1525123|Brst-R Mam Mag
C1525123|View magnification:Finding:Point in time:Breast.right:Document:Mam
C1525123|View magnification:Find:Pt:Breast.right:Doc:Mam
C1526091|Sacroiliac joint - right X-ray
C1526091|SIJ-R XR
C1526091|Views:Finding:Point in time:Sacroiliac joint.right:Document:XR
C1526091|Views:Find:Pt:Sacroiliac joint.right:Doc:XR
C1526093|Scapula-R XR AP+Lat
C1526093|Scapula - right X-ray AP and lateral
C1526093|Views AP & lateral:Find:Pt:Scapula.right:Doc:XR
C1526093|Views AP & lateral:Finding:Point in time:Scapula.right:Document:XR
C1526098|Shoulder - right X-ray 2 views
C1526098|Should-R XR 2V
C1526098|Views 2:Find:Pt:Shoulder.right:Doc:XR
C1526098|Views 2:Finding:Point in time:Shoulder.right:Document:XR
C1526152|Sinuses XR PA+Lat+Caldwell+Waters
C1526152|Sinuses X-ray PA and lateral and Caldwell and Waters
C1526152|Views PA & lateral & Caldwell & Waters:Find:Pt:Sinuses:Doc:XR
C1526152|Views PA & lateral & Caldwell & Waters:Finding:Point in time:Sinuses:Document:XR
C1524268|Spine X-ray 2 views
C1524268|Spine XR 2V
C1524268|Views 2:Find:Pt:Spine:Doc:XR
C1524268|Views 2:Finding:Point in time:Spine:Document:XR
C1526174|Tib+Fib XR 1V
C1526174|Tibia and Fibula X-ray Single view
C1526174|View 1:Finding:Point in time:Tibia+Fibula:Document:XR
C1526174|View 1:Find:Pt:Tibia+Fibula:Doc:XR
C1524705|Wrist XR AP+Lat+Obl
C1524705|Wrist X-ray AP and lateral and oblique
C1524705|Views AP & lateral & oblique:Find:Pt:Wrist:Doc:XR
C1524705|Views AP & lateral & oblique:Finding:Point in time:Wrist:Document:XR
C1524706|Wrist X-ray Brewerton
C1524706|Wrist XR Brewerton
C1524706|View Brewerton:Finding:Point in time:Wrist:Document:XR
C1524706|View Brewerton:Find:Pt:Wrist:Doc:XR
C1526222|Jugular v-R XRA W contr IV
C1526222|Jugular vein - right Fluoroscopic angiogram W contrast IV
C1526222|Views^W contrast Intravenous:Finding:Point in time:Jugular vein.right:Document:XR.fluor.angio
C1526222|Views^W contrast IV:Find:Pt:Jugular vein.right:Doc:XR.fluor.angio
C1526267|Brst-L US FNA Asp
C1526267|US Guidance for fine needle aspiration of Breast - left
C1526267|Guidance for aspiration.fine needle:Finding:Point in time:Breast.left:Document:Ultrasound
C1526267|Guidance for aspiration.fine needle:Find:Pt:Breast.left:Doc:US
C1525910|C+T+L-spine Flr Ltd W contr IT
C1525910|Spine Cervical and Thoracic and Lumbar Fluoroscopy limited W contrast IT
C1525910|Views limited^W contrast IT:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:XR.fluor
C1525910|Views limited^W contrast Intrathecal:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:XR.fluor
C1525911|Kidney US Cyst Asp guid
C1525911|US Guidance for aspiration of cyst of Kidney
C1525911|Guidance for aspiration of cyst:Finding:Point in time:Kidney:Document:Ultrasound
C1525911|Guidance for aspiration of cyst:Find:Pt:Kidney:Doc:US
C1525913|Femoral vessels - bilateral US
C1525913|Fem ves-Bl US
C1525913|Multisection:Finding:Point in time:Femoral vessels.bilateral:Document:Ultrasound
C1525913|Multisection:Find:Pt:Femoral vessels.bilateral:Doc:US
C1525919|Fem ves US
C1525919|Femoral vessels US
C1525919|Multisection:Find:Pt:Femoral vessels:Doc:US
C1525919|Multisection:Finding:Point in time:Femoral vessels:Document:Ultrasound
C1526298|Breast implant Mammogram
C1526298|Brst implant Mam
C1526298|Views:Find:Pt:Breast implant:Doc:Mam
C1526298|Views:Finding:Point in time:Breast implant:Document:Mam
C1526306|C-spine XR AP+Lat+Obl+Odont+Swimmer
C1526306|Views AP & lateral & oblique & odontoid & swimmer:Find:Pt:Spine.cervical:Doc:XR
C1526306|Views AP & lateral & oblique & odontoid & swimmer:Finding:Point in time:Spine.cervical:Document:XR
C1526306|Cervical spine X-ray AP and lateral and oblique and odontoid and swimmer
C1526311|Chest XR W nipple markers
C1526311|Chest X-ray W nipple markers
C1526311|Views^W nipple markers:Finding:Point in time:Chest:Document:XR
C1526311|Views^W nipple markers:Find:Pt:Chest:Doc:XR
C1526317|Lacrimal duct - left Fluoroscopy W contrast intra lacrimal duct
C1526317|Lacrimal duct-L Flr W contr intra LD
C1526317|Views^W contrast intra lacrimal duct:Find:Pt:Lacrimal duct.left:Doc:XR.fluor
C1526317|Views^W contrast intra lacrimal duct:Finding:Point in time:Lacrimal duct.left:Document:XR.fluor
C1526320|Kidney XR W contr Ante via Pyelostomy
C1526320|Views^W contrast antegrade via pyelostomy:Find:Pt:Kidney:Doc:XR
C1526320|Views^W contrast antegrade via pyelostomy:Finding:Point in time:Kidney:Document:XR
C1526320|Kidney X-ray W contrast antegrade via pyelostomy
C1524496|Brst-R MRI W contr IV
C1524496|Breast - right MRI W contrast IV
C1524496|Multisection^W contrast IV:Find:Pt:Breast.right:Doc:MRI
C1524496|Multisection^W contrast Intravenous:Finding:Point in time:Breast.right:Document:MRI
C1524510|LE-R CT W contr IV
C1524510|Lower extremity - right CT W contrast IV
C1524510|Multisection^W contrast IV:Find:Pt:Lower extremity.right:Doc:CT
C1524510|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.right:Document:Computerized Tomography
C1524863|Hand-L CT WO contr
C1524863|Hand - left CT WO contrast
C1524863|Multisection^WO contrast:Finding:Point in time:Hand.left:Document:Computerized Tomography
C1524863|Multisection^WO contrast:Find:Pt:Hand.left:Doc:CT
C1524528|Ft-R MRI W contr IV
C1524528|Foot - right MRI W contrast IV
C1524528|Multisection^W contrast IV:Find:Pt:Foot.right:Doc:MRI
C1524528|Multisection^W contrast Intravenous:Finding:Point in time:Foot.right:Document:MRI
C1524934|Femur - left X-ray Single view
C1524934|Femur-L XR 1V
C1524934|View 1:Finding:Point in time:Femur.left:Document:XR
C1524934|View 1:Find:Pt:Femur.left:Doc:XR
C1524944|Finger second X-ray lateral
C1524944|Finger.2nd XR Lat
C1524944|View lateral:Find:Pt:Finger.second:Doc:XR
C1524944|View lateral:Finding:Point in time:Finger.second:Document:XR
C1524287|Fluoroscopy Guidance for aspiration of Hip
C1524287|Hip Flr Asp guid
C1524287|Guidance for aspiration:Find:Pt:Hip:Doc:XR.fluor
C1524287|Guidance for aspiration:Finding:Point in time:Hip:Document:XR.fluor
C1524612|Elbow - left CT WO and W contrast IV
C1524612|Multisection^WO & W contrast Intravenous:Finding:Point in time:Elbow.left:Document:Computerized Tomography
C1524612|Elbow-L CT WO+W contr IV
C1524612|Multisection^WO & W contrast IV:Find:Pt:Elbow.left:Doc:CT
C1524972|Wrist - bilateral X-ray PA
C1524972|Wrist-Bl XR PA V1
C1524972|View PA:Find:Pt:Wrist.bilateral:Doc:XR
C1524972|View PA:Finding:Point in time:Wrist.bilateral:Document:XR
C1524342|Ankle - right CT
C1524342|Ankle-R CT
C1524342|Multisection:Finding:Point in time:Ankle.right:Document:Computerized Tomography
C1524342|Multisection:Find:Pt:Ankle.right:Doc:CT
C1525000|Femur X-ray 2 views
C1525000|Femur XR 2V
C1525000|Views 2:Find:Pt:Femur:Doc:XR
C1525000|Views 2:Finding:Point in time:Femur:Document:XR
C1525015|Knee - left X-ray 5 views
C1525015|Knee-L XR 5V
C1525015|Views 5:Find:Pt:Knee.left:Doc:XR
C1525015|Views 5:Finding:Point in time:Knee.left:Document:XR
C1525018|Should-L XR 6V
C1525018|Shoulder - left X-ray 6 views
C1525018|Views 6:Find:Pt:Shoulder.left:Doc:XR
C1525018|Views 6:Finding:Point in time:Shoulder.left:Document:XR
C1524369|Lower extremity - bilateral MRI
C1524369|LE-Bl MRI
C1524369|Multisection:Find:Pt:Lower extremity.bilateral:Doc:MRI
C1524369|Multisection:Finding:Point in time:Lower extremity.bilateral:Document:MRI
C1525026|Chest XR AP+Lat
C1525026|Chest X-ray AP and lateral
C1525026|Views AP & lateral:Finding:Point in time:Chest:Document:XR
C1525026|Views AP & lateral:Find:Pt:Chest:Doc:XR
C1524397|Hand - left X-ray tomograph
C1524397|Hand-L XRTomo
C1524397|Multisection:Find:Pt:Hand.left:Doc:XR.tomo
C1524397|Multisection:Finding:Point in time:Hand.left:Document:XR.tomo
C1527046|Hip CT
C1527046|Multisection:Find:Pt:Hip:Doc:CT
C1527046|Multisection:Finding:Point in time:Hip:Document:Computerized Tomography
C1524768|Larynx MRI WO+W contr IV
C1524768|Multisection^WO & W contrast IV:Find:Pt:Larynx:Doc:MRI
C1524768|Larynx MRI WO and W contrast IV
C1524768|Multisection^WO & W contrast Intravenous:Finding:Point in time:Larynx:Document:MRI
C1525087|Chest XR PA+Lordotic
C1525087|Chest X-ray PA and lordotic
C1525087|Views PA & lordotic:Find:Pt:Chest:Doc:XR
C1525087|Views PA & lordotic:Finding:Point in time:Chest:Document:XR
C1830218|Chest CT WO+W red contr vol IV
C1830218|Multisection^WO & W reduced contrast volume Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C1830218|Multisection^WO & W reduced contrast volume IV:Find:Pt:Chest:Doc:CT
C1830218|Chest CT WO and W reduced contrast volume IV
C1830222|Orbit+Face+Neck MRI W contr IV
C1830222|Orbit and Face and Neck MRI W contrast IV
C1830222|Multisection^W contrast IV:Find:Pt:Orbit+Face+Neck:Doc:MRI
C1830222|Multisection^W contrast Intravenous:Finding:Point in time:Orbit+Face+Neck:Document:MRI
C1830225|LE ves MRI.Angio W contr IV
C1830225|Lower extremity vessels MRI angiogram W contrast IV
C1830225|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity vessels:Document:MRI.angio
C1830225|Multisection^W contrast IV:Find:Pt:Lower extremity vessels:Doc:MRI.angio
C1830231|Abd CT W red contr vol IV
C1830231|Abdomen CT W reduced contrast volume IV
C1830231|Multisection^W reduced contrast volume IV:Find:Pt:Abdomen:Doc:CT
C1830231|Multisection^W reduced contrast volume Intravenous:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1830249|Chest XR GE 2 & PA+Lat
C1830249|Chest X-ray GE 2 and PA and Lateral views
C1830249|Views GE 2 & PA & lateral:Find:Pt:Chest:Doc:XR
C1830249|Views GE 2 & PA & lateral:Finding:Point in time:Chest:Document:XR
C1830252|Breast implant - bilateral Mammogram displacement
C1830252|Brst implant-Bl Mam Displacement
C1830252|Views displacement:Finding:Point in time:Breast implant.bilateral:Document:Mam
C1830252|Views displacement:Find:Pt:Breast implant.bilateral:Doc:Mam
C1830282|Liver CT W 133Xe IH
C1830282|Multisection^W Xe-133 IH:Find:Pt:Abdomen>Liver:Doc:CT
C1830282|Multisection^W Xe-133 Inhalation:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1830282|Liver CT W Xe-133 IH
C1715443|L-spine XR Obl1V+(views W R+L-bending)
C1715443|View oblique & (Views^W R-bending & W L-bending):Find:Pt:Spine.lumbar:Doc:XR
C1715443|View oblique & (Views^W R-bending & W L-bending):Finding:Point in time:Spine.lumbar:Document:XR
C1715443|Lumbar spine X-ray oblique view and (views W right bending and W left bending)
C1715453|Sacroiliac Joint X-ray GE 3 views
C1715453|SIJ XR GE 3V
C1715453|Views GE 3:Find:Pt:Sacroiliac joint:Doc:XR
C1715453|Views GE 3:Finding:Point in time:Sacroiliac joint:Document:XR
C1651656|Deprecated Views:Finding:Point in time:Tibia.left:Narrative:XR
C1651656|Views:Find:Pt:Tibia.left:Nar:XR
C1651656|Deprecated Tib-L XR
C1651656|Views:Finding:Point in time:Tibia.left:Narrative:XR
C1651656|Deprecated Tibia Left X-ray
C1714804|Chest XR 2V+R-Obl+L-Obl
C1714804|Chest X-ray 2 views and right oblique and left oblique
C1714804|Views 2 & R-Oblique & L-Oblique:Find:Pt:Chest:Doc:XR
C1714804|Views 2 & R-Oblique & L-Oblique:Finding:Point in time:Chest:Document:XR
C1706620|Finger fifth - right X-ray GE 3 views
C1706620|Finger.5th-R XR GE 3V
C1706620|Finger fifth - right Narrative X-ray GE 3 views
C1706620|Views GE 3:Finding:Point in time:Finger.fifth.right:Document:XR
C1706620|Views GE 3:Find:Pt:Finger.fifth.right:Doc:XR
C1717259|Views:Find:Pt:Mandible.right:Doc:XR
C1717259|Deprecated Mandible - right X-ray
C1717259|Views:Finding:Point in time:Mandible.right:Document:XR
C1717259|Deprecated Mandible-R XR
C1714940|Guidance for abscess drainage:Find:Pt:Peritoneal cavity:Nar:US
C1714940|Deprecated Perit Cavity US Abs drain gui
C1714940|Deprecated US Guidance for abscess drainage of Peritoneal cavity
C1714940|Guidance for abscess drainage:Finding:Point in time:Peritoneal cavity:Narrative:Ultrasound
C1714507|Kidney CT FNA Asp
C1714507|CT Guidance for fine needle aspiration of Kidney
C1714507|Guidance for aspiration.fine needle:Finding:Point in time:Kidney:Document:Computerized Tomography
C1714507|Guidance for aspiration.fine needle:Find:Pt:Kidney:Doc:CT
C1715112|Views AP (supine KUB & upright) & PA upright chest:Find:Pt:Abdomen+Chest:Nar:XR
C1715112|Deprecated Abdomen & Chest X-ray AP (supine & upright) & PA chest
C1715112|Deprecated Abd+Chest XR AP(supKUB+Upr)+P
C1715112|Views AP (supine KUB & upright) & PA upright chest:Finding:Point in time:Abdomen+Chest:Narrative:XR
C1715113|Skull+Face+Mandible XR For Dent Meas
C1715113|Skull and Facial bones and Mandible X-ray for dental measurement
C1715113|Views for dental measurement:Find:Pt:Skull+Facial bones+Mandible:Doc:XR
C1715113|Views for dental measurement:Finding:Point in time:Skull+Facial bones+Mandible:Document:XR
C1637284|Spine XR Lat stand
C1637284|Spine X-ray lateral standing
C1637284|View lateral^standing:Finding:Point in time:Spine:Document:XR
C1637284|View lateral^standing:Find:Pt:Spine:Doc:XR
C1623575|Gastrointestine upper Fluoroscopy W water soluble contrast PO
C1623575|UGI Flr W H2O soluble contr PO
C1623575|Views^W water soluble contrast Oral:Finding:Point in time:Gastrointestine.upper:Document:XR.fluor
C1623575|Views^W water soluble contrast PO:Find:Pt:Gastrointestine.upper:Doc:XR.fluor
C1635017|Submandib gland-L Flr W contr intra SD
C1635017|Submandibular gland - left Fluoroscopy W contrast intra salivary duct
C1635017|Views^W contrast intra salivary duct:Find:Pt:Submandibular gland.left:Doc:XR.fluor
C1635017|Views^W contrast intra salivary duct:Finding:Point in time:Submandibular gland.left:Document:XR.fluor
C1626843|UGI+SB+GB Flr W contr PO
C1626843|Gastrointestine upper and Small bowel and Gallbladder Fluoroscopy W contrast PO
C1626843|View^W contrast Oral:Finding:Point in time:Gastrointestine.upper+Small bowel+Gallbladder:Document:XR.fluor
C1626843|View^W contrast PO:Find:Pt:Gastrointestine.upper+Small bowel+Gallbladder:Doc:XR.fluor
C1645732|T+L-spine XR Scoli AP In Traction
C1645732|Views scoliosis AP^in traction:Find:Pt:Spine.thoracic+Spine.lumbar:Doc:XR
C1645732|Spine Thoracic and Lumbar X-ray scoliosis AP in traction
C1645732|Views scoliosis AP^in traction:Finding:Point in time:Spine.thoracic+Spine.lumbar:Document:XR
C1631255|Deprecated L-spine W Non-ionic contr IT
C1631255|Views^W non-ionic contrast IT:Find:Pt:Spine.lumbar:Nar
C1631255|Deprecated Spine Lumbar X-ray fluoroscopy W contrast IT
C1631255|Views^W non-ionic contrast Intrathecal:Finding:Point in time:Spine.lumbar:Narrative
C1632225|Mammogram Guidance for localization of Breast - left
C1632225|Brst-L Mam Localization guid
C1632225|Guidance for localization:Find:Pt:Breast.left:Doc:Mam
C1632225|Guidance for localization:Finding:Point in time:Breast.left:Document:Mam
C1953977|Mastoid - left X-ray 3 views
C1953977|Mastoid-L XR 3V
C1953977|Views 3:Find:Pt:Mastoid.left:Doc:XR
C1953977|Views 3:Finding:Point in time:Mastoid.left:Document:XR
C3262935|Multisection^W contrast Intrasynovial:Finding:Point in time:Hip.right:Document:Computerized Tomography
C3262935|Multisection^W contrast IS:Find:Pt:Hip.right:Doc:CT
C3262935|Hip-R CT W contr IS
C3262935|Hip - right CT W contrast IS
C3262971|Patella - left X-ray Single view
C3262971|Patella-L XR 1V
C3262971|View 1:Find:Pt:Patella.left:Doc:XR
C3262971|View 1:Finding:Point in time:Patella.left:Document:XR
C3262979|Brst Mam Bx needle Str Guid
C3262979|Guidance for stereotactic biopsy.needle:Finding:Point in time:Breast:Document:Mam
C3262979|Guidance for stereotactic biopsy.needle:Find:Pt:Breast:Doc:Mam
C3262979|Mammogram Guidance for stereotactic needle biopsy of Breast
C3263070|LE-R XR AP+Lat
C3263070|Lower extremity - right X-ray AP and lateral
C3263070|Views AP & lateral:Finding:Point in time:Lower extremity.right:Document:XR
C3263070|Views AP & lateral:Find:Pt:Lower extremity.right:Doc:XR
C3262901|Fluoroscopy Guidance for drainage of Chest
C3262901|Chest Flr Drain guid
C3262901|Guidance for drainage:Find:Pt:Chest:Doc:XR.fluor
C3262901|Guidance for drainage:Finding:Point in time:Chest:Document:XR.fluor
C3262928|Multisection^W contrast Intrasynovial:Finding:Point in time:Hip.left:Document:Computerized Tomography
C3262928|Multisection^W contrast IS:Find:Pt:Hip.left:Doc:CT
C3262928|Hip-L CT W contr IS
C3262928|Hip - left CT W contrast IS
C0942219|Brst-L US
C0942219|Breast - left US
C0942219|Multisection:Finding:Point in time:Breast.left:Document:Ultrasound
C0942219|Multisection:Find:Pt:Breast.left:Doc:US
C0942221|Carotid artery - left US
C0942221|Carot a-L US
C0942221|Multisection:Finding:Point in time:Carotid artery.left:Document:Ultrasound
C0942221|Multisection:Find:Pt:Carotid artery.left:Doc:US
C0945335|Fluoroscopic angiogram Guidance for placement of stent in Vein - right
C0945335|Vein-R XRA Stent plac guid
C0945335|Guidance for placement of stent:Finding:Point in time:Vein.right:Document:XR.fluor.angio
C0945335|Guidance for placement of stent:Find:Pt:Vein.right:Doc:XR.fluor.angio
C0942360|Hand-R XR 3V
C0942360|Hand - right X-ray 3 views
C0942360|Views 3:Find:Pt:Hand.right:Doc:XR
C0942360|Views 3:Finding:Point in time:Hand.right:Document:XR
C0882026|Meckels divertic RI W Tc99mM04 IV
C0882026|Meckels diverticulum Scan W Tc-99m M04 IV
C0882026|Views^W Tc-99m M04 Intravenous:Finding:Point in time:Meckels diverticulum:Document:Radnuc
C0882026|Views^W Tc-99m M04 IV:Find:Pt:Meckels diverticulum:Doc:Radnuc
C0882051|Pancreas CT W contr IV
C0882051|Pancreas CT W contrast IV
C0882051|Multisection^W contrast IV:Find:Pt:Abdomen>Pancreas:Doc:CT
C0882051|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen>Pancreas:Document:Computerized Tomography
C0882102|Skull XR AP+Lat
C0882102|Skull X-ray AP and lateral
C0882102|Views AP & lateral:Finding:Point in time:Skull:Document:XR
C0882102|Views AP & lateral:Find:Pt:Skull:Doc:XR
C0882550|SB Flr W Pos Cntrst Enteroclysis Tube
C0882550|Views^W positive contrast via enteroclysis tube:Finding:Point in time:Small bowel:Document:XR.fluor
C0882550|Views^W positive contrast via enteroclysis tube:Find:Pt:Small bowel:Doc:XR.fluor
C0882550|Small bowel Fluoroscopy W positive contrast via enteroclysis tube
C3853709|C-spine XR
C3853709|Views:Finding:Point in time:Spine.cervical:Document:XR
C3853709|Views:Find:Pt:Spine.cervical:Doc:XR
C3853709|Cervical spine X-ray
C0882126|L-spine CT
C0882126|Multisection:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C0882126|Multisection:Find:Pt:Spine.lumbar:Doc:CT
C0882126|Lumbar spine CT
C0882131|L-spine XR Lat
C0882131|View lateral:Finding:Point in time:Spine.lumbar:Document:XR
C0882131|View lateral:Find:Pt:Spine.lumbar:Doc:XR
C0882131|Lumbar spine X-ray lateral
C0882148|Multisection:Finding:Point in time:Spleen:Narrative:COMPUTERIZED TOMOGRAPHY
C0882148|Spleen CT
C0882148|Multisection:Find:Pt:Abdomen>Spleen:Doc:CT
C0882148|Multisection:Finding:Point in time:Abdomen>Spleen:Document:Computerized Tomography
C0882160|Views:Finding:Point in time:Temporomandibular joint:Narrative:XR
C0882160|TMJ XR
C0882160|Temporomandibular joint X-ray
C0882160|Views:Find:Pt:Temporomandibular joint:Doc:XR
C0882160|Views:Finding:Point in time:Temporomandibular joint:Document:XR
C0882182|IVC XRA Filter plac guid W contr IV
C0882182|Fluoroscopic angiogram Guidance for placement of IVC filter in Inferior vena cava-- W contrast IV
C0882182|Guidance for placement of IVC filter^W contrast Intravenous:Finding:Point in time:Vena cava.inferior:Document:XR.fluor.angio
C0882182|Guidance for placement of IVC filter^W contrast IV:Find:Pt:Vena cava.inferior:Doc:XR.fluor.angio
C0882565|Unspecified body region Fluoroscopy 1 hour
C0882565|XXX Flr 1h
C0882565|View:Find:1H:XXX:Doc:XR.fluor
C0882565|View:Finding:1 hour:To be specified in another part of the message:Document:XR.fluor
C0882221|XXX XRTomo
C0882221|Unspecified body region X-ray tomograph
C0882221|Multisection:Find:Pt:XXX:Doc:XR.tomo
C0882221|Multisection:Finding:Point in time:To be specified in another part of the message:Document:XR.tomo
C0945305|Salivary gland-Bl Flr W contr intra SD
C0945305|Salivary gland - bilateral Fluoroscopy W contrast intra salivary duct
C0945305|Views^W contrast intra salivary duct:Finding:Point in time:Salivary gland.bilateral:Document:XR.fluor
C0945305|Views^W contrast intra salivary duct:Find:Pt:Salivary gland.bilateral:Doc:XR.fluor
C0945309|Elbow-L XR
C0945309|Elbow - left X-ray
C0945309|Views:Find:Pt:Elbow.left:Doc:XR
C0945309|Views:Finding:Point in time:Elbow.left:Document:XR
C0881781|Views:Finding:Point in time:Ankle:Narrative:XR
C0881781|Ankle XR
C0881781|Ankle X-ray
C0881781|Views:Find:Pt:Ankle:Doc:XR
C0881781|Views:Finding:Point in time:Ankle:Document:XR
C0881792|IC ves XRA Embolectomy W contr IV
C0881792|Vessel intracranial Fluoroscopic angiogram Embolectomy W contrast IV
C0881792|Embolectomy^W contrast IV:Find:Pt:Intracranial vessel:Doc:XR.fluor.angio
C0881792|Embolectomy^W contrast Intravenous:Finding:Point in time:Intracranial vessel:Document:XR.fluor.angio
C0881794|Fluoroscopic angiogram Guidance for placement of stent in Artery
C0881794|Artery XRA Stent plac guid
C0881794|Guidance for placement of stent:Finding:Point in time:To be specified in another part of the message artery:Document:XR.fluor.angio
C0881794|Guidance for placement of stent:Find:Pt:XXX artery:Doc:XR.fluor.angio
C0881802|Abd XR AP R-Lat Decub
C0881802|Abdomen X-ray AP right lateral-decubitus
C0881802|View AP R-lateral-decubitus:Find:Pt:Abdomen:Doc:XR
C0881802|View AP R-lateral-decubitus:Finding:Point in time:Abdomen:Document:XR
C0881809|Fluoroscopy Guidance for stone removal of Biliary duct common-- W contrast intra biliary duct
C0881809|CBD Flr Stone rem guid W contr intra BD
C0881809|Guidance for stone removal^W contrast intra biliary duct:Find:Pt:Biliary duct.common:Doc:XR.fluor
C0881809|Guidance for stone removal^W contrast intra biliary duct:Finding:Point in time:Biliary duct.common:Document:XR.fluor
C0881810|BDs+GB RI for Bil Pat W Tc99mIV
C0881810|Biliary ducts and Gallbladder Scan for patency of biliary structures W Tc-99m IV
C0881810|Views for patency of biliary structures^W Tc-99m IV:Find:Pt:Biliary ducts+Gallbladder:Doc:Radnuc
C0881810|Views for patency of biliary structures^W Tc-99m Intravenous:Finding:Point in time:Biliary ducts+Gallbladder:Document:Radnuc
C0881826|Brain MRI W contr IV
C0881826|Brain MRI W contrast IV
C0881826|Multisection^W contrast IV:Find:Pt:Brain:Doc:MRI
C0881826|Multisection^W contrast Intravenous:Finding:Point in time:Brain:Document:MRI
C0881894|Views^W water soluble contrast Rectal:Finding:Point in time:Colon:Narrative:XR.fluor
C0881894|Colon Fluoroscopy W water soluble contrast PR
C0881894|Colon Flr W H2O sol contr PR
C0881894|Views^W water soluble contrast PR:Find:Pt:Colon:Doc:XR.fluor
C0881894|Views^W water soluble contrast Rectal:Finding:Point in time:Colon:Document:XR.fluor
C0881909|Extracranial vessels Fluoroscopic angiogram Embolectomy W contrast IA
C0881909|Embolectomy^W contrast IA:Find:Pt:Extracranial vessels:Doc:XR.fluor.angio
C0881909|EC vess XRA Embolectomy W contr IA
C0881909|Embolectomy^W contrast Intra-arterial:Finding:Point in time:Extracranial vessels:Document:XR.fluor.angio
C0882529|Extr CT
C0882529|Extremity CT
C0882529|Multisection:Finding:Point in time:Extremity:Document:Computerized Tomography
C0882529|Multisection:Find:Pt:Extremity:Doc:CT
C0882002|Multisection^WO & W contrast IV:Find:Pt:Knee:Doc:MRI
C0882002|Multisection^WO & W contrast Intravenous:Finding:Point in time:Knee:Document:MRI
C0882002|Knee MRI WO+W contr IV
C0882002|Knee MRI WO and W contrast IV
C1114502|Ft MRI WO contr
C1114502|Foot MRI WO contrast
C1114502|Multisection^WO contrast:Find:Pt:Foot:Doc:MRI
C1114502|Multisection^WO contrast:Finding:Point in time:Foot:Document:MRI
C1114507|Hip MRI WO contrast
C1114507|Hip MRI WO contr
C1114507|Multisection^WO contrast:Find:Pt:Hip:Doc:MRI
C1114507|Multisection^WO contrast:Finding:Point in time:Hip:Document:MRI
C1114509|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper arm:Document:MRI
C1114509|Upper arm MRI WO+W contr IV
C1114509|Multisection^WO & W contrast IV:Find:Pt:Upper arm:Doc:MRI
C1114509|Upper arm MRI WO and W contrast IV
C1114520|Abd US Ltd
C1114520|Abdomen US limited
C1114520|Multisection limited:Find:Pt:Abdomen:Doc:US
C1114520|Multisection limited:Finding:Point in time:Abdomen:Document:Ultrasound
C1114554|Chest XR PA+Lat+Lordotic Upr
C1114554|Chest X-ray PA and lateral and lordotic upright
C1114554|Views PA & lateral & lordotic upright:Find:Pt:Chest:Doc:XR
C1114554|Views PA & lateral & lordotic upright:Finding:Point in time:Chest:Document:XR
C1114575|Pelvis+Hip-Bl XR Max abd
C1114575|Pelvis and Hip - bilateral X-ray max abduction
C1114575|Views max abduction:Finding:Point in time:Pelvis+Hip.bilateral:Document:XR
C1114575|Views max abduction:Find:Pt:Pelvis+Hip.bilateral:Doc:XR
C1114603|VIEWS^W CONTRAST.XXX INTRAVENOUS:FINDING:POINT IN TIME:KIDNEY.BILATERAL AND COLLECTING SYSTEM:NARRATIVE:XR.TOMO
C1114603|Deprecated Kidney Bilateral & Collecting system X-ray tomograph Multisection W contrast IV
C1114603|Views^W contrast.XXX IV:Find:Pt:Kidney.bilateral+Collecting system:Nar:XR.tomo
C1114603|Deprecated KD-Bl+CS XR.Tomo
C1114603|Views^W contrast.XXX Intravenous:Finding:Point in time:Kidney.bilateral+Collecting system:Narrative:XR.tomo
C1114457|Head Cistern Fluoroscopy video W contrast
C1114457|Head.cistern XRVideo W contr
C1114457|Views^W contrast:Find:Pt:Head.cistern:Doc:XR.fluor.video
C1114457|Views^W contrast:Finding:Point in time:Head.cistern:Document:XR.fluor.video
C1114469|Fluoroscopy Guidance for change of tube in Sinus tract-- W contrast
C1114469|Sinus tr Flr Tube chnge guid W contr
C1114469|Guidance for change of tube^W contrast:Find:Pt:Sinus tract:Doc:XR.fluor
C1114469|Guidance for change of tube^W contrast:Finding:Point in time:Sinus tract:Document:XR.fluor
C1526828|Views^W contrast via nephrostomy tube:Find:Pt:Kidney.left:Doc:XR.fluor
C1526828|Kidney-L Flr W contr via NT
C1526828|Views^W contrast via nephrostomy tube:Finding:Point in time:Kidney.left:Document:XR.fluor
C1526828|Kidney - left Fluoroscopy W contrast via nephrostomy tube
C1543425|L-spine XR Lat Stand+W FE
C1543425|Views lateral^standing & W flexion & W extension:Finding:Point in time:Spine.lumbar:Document:XR
C1543425|Views lateral^standing & W flexion & W extension:Find:Pt:Spine.lumbar:Doc:XR
C1543425|Lumbar spine X-ray lateral standing and W flexion and W extension
C1543430|Knee-L XR Sunrise+Tunnel stand
C1543430|Knee - left X-ray Sunrise and tunnel standing
C1543430|Views Sunrise & tunnel^standing:Find:Pt:Knee.left:Doc:XR
C1543430|Views Sunrise & tunnel^standing:Finding:Point in time:Knee.left:Document:XR
C1543432|Should-L XR AP(w IR)+West Point
C1543432|Shoulder - left X-ray AP (W internal rotation) and West Point
C1543432|Views AP (W internal rotation) & West Point:Find:Pt:Shoulder.left:Doc:XR
C1543432|Views AP (W internal rotation) & West Point:Finding:Point in time:Shoulder.left:Document:XR
C1543445|Liver Flr Abscess drain guid
C1543445|Fluoroscopy Guidance for drainage of abscess of Liver
C1543445|Guidance for drainage of abscess:Find:Pt:Liver:Doc:XR.fluor
C1543445|Guidance for drainage of abscess:Finding:Point in time:Liver:Document:XR.fluor
C1543464|Knee - right X-ray 4 views and AP standing
C1543464|Knee-R XR 4V+AP stand
C1543464|Views 4 & AP^standing:Finding:Point in time:Knee.right:Document:XR
C1543464|Views 4 & AP^standing:Find:Pt:Knee.right:Doc:XR
C1543805|RI Tum local guid W RNC IV
C1543805|Scan Guidance for localization of tumor
C1543805|Guidance for localization of tumor^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543805|Guidance for localization of tumor^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C1543806|Vein RI W Tc99mSC IV
C1543806|Vein Scan W Tc-99m SC IV
C1543806|Views^W Tc-99m Subcutaneous Intravenous:Finding:Point in time:Vein:Document:Radnuc
C1543806|Views^W Tc-99m SC IV:Find:Pt:Vein:Doc:Radnuc
C1543808|Vein RI W Tc99mHDP IV
C1543808|Vein Scan W Tc-99m HDP IV
C1543808|Views^W Tc-99m HDP IV:Find:Pt:Vein:Doc:Radnuc
C1543808|Views^W Tc-99m HDP Intravenous:Finding:Point in time:Vein:Document:Radnuc
C1543883|Views static^W radionuclide Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1543883|Views static^W radionuclide IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1543883|Kidney - bilateral Scan static
C1543883|Kdny-Bl RI Static W RNC IV
C1542920|LV RI FP W RNC IV
C1542920|Left ventricle Scan first pass
C1542920|Views first pass^W radionuclide Intravenous:Finding:Point in time:Heart.ventricle.left:Document:Radnuc
C1542920|Views first pass^W radionuclide IV:Find:Pt:Heart.ventricle.left:Doc:Radnuc
C1543912|Hrt RI FP+WM W RNC IV
C1543912|Heart Scan first pass and wall motion
C1543912|Views first pass & wall motion^W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543912|Views first pass & wall motion^W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543950|Hrt RI Gated W Stress+W RNC IV
C1543950|Heart Scan gated W stress and W radionuclide IV
C1543950|Views gated^W stress & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1543950|Views gated^W stress & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543512|Renal ves DOP Ltd
C1543512|Renal vessels US.doppler limited
C1543512|Multisection limited:Find:Pt:Renal vessels:Doc:US.doppler
C1543512|Multisection limited:Finding:Point in time:Renal vessels:Document:Ultrasound.doppler
C1543147|XXX CT Needle local guid
C1543147|CT Guidance for needle localization of Unspecified body region
C1543147|Guidance for needle localization:Find:Pt:XXX:Doc:CT
C1543147|Guidance for needle localization:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1543565|Ribs lower post XR
C1543565|Ribs lower posterior X-ray
C1543565|Views:Finding:Point in time:Ribs.lower.posterior:Document:XR
C1543565|Views:Find:Pt:Ribs.lower.posterior:Doc:XR
C1526355|Deprecated Heel DXA T-score BDM
C1526355|Bone density:T Score:Point in time:Calcaneus:Quantitative:XR.DXA
C1526355|Bone density:Tscore:Pt:Calcaneus:Qn:XR.DXA
C1526355|Deprecated Calcaneus DXA [T-score] Bone density
C1543169|Scapula X-ray AP single view
C1543169|Scapula XR AP 1V
C1543169|View AP:Finding:Point in time:Scapula:Document:XR
C1543169|View AP:Find:Pt:Scapula:Doc:XR
C1543584|Umbilical vessels US.doppler
C1543584|Umb ves DOP
C1543584|Multisection:Find:Pt:Umbilical vessels:Doc:US.doppler
C1543584|Multisection:Finding:Point in time:Umbilical vessels:Document:Ultrasound.doppler
C1543594|Skull XR PA+R-Lat+L-Lat
C1543594|Skull X-ray PA and right lateral and left lateral
C1543594|Views PA & R-lateral & L-lateral:Finding:Point in time:Skull:Document:XR
C1543594|Views PA & R-lateral & L-lateral:Find:Pt:Skull:Doc:XR
C1543596|Skull XR PA+R-Lat+L-Lat+Caldwell+Towne
C1543596|Skull X-ray PA and right lateral and left lateral and Caldwell and Towne
C1543596|Views PA & R-lateral & L-lateral & Caldwell & Towne:Find:Pt:Skull:Doc:XR
C1543596|Views PA & R-lateral & L-lateral & Caldwell & Towne:Finding:Point in time:Skull:Document:XR
C1525167|Pelvis+Hip-R XR
C1525167|Pelvis and Hip - right X-ray
C1525167|Views:Find:Pt:Pelvis+Hip.right:Doc:XR
C1525167|Views:Finding:Point in time:Pelvis+Hip.right:Document:XR
C1525929|Deprecated Heel-R XR Harris
C1525929|View Harris:Finding:Point in time:Calcaneus.right:Document:XR
C1525929|View Harris:Find:Pt:Calcaneus.right:Doc:XR
C1525929|Deprecated Calcaneus - right X-ray Harris
C1542863|Breast FFD mammogram diagnostic
C1542863|Brst FFDM Dx
C1542863|Views diagnostic:Find:Pt:Breast:Doc:Mam.FFD
C1542863|Views diagnostic:Finding:Point in time:Breast:Document:Mam.FFD
C1543694|Brain SPECT
C1543694|Brain SPECT W RNC IV
C1543694|Multisection^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc.SPECT
C1543694|Multisection^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc.SPECT
C1526749|Should-R XR Grashey+Ax
C1526749|Shoulder - right X-ray Grashey and axillary
C1526749|Views Grashey & axillary:Find:Pt:Shoulder.right:Doc:XR
C1526749|Views Grashey & axillary:Finding:Point in time:Shoulder.right:Document:XR
C1526791|Temporal bone-L CT W contr IV
C1526791|Temporal bone - left CT W contrast IV
C1526791|Multisection^W contrast IV:Find:Pt:Temporal bone.left:Doc:CT
C1526791|Multisection^W contrast Intravenous:Finding:Point in time:Temporal bone.left:Document:Computerized Tomography
C1543412|Ribs-L+Chest XR
C1543412|Ribs - left and Chest X-ray
C1543412|Views:Finding:Point in time:Ribs.left+Chest:Document:XR
C1543412|Views:Find:Pt:Ribs.left+Chest:Doc:XR
C1543413|Should-L XR AP(w IR+ER)
C1543413|Shoulder - left X-ray AP (W internal rotation and W external rotation)
C1543413|Views AP (W internal rotation & W external rotation):Find:Pt:Shoulder.left:Doc:XR
C1543413|Views AP (W internal rotation & W external rotation):Finding:Point in time:Shoulder.left:Document:XR
C1543416|Ft-Bl XR AP+Lat stand
C1543416|Foot - bilateral X-ray AP and lateral standing
C1543416|Views AP & lateral^standing:Find:Pt:Foot.bilateral:Doc:XR
C1543416|Views AP & lateral^standing:Finding:Point in time:Foot.bilateral:Document:XR
C1543419|Ft-L XR AP+Lat+Obl stand
C1543419|Foot - left X-ray AP and lateral and oblique standing
C1543419|Views AP & lateral & oblique^standing:Finding:Point in time:Foot.left:Document:XR
C1543419|Views AP & lateral & oblique^standing:Find:Pt:Foot.left:Doc:XR
C1524428|Knee - left CT
C1524428|Knee-L CT
C1524428|Multisection:Find:Pt:Knee.left:Doc:CT
C1524428|Multisection:Finding:Point in time:Knee.left:Document:Computerized Tomography
C1524179|Shoulder - left X-ray tomograph
C1524179|Should-L XRTomo
C1524179|Multisection:Finding:Point in time:Shoulder.left:Document:XR.tomo
C1524179|Multisection:Find:Pt:Shoulder.left:Doc:XR.tomo
C1524821|Brst MRI WO contr
C1524821|Breast MRI WO contrast
C1524821|Multisection^WO contrast:Finding:Point in time:Breast:Document:MRI
C1524821|Multisection^WO contrast:Find:Pt:Breast:Doc:MRI
C1524446|Heart MRI limited
C1524446|Hrt MRI Ltd
C1524446|Multisection limited:Finding:Point in time:Heart:Document:MRI
C1524446|Multisection limited:Find:Pt:Heart:Doc:MRI
C1524455|L-spine MRI Ltd W contr IV
C1524455|Multisection limited^W contrast IV:Find:Pt:Spine.lumbar:Doc:MRI
C1524455|Multisection limited^W contrast Intravenous:Finding:Point in time:Spine.lumbar:Document:MRI
C1524455|Lumbar spine MRI limited W contrast IV
C1525296|Should-L XR Ax
C1525296|Shoulder - left X-ray axillary
C1525296|View axillary:Finding:Point in time:Shoulder.left:Document:XR
C1525296|View axillary:Find:Pt:Shoulder.left:Doc:XR
C1525237|Pelvis vessels MRI angiogram WO and W contrast IV
C1525237|Multisection^WO & W contrast IV:Find:Pt:Pelvis vessels:Doc:MRI.angio
C1525237|Multisection^WO & W contrast Intravenous:Finding:Point in time:Pelvis vessels:Document:MRI.angio
C1525237|Pelvis ves MRI.Angio WO+W contr IV
C1525252|Ankle ves MRI.Angio WO contr
C1525252|Ankle vessels MRI angiogram WO contrast
C1525252|Multisection^WO contrast:Find:Pt:Ankle vessels:Doc:MRI.angio
C1525252|Multisection^WO contrast:Finding:Point in time:Ankle vessels:Document:MRI.angio
C1525278|L-spine XR 2V stand
C1525278|Views 2^standing:Finding:Point in time:Spine.lumbar:Document:XR
C1525278|Views 2^standing:Find:Pt:Spine.lumbar:Doc:XR
C1525278|Lumbar spine X-ray 2 views standing
C1525279|Foot - bilateral X-ray 3 views standing
C1525279|Ft-Bl XR 3V stand
C1525279|Views 3^standing:Finding:Point in time:Foot.bilateral:Document:XR
C1525279|Views 3^standing:Find:Pt:Foot.bilateral:Doc:XR
C1524686|Knee X-ray Rosenberg standing
C1524686|Knee XR Rosenberg stand
C1524686|View Rosenberg^standing:Find:Pt:Knee:Doc:XR
C1524686|View Rosenberg^standing:Finding:Point in time:Knee:Document:XR
C1525459|Humerus - bilateral X-ray transthoracic
C1525459|Humerus-Bl XR Transthoracic
C1525459|View transthoracic:Finding:Point in time:Humerus.bilateral:Document:XR
C1525459|View transthoracic:Find:Pt:Humerus.bilateral:Doc:XR
C1524225|Shoulder - bilateral X-ray West Point
C1524225|Should-Bl XR West Point
C1524225|View West Point:Finding:Point in time:Shoulder.bilateral:Document:XR
C1524225|View West Point:Find:Pt:Shoulder.bilateral:Doc:XR
C1524250|Knee-Bl XR AP+Lat+Obl+Sunrise
C1524250|Knee - bilateral X-ray AP and lateral and oblique and Sunrise
C1524250|Views AP & lateral & oblique & Sunrise:Find:Pt:Knee.bilateral:Doc:XR
C1524250|Views AP & lateral & oblique & Sunrise:Finding:Point in time:Knee.bilateral:Document:XR
C1525529|Deprecated Views AP & axillary & Y:Finding:Point in time:Shoulder.left:Narrative:XR
C1525529|Views AP & axillary & Y:Find:Pt:Shoulder.left:Nar:XR
C1525529|Deprecated Shoulder Left X-ray AP & axillary & Y
C1525529|Deprecated Should-L XR AP+Ax+Y
C1525529|Views AP & axillary & Y:Finding:Point in time:Shoulder.left:Narrative:XR
C1525585|Elbow - left Fluoroscopy W contrast IS
C1525585|Views^W contrast IS:Find:Pt:Elbow.left:Doc:XR.fluor
C1525585|Elbow-L Flr W contr IS
C1525585|Views^W contrast Intrasynovial:Finding:Point in time:Elbow.left:Document:XR.fluor
C1525653|Multisection^WO & W contrast Intravenous:Finding:Point in time:Temporomandibular joint:Document:Computerized Tomography
C1525653|Temporomandibular joint CT WO and W contrast IV
C1525653|Multisection^WO & W contrast IV:Find:Pt:Temporomandibular joint:Doc:CT
C1525653|TMJ CT WO+W contr IV
C1525672|Multisection & 3D reconstruction:Finding:Point in time:Head:Document:Computerized Tomography
C1525672|Deprecated Head CT +3DR
C1525672|Deprecated Head CT and 3D reconstruction
C1525672|Multisection & 3D reconstruction:Find:Pt:Head:Doc:CT
C1525722|UE aa-Bl XRA W contr IA
C1525722|Upper extremity arteries - bilateral Fluoroscopic angiogram W contrast IA
C1525722|Views^W contrast IA:Find:Pt:Upper extremity arteries.bilateral:Doc:XR.fluor.angio
C1525722|Views^W contrast Intra-arterial:Finding:Point in time:Upper extremity arteries.bilateral:Document:XR.fluor.angio
C1525745|Renal v-L XRA W contr IV
C1525745|Renal vein - left Fluoroscopic angiogram W contrast IV
C1525745|Views^W contrast Intravenous:Finding:Point in time:Renal vein.left:Document:XR.fluor.angio
C1525745|Views^W contrast IV:Find:Pt:Renal vein.left:Doc:XR.fluor.angio
C1524696|Wrist-L CT W contr IV
C1524696|Wrist - left CT W contrast IV
C1524696|Multisection^W contrast IV:Find:Pt:Wrist.left:Doc:CT
C1524696|Multisection^W contrast Intravenous:Finding:Point in time:Wrist.left:Document:Computerized Tomography
C1525784|Knee XR PA V1 Stand+W 45 deg Flx
C1525784|Knee X-ray PA standing and W 45 degree flexion
C1525784|View PA^standing & W 45 degree flexion:Finding:Point in time:Knee:Document:XR
C1525784|View PA^standing & W 45 degree flexion:Find:Pt:Knee:Doc:XR
C1524136|Ac arch+Carot a.ext-R XRA W contr IA
C1524136|Aortic arch and Carotid artery.external - right Fluoroscopic angiogram W contrast IA
C1524136|Views^W contrast Intra-arterial:Finding:Point in time:Aortic arch+Carotid artery.external.right:Document:XR.fluor.angio
C1524136|Views^W contrast IA:Find:Pt:Aortic arch+Carotid artery.external.right:Doc:XR.fluor.angio
C1524139|Lymph Abd+Pelvic-L Flr W contr IL
C1524139|Lymphatics abdominal and Lymphatics pelvic - left Fluoroscopy W contrast intra lymphatic
C1524139|Views^W contrast intra lymphatic:Find:Pt:Lymphatics.abdominal+Lymphatics.pelvic.left:Doc:XR.fluor
C1524139|Views^W contrast intra lymphatic:Finding:Point in time:Lymphatics.abdominal+Lymphatics.pelvic.left:Document:XR.fluor
C1525945|Pelvis XR Inlet+Outlet+Obl
C1525945|Pelvis X-ray inlet and outlet and oblique
C1525945|Views inlet & outlet & oblique:Find:Pt:Pelvis:Doc:XR
C1525945|Views inlet & outlet & oblique:Finding:Point in time:Pelvis:Document:XR
C1525838|Brst Mam Mag
C1525838|Breast Mammogram magnification
C1525838|Views magnification:Find:Pt:Breast:Doc:Mam
C1525838|Views magnification:Finding:Point in time:Breast:Document:Mam
C1525955|Extr XR
C1525955|Extremity X-ray
C1525955|Views:Find:Pt:Extremity:Doc:XR
C1525955|Views:Finding:Point in time:Extremity:Document:XR
C1525958|Views^W contrast Intrasynovial:Finding:Point in time:Wrist.right:Document:XR.fluor
C1525958|Views^W contrast IS:Find:Pt:Wrist.right:Doc:XR.fluor
C1525958|Wrist-R Flr W contr IS
C1525958|Wrist - right Fluoroscopy W contrast IS
C1525985|Ankle - right X-ray lateral W manual stress
C1525985|Ankle-R XR Lat W Stress
C1525985|Views lateral^W manual stress:Find:Pt:Ankle.right:Doc:XR
C1525985|Views lateral^W manual stress:Finding:Point in time:Ankle.right:Document:XR
C1526019|Ft-R XR Lat
C1526019|Foot - right X-ray lateral
C1526019|View lateral:Find:Pt:Foot.right:Doc:XR
C1526019|View lateral:Finding:Point in time:Foot.right:Document:XR
C1526129|UE vv-R XRA W contr IV
C1526129|Upper extremity veins - right Fluoroscopic angiogram W contrast IV
C1526129|Views^W contrast IV:Find:Pt:Upper extremity veins.right:Doc:XR.fluor.angio
C1526129|Views^W contrast Intravenous:Finding:Point in time:Upper extremity veins.right:Document:XR.fluor.angio
C1525899|Wrist-R XR 5V
C1525899|Wrist - right X-ray 5 views
C1525899|Views 5:Find:Pt:Wrist.right:Doc:XR
C1525899|Views 5:Finding:Point in time:Wrist.right:Document:XR
C1526032|Hand-R XR
C1526032|Hand - right X-ray
C1526032|Views:Find:Pt:Hand.right:Doc:XR
C1526032|Views:Finding:Point in time:Hand.right:Document:XR
C1526154|Sinuses XR Lat+Waters
C1526154|Sinuses X-ray lateral and Waters
C1526154|Views lateral & Waters:Find:Pt:Sinuses:Doc:XR
C1526154|Views lateral & Waters:Finding:Point in time:Sinuses:Document:XR
C1524269|SC joint XR AP 1V
C1524269|Sternoclavicular Joint X-ray AP single view
C1524269|View AP:Find:Pt:Sternoclavicular joint:Doc:XR
C1524269|View AP:Finding:Point in time:Sternoclavicular joint:Document:XR
C1524704|Wrist X-ray 3 views
C1524704|Wrist XR 3V
C1524704|Views 3:Find:Pt:Wrist:Doc:XR
C1524704|Views 3:Finding:Point in time:Wrist:Document:XR
C1526282|Kidney - right US
C1526282|Kidney-R US
C1526282|Multisection:Find:Pt:Kidney.right:Doc:US
C1526282|Multisection:Finding:Point in time:Kidney.right:Document:Ultrasound
C1526295|Hip-L XR in Surg
C1526295|Hip - left X-ray during surgery
C1526295|View^during surgery:Find:Pt:Hip.left:Doc:XR
C1526295|View^during surgery:Finding:Point in time:Hip.left:Document:XR
C1525143|Penis US
C1525143|Multisection:Finding:Point in time:Penis:Document:Ultrasound
C1525143|Multisection:Find:Pt:Penis:Doc:US
C1524475|Multisection^W contrast IS:Find:Pt:Shoulder.right:Doc:CT
C1524475|Multisection^W contrast Intrasynovial:Finding:Point in time:Shoulder.right:Document:Computerized Tomography
C1524475|Shoulder - right CT W contrast IS
C1524475|Should-R CT W contr IS
C1524480|Ankle MRI W contr IV
C1524480|Ankle MRI W contrast IV
C1524480|Multisection^W contrast IV:Find:Pt:Ankle:Doc:MRI
C1524480|Multisection^W contrast Intravenous:Finding:Point in time:Ankle:Document:MRI
C1524874|Hip-R CT WO contr
C1524874|Hip - right CT WO contrast
C1524874|Multisection^WO contrast:Finding:Point in time:Hip.right:Document:Computerized Tomography
C1524874|Multisection^WO contrast:Find:Pt:Hip.right:Doc:CT
C1524875|Hip - right MRI WO contrast
C1524875|Hip-R MRI WO contr
C1524875|Multisection^WO contrast:Find:Pt:Hip.right:Doc:MRI
C1524875|Multisection^WO contrast:Finding:Point in time:Hip.right:Document:MRI
C1524890|Knee CT WO contrast
C1524890|Knee CT WO contr
C1524890|Multisection^WO contrast:Find:Pt:Knee:Doc:CT
C1524890|Multisection^WO contrast:Finding:Point in time:Knee:Document:Computerized Tomography
C1524166|Hip CT W contr IV
C1524166|Hip CT W contrast IV
C1524166|Multisection^W contrast IV:Find:Pt:Hip:Doc:CT
C1524166|Multisection^W contrast Intravenous:Finding:Point in time:Hip:Document:Computerized Tomography
C1524153|Sinuses CT WO contrast
C1524153|Sinuses CT WO contr
C1524153|Multisection^WO contrast:Finding:Point in time:Head>Sinuses:Document:Computerized Tomography
C1524153|Multisection^WO contrast:Find:Pt:Head>Sinuses:Doc:CT
C1524571|Pelvis MRI W contr IV
C1524571|Pelvis MRI W contrast IV
C1524571|Multisection^W contrast Intravenous:Finding:Point in time:Pelvis:Document:MRI
C1524571|Multisection^W contrast IV:Find:Pt:Pelvis:Doc:MRI
C1524930|Elbow X-ray Single view
C1524930|Elbow XR 1V
C1524930|View 1:Find:Pt:Elbow:Doc:XR
C1524930|View 1:Finding:Point in time:Elbow:Document:XR
C1524200|Wrist - left X-ray Single view
C1524200|Wrist-L XR 1V
C1524200|View 1:Find:Pt:Wrist.left:Doc:XR
C1524200|View 1:Finding:Point in time:Wrist.left:Document:XR
C1524624|Chest X-ray 3 views
C1524624|Chest XR 3V
C1524624|Views 3:Finding:Point in time:Chest:Document:XR
C1524624|Views 3:Find:Pt:Chest:Doc:XR
C1524642|Toes - left X-ray 3 views
C1524642|Toes-L XR 3V
C1524642|Views 3:Find:Pt:Toes.left:Doc:XR
C1524642|Views 3:Finding:Point in time:Toes.left:Document:XR
C1524643|Ankle X-ray 4 views
C1524643|Ankle XR 4V
C1524643|Views 4:Finding:Point in time:Ankle:Document:XR
C1524643|Views 4:Find:Pt:Ankle:Doc:XR
C1525009|L-spine XR 2V
C1525009|Views 2:Finding:Point in time:Spine.lumbar:Document:XR
C1525009|Views 2:Find:Pt:Spine.lumbar:Doc:XR
C1525009|Lumbar spine X-ray 2 views
C1524755|Upper arm-R CT WO+W contr IV
C1524755|Multisection^WO & W contrast IV:Find:Pt:Upper arm.right:Doc:CT
C1524755|Upper arm - right CT WO and W contrast IV
C1524755|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper arm.right:Document:Computerized Tomography
C1525047|Humerus-L XR AP+Lat
C1525047|Humerus - left X-ray AP and lateral
C1525047|Views AP & lateral:Finding:Point in time:Humerus.left:Document:XR
C1525047|Views AP & lateral:Find:Pt:Humerus.left:Doc:XR
C1525051|Patella-Bl XR AP+Lat
C1525051|Patella - bilateral X-ray AP and lateral
C1525051|Views AP & lateral:Find:Pt:Patella.bilateral:Doc:XR
C1525051|Views AP & lateral:Finding:Point in time:Patella.bilateral:Document:XR
C1525061|Elbow XR AP+Lat+Obl
C1525061|Elbow X-ray AP and lateral and oblique
C1525061|Views AP & lateral & oblique:Finding:Point in time:Elbow:Document:XR
C1525061|Views AP & lateral & oblique:Find:Pt:Elbow:Doc:XR
C1524411|Hip - right MRI
C1524411|Hip-R MRI
C1524411|Multisection:Find:Pt:Hip.right:Doc:MRI
C1524411|Multisection:Finding:Point in time:Hip.right:Document:MRI
C1524423|Kidney - left MRI
C1524423|Kidney-L MRI
C1524423|Multisection:Find:Pt:Kidney.left:Doc:MRI
C1524423|Multisection:Finding:Point in time:Kidney.left:Document:MRI
C1524424|Kidney-R MRI
C1524424|Kidney - right MRI
C1524424|Multisection:Finding:Point in time:Kidney.right:Document:MRI
C1524424|Multisection:Find:Pt:Kidney.right:Doc:MRI
C1524772|Multisection^WO & W contrast Intravenous:Finding:Point in time:Posterior fossa:Document:Computerized Tomography
C1524772|Posterior fossa CT WO and W contrast IV
C1524772|Multisection^WO & W contrast IV:Find:Pt:Posterior fossa:Doc:CT
C1524772|Post fossa CT WO+W contr IV
C1525093|Vessel Fluoroscopic angiogram Atherectomy W contrast
C1525093|Atherectomy^W contrast:Finding:Point in time:Vessel:Document:XR.fluor.angio
C1525093|Atherectomy^W contrast:Find:Pt:Vessel:Doc:XR.fluor.angio
C1525093|Vesl XRA Atherect W contr
C1830185|Mammogram Guidance for fine needle aspiration of Breast - left
C1830185|Brst-L Mam FNA Asp
C1830185|Guidance for aspiration.fine needle:Find:Pt:Breast.left:Doc:Mam
C1830185|Guidance for aspiration.fine needle:Finding:Point in time:Breast.left:Document:Mam
C1830207|Multisection^W contrast IV:Find:Pt:Whole body:Doc:CT
C1830207|Whole body CT W contr IV
C1830207|Whole body CT W contrast IV
C1830207|Multisection^W contrast Intravenous:Finding:Point in time:Whole body:Document:Computerized Tomography
C1830227|Maxillofacial region CT W reduced contrast volume IV
C1830227|Maxillofacial CT W red contr vol IV
C1830227|Multisection^W reduced contrast volume Intravenous:Finding:Point in time:Head>Maxillofacial region:Document:Computerized Tomography
C1830227|Multisection^W reduced contrast volume IV:Find:Pt:Head>Maxillofacial region:Doc:CT
C1830094|Breast Implant - unilateral Mammogram
C1830094|Brst implant-Ul Mam
C1830094|Views:Finding:Point in time:Breast implant.unilateral:Document:Mam
C1830094|Views:Find:Pt:Breast implant.unilateral:Doc:Mam
C1715411|Liver+Spleen RI W Tc99mMAA IV
C1715411|Liver and Spleen Scan W Tc-99m MAA IV
C1715411|Views^W Tc-99m MAA Intravenous:Finding:Point in time:Liver+Spleen:Document:Radnuc
C1715411|Views^W Tc-99m MAA IV:Find:Pt:Liver+Spleen:Doc:Radnuc
C1717313|Bone RI W Tc99mMedronate IV
C1717313|Bone Scan W Tc-99m medronate IV
C1717313|Views^W Tc-99m medronate IV:Find:Pt:Bone:Doc:Radnuc
C1717313|Views^W Tc-99m medronate Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1715454|Wrist X-ray GE 3 views
C1715454|Wrist XR GE 3V
C1715454|Views GE 3:Finding:Point in time:Wrist:Document:XR
C1715454|Views GE 3:Find:Pt:Wrist:Doc:XR
C1635663|Brain+Pituitary+ST MRI W contr IV
C1635663|Brain and Pituitary and Sella turcica MRI W contrast IV
C1635663|Multisection^W contrast IV:Find:Pt:Brain+Pituitary+Sella turcica:Doc:MRI
C1635663|Multisection^W contrast Intravenous:Finding:Point in time:Brain+Pituitary+Sella turcica:Document:MRI
C1632801|Brain and Pituitary and Sella turcica MRI WO and W contrast IV
C1632801|Brain+Pituitary+ST MRI WO+W contr IV
C1632801|Multisection^WO & W contrast IV:Find:Pt:Brain+Pituitary+Sella turcica:Doc:MRI
C1632801|Multisection^WO & W contrast Intravenous:Finding:Point in time:Brain+Pituitary+Sella turcica:Document:MRI
C1714901|Vessel Scan flow
C1714901|Views flow^W radionuclide Intravenous:Finding:Point in time:Vessel:Document:Radnuc
C1714901|Views flow^W radionuclide IV:Find:Pt:Vessel:Doc:Radnuc
C1714901|Vesl RI Flow W RNC IV
C1717260|XXX Flr Drain guid
C1717260|Fluoroscopy Guidance for drainage of Unspecified body region
C1717260|Guidance for drainage:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1717260|Guidance for drainage:Find:Pt:XXX:Doc:XR.fluor
C1714946|Liver+BDs+GB RI W RNC IV
C1714946|Liver and Biliary ducts and Gallbladder Scan
C1714946|Views^W radionuclide Intravenous:Finding:Point in time:Liver+Biliary ducts+Gallbladder:Document:Radnuc
C1714946|Views^W radionuclide IV:Find:Pt:Liver+Biliary ducts+Gallbladder:Doc:Radnuc
C1714961|UGI+SB Flr W Ba PO
C1714961|Upper Gastrointestine and Small bowel Fluoroscopy W barium contrast PO
C1714961|Views^W barium contrast PO:Find:Pt:Gastrointestine.upper+Small bowel:Doc:XR.fluor
C1714961|Views^W barium contrast Oral:Finding:Point in time:Gastrointestine.upper+Small bowel:Document:XR.fluor
C1715017|Brain RI Flow Ltd W RNC IV
C1715017|Brain Scan flow limited
C1715017|Views flow limited^W radionuclide Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1715017|Views flow limited^W radionuclide IV:Find:Pt:Brain:Doc:Radnuc
C1714495|Hrt RI PF Qn Rest+W RNC IV
C1714495|Heart Scan perfusion quantitative at rest and W radionuclide IV
C1714495|Views perfusion quantitative^at rest & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1714495|Views perfusion quantitative^at rest & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc
C1630769|Pelvis X-ray AP single view standing
C1630769|Pelvis XR AP 1V stand
C1630769|View AP^standing:Finding:Point in time:Pelvis:Document:XR
C1630769|View AP^standing:Find:Pt:Pelvis:Doc:XR
C1625791|Foot sesamoid bones - right X-ray
C1625791|Ft.sesamoids-R XR
C1625791|Views:Finding:Point in time:Foot.sesamoid bones.right:Document:XR
C1625791|Views:Find:Pt:Foot.sesamoid bones.right:Doc:XR
C1633398|Vein Fluoroscopic angiogram Percutaneous transluminal angioplasty of vessel W contrast IA
C1633398|Vein XRA PTA of ves W contr IA
C1633398|Percutaneous transluminal angioplasty of vessel^W contrast Intra-arterial:Finding:Point in time:Vein:Document:XR.fluor.angio
C1633398|Percutaneous transluminal angioplasty of vessel^W contrast IA:Find:Pt:Vein:Doc:XR.fluor.angio
C1646317|Pelvis XR Stereo
C1646317|Pelvis X-ray stereo
C1646317|View stereo:Find:Pt:Pelvis:Doc:XR
C1646317|View stereo:Finding:Point in time:Pelvis:Document:XR
C1641047|Uterus+FT US W saline IU
C1641047|Multisection^W saline Intrauterine:Finding:Point in time:Uterus+Fallopian tubes:Document:Ultrasound
C1641047|Multisection^W saline IU:Find:Pt:Uterus+Fallopian tubes:Doc:US
C1641047|Uterus and Fallopian tubes US W saline IU
C1627299|Pelvis+Hip-Bl XR AP+Lat Frog
C1627299|Pelvis and Hip - bilateral X-ray AP and lateral frog
C1627299|Views AP & lateral frog:Find:Pt:Pelvis+Hip.bilateral:Doc:XR
C1627299|Views AP & lateral frog:Finding:Point in time:Pelvis+Hip.bilateral:Document:XR
C1644659|Scan for lymphoma
C1644659|RI for Lymphoma W RNC IV
C1644659|Views for lymphoma^W radionuclide IV:Find:Pt:^Patient:Doc:Radnuc
C1644659|Views for lymphoma^W radionuclide Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1630175|CT Guidance for needle biopsy of Lymph node
C1630175|LN CT Bx needle guid
C1630175|Guidance for biopsy.needle:Find:Pt:Lymph node:Doc:CT
C1630175|Guidance for biopsy.needle:Finding:Point in time:Lymph node:Document:Computerized Tomography
C1633390|Guidance for nerve block:Find:Pt:Spine:Doc:CT
C1633390|Spine CT Nerve Block guid
C1633390|CT Guidance for nerve block of Spine
C1633390|Guidance for nerve block:Finding:Point in time:Spine:Document:Computerized Tomography
C1641529|Neck XR Lat Port
C1641529|Neck X-ray lateral portable
C1641529|View lateral portable:Finding:Point in time:Neck:Document:XR
C1641529|View lateral portable:Find:Pt:Neck:Doc:XR
C1646782|Humerus - right X-ray portable
C1646782|Humerus-R XR port
C1646782|Views portable:Find:Pt:Humerus.right:Doc:XR
C1646782|Views portable:Finding:Point in time:Humerus.right:Document:XR
C1625217|Lower leg-Bl MRI W contr IV
C1625217|Lower leg - bilateral MRI W contrast IV
C1625217|Multisection^W contrast IV:Find:Pt:Lower leg.bilateral:Doc:MRI
C1625217|Multisection^W contrast Intravenous:Finding:Point in time:Lower leg.bilateral:Document:MRI
C1978448|Ankle+Foot-L XR
C1978448|Ankle - left and Foot.left X-ray
C1978448|Views:Find:Pt:Ankle.left+Foot.left:Doc:XR
C1978448|Views:Finding:Point in time:Ankle.left+Foot.left:Document:XR
C1977260|Brst.duct-R Mam 1V W contr intra Dct
C1977260|Breast duct - right Mammogram Single view W contrast intra duct
C1977260|View 1^W contrast intra duct:Find:Pt:Breast.duct.right:Doc:Mam
C1977260|View 1^W contrast intra duct:Finding:Point in time:Breast.duct.right:Document:Mam
C1953984|Foot - right X-ray GE 3 views
C1953984|Ft-R XR GE 3V
C1953984|Views GE 3:Finding:Point in time:Foot.right:Document:XR
C1953984|Views GE 3:Find:Pt:Foot.right:Doc:XR
C3174371|Sagittal sinus vein - left Fluoroscopic angiogram W contrast IV
C3174371|SS v-L XRA W contr IV
C3174371|Views^W contrast Intravenous:Finding:Point in time:Sagittal sinus vein.left:Document:XR.fluor.angio
C3174371|Views^W contrast IV:Find:Pt:Sagittal sinus vein.left:Doc:XR.fluor.angio
C3169523|Renal artery - left Fluoroscopic angiogram W contrast IA
C3169523|Renal a-L XRA W contr IA
C3169523|Views^W contrast IA:Find:Pt:Renal artery.left:Doc:XR.fluor.angio
C3169523|Views^W contrast Intra-arterial:Finding:Point in time:Renal artery.left:Document:XR.fluor.angio
C3533906|Multisection diagnostic:Finding:Point in time:Breast.bilateral:Document:Mam.FFD.tomosynthesis
C3533906|Breast - bilateral FFD mammogram-tomosynthesis diagnostic
C3533906|Multisection diagnostic:Find:Pt:Breast.bilateral:Doc:Mam.FFD.tomosynthesis
C3533906|Brst-Bl FFDM-DBT Dx
C3533799|Abdomen and Pelvis MRI W contrast PO and WO contrast IV
C3533799|Abd+Pelvis MRI W contr PO+WO IV
C3533799|Multisection^W contrast PO+WO contrast IV:Find:Pt:Abdomen+Pelvis:Doc:MRI
C3533799|Multisection^W contrast Oral+WO contrast Intravenous:Finding:Point in time:Abdomen+Pelvis:Document:MRI
C3655082|Extr aa-Bl DOP Ltd+Phys stdy
C3655082|Multisection limited & physiologic artery study:Finding:Point in time:Extremity arteries.bilateral:Document:Ultrasound.doppler
C3655082|Extremity arteries - bilateral US.doppler Multisection limited and physiologic artery study
C3655082|Multisection limited & physiologic artery study:Find:Pt:Extremity arteries.bilateral:Doc:US.doppler
C3262958|Knee X-ray Sunrise and tunnel
C3262958|Knee XR Sunrise+Tunnel
C3262958|Views Sunrise & tunnel:Finding:Point in time:Knee:Document:XR
C3262958|Views Sunrise & tunnel:Find:Pt:Knee:Doc:XR
C3262960|Ankle - left X-ray 3 views standing
C3262960|Ankle-L XR 3V stand
C3262960|Views 3^standing:Find:Pt:Ankle.left:Doc:XR
C3262960|Views 3^standing:Finding:Point in time:Ankle.left:Document:XR
C3262990|Elbow-Bl MRI W contr IV
C3262990|Elbow - bilateral MRI W contrast IV
C3262990|Multisection^W contrast IV:Find:Pt:Elbow.bilateral:Doc:MRI
C3262990|Multisection^W contrast Intravenous:Finding:Point in time:Elbow.bilateral:Document:MRI
C3263043|Liver Scan W Tc-99m SC IV
C3263043|Liver RI W Tc99mSC IV
C3263043|Views^W Tc-99m Subcutaneous Intravenous:Finding:Point in time:Liver:Document:Radnuc
C3263043|Views^W Tc-99m SC IV:Find:Pt:Liver:Doc:Radnuc
C3263069|LE-R XR 2V
C3263069|Lower extremity - right X-ray 2 views
C3263069|Views 2:Finding:Point in time:Lower extremity.right:Document:XR
C3263069|Views 2:Find:Pt:Lower extremity.right:Doc:XR
C3261716|Chest US limited
C3261716|Chest US Ltd
C3261716|Multisection limited:Find:Pt:Chest:Doc:US
C3261716|Multisection limited:Finding:Point in time:Chest:Document:Ultrasound
C3263090|US Guidance for needle biopsy of Breast - right
C3263090|Brst-R US Bx needle guid
C3263090|Guidance for biopsy.needle:Finding:Point in time:Breast.right:Document:Ultrasound
C3263090|Guidance for biopsy.needle:Find:Pt:Breast.right:Doc:US
C3263091|Salivary gland US Bx needle guid
C3263091|US Guidance for needle biopsy of Salivary gland
C3263091|Guidance for biopsy.needle:Finding:Point in time:Salivary gland:Document:Ultrasound
C3263091|Guidance for biopsy.needle:Find:Pt:Salivary gland:Doc:US
C0942171|Thumb-L XR
C0942171|Thumb - left X-ray
C0942171|Views:Finding:Point in time:Thumb.left:Document:XR
C0942171|Views:Find:Pt:Thumb.left:Doc:XR
C0942261|Should-Bl MRI
C0942261|Shoulder - bilateral MRI
C0942261|Multisection:Find:Pt:Shoulder.bilateral:Doc:MRI
C0942261|Multisection:Finding:Point in time:Shoulder.bilateral:Document:MRI
C0942276|Wrist - right US
C0942276|Wrist-R US
C0942276|Multisection:Find:Pt:Wrist.right:Doc:US
C0942276|Multisection:Finding:Point in time:Wrist.right:Document:Ultrasound
C0945331|Brst-L US Ltd
C0945331|Breast - left US limited
C0945331|Multisection limited:Find:Pt:Breast.left:Doc:US
C0945331|Multisection limited:Finding:Point in time:Breast.left:Document:Ultrasound
C0942314|US Guidance for drainage of Extremity - right
C0942314|Extr-R US Drain guid
C0942314|Guidance for drainage:Finding:Point in time:Extremity.right:Document:Ultrasound
C0942314|Guidance for drainage:Find:Pt:Extremity.right:Doc:US
C0945340|Brst-Bl Mam Cyst Asp guid
C0945340|Mammogram Guidance for aspiration of cyst of Breast - bilateral
C0945340|Guidance for aspiration of cyst:Find:Pt:Breast.bilateral:Doc:Mam
C0945340|Guidance for aspiration of cyst:Finding:Point in time:Breast.bilateral:Document:Mam
C0942334|Breast - right Mammogram diagnostic limited
C0942334|Brst-R Mam Dx Ltd
C0942334|Views diagnostic limited:Find:Pt:Breast.right:Doc:Mam
C0942334|Views diagnostic limited:Finding:Point in time:Breast.right:Document:Mam
C0942339|View AP^standing:Finding:Point in time:Knee.bilateral:Narrative:XR
C0942339|Knee-Bl XR AP 1V stand
C0942339|Knee - bilateral X-ray AP single view standing
C0942339|View AP^standing:Find:Pt:Knee.bilateral:Doc:XR
C0942339|View AP^standing:Finding:Point in time:Knee.bilateral:Document:XR
C0942357|Administration of vasodilator into catheter of Vein - right
C0942357|Vein-R VD admin into cath
C0942357|Administration of vasodilator into catheter:Find:Pt:Vein.right:Doc
C0942357|Administration of vasodilator into catheter:Finding:Point in time:Vein.right:Document
C0882040|Optic foramen X-ray
C0882040|Optic foramen XR
C0882040|Views:Finding:Point in time:Optic foramen:Document:XR
C0882040|Views:Find:Pt:Optic foramen:Doc:XR
C0882087|Multisection^WO & W contrast IV:Find:Pt:Head>Pituitary+Sella turcica:Doc:CT
C0882087|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head>Pituitary+Sella turcica:Document:Computerized Tomography
C0882087|Pituitary and Sella turcica CT WO and W contrast IV
C0882087|Head Pit+Slla turc CT WO+W contr IV
C0882194|Unspecified body region Courtesy consultation
C0882194|XXX Courtesy consult
C0882194|Courtesy consultation.XXX:Find:Pt:XXX:Doc
C0882194|Courtesy consultation.XXX:Finding:Point in time:To be specified in another part of the message:Document
C0882216|XXX Flr 15M
C0882216|Unspecified body region Fluoroscopy 15 minutes
C0882216|View:Find:15M:XXX:Doc:XR.fluor
C0882216|View:Finding:15 minutes:To be specified in another part of the message:Document:XR.fluor
C0882225|Hep a XRA Cath plac guid W contr IA
C0882225|Fluoroscopic angiogram Guidance for placement of catheter in Hepatic artery-- W contrast IA
C0882225|Guidance for placement of catheter^W contrast Intra-arterial:Finding:Point in time:Hepatic artery:Document:XR.fluor.angio
C0882225|Guidance for placement of catheter^W contrast IA:Find:Pt:Hepatic artery:Doc:XR.fluor.angio
C0942098|Views^W contrast IS:Find:Pt:Shoulder.bilateral:Doc:XR.fluor
C0942098|Shoulder - bilateral Fluoroscopy W contrast IS
C0942098|Views^W contrast Intrasynovial:Finding:Point in time:Shoulder.bilateral:Document:XR.fluor
C0942098|Should-Bl Flr W contr IS
C0942104|Spinal artery - left Fluoroscopic angiogram W contrast IA
C0942104|Spinal a-L XRA W contr IA
C0942104|Views^W contrast IA:Find:Pt:Spinal artery.left:Doc:XR.fluor.angio
C0942104|Views^W contrast Intra-arterial:Finding:Point in time:Spinal artery.left:Document:XR.fluor.angio
C0942118|Ankle-L XR
C0942118|Ankle - left X-ray
C0942118|Views:Finding:Point in time:Ankle.left:Document:XR
C0942118|Views:Find:Pt:Ankle.left:Doc:XR
C0942124|Deprecated Carpal bones-L XR
C0942124|Views:Finding:Point in time:Carpal bones.left:Narrative:XR
C0942124|Deprecated Carpal bones - left X-ray
C0942124|Views:Find:Pt:Carpal bones.left:Nar:XR
C0881782|Anus US
C0881782|Multisection:Finding:Point in time:Anus:Document:Ultrasound
C0881782|Multisection:Find:Pt:Anus:Doc:US
C0881789|UE vv XRA W contr IV
C0881789|Upper extremity veins Fluoroscopic angiogram W contrast IV
C0881789|Views^W contrast Intravenous:Finding:Point in time:Upper extremity veins:Document:XR.fluor.angio
C0881789|Views^W contrast IV:Find:Pt:Upper extremity veins:Doc:XR.fluor.angio
C0881813|BDs+GB Flr W contr PC transhepatic
C0881813|Biliary ducts and Gallbladder Fluoroscopy W contrast percutaneous transhepatic
C0881813|Views^W contrast percutaneous transhepatic:Finding:Point in time:Biliary ducts+Gallbladder:Document:XR.fluor
C0881813|Views^W contrast percutaneous transhepatic:Find:Pt:Biliary ducts+Gallbladder:Doc:XR.fluor
C0882523|Chest X-ray AP left lateral-decubitus portable
C0882523|Chest XR AP L-Lat Decub Port
C0882523|View AP L-lateral-decubitus portable:Find:Pt:Chest:Doc:XR
C0882523|View AP L-lateral-decubitus portable:Finding:Point in time:Chest:Document:XR
C0881901|Views:Finding:Point in time:Elbow:Narrative:XR
C0881901|Elbow X-ray
C0881901|Elbow XR
C0881901|Views:Find:Pt:Elbow:Doc:XR
C0881901|Views:Finding:Point in time:Elbow:Document:XR
C0881982|Guidance for placement of percutaneous nephroureteral stent^W contrast via stent:Find:Pt:Kidney.bilateral:Doc:XR.fluor
C0881982|Guidance for placement of percutaneous nephroureteral stent^W contrast via stent:Finding:Point in time:Kidney.bilateral:Document:XR.fluor
C0881982|Fluoroscopy Guidance for placement of percutaneous nephroureteral stent in Kidney - bilateral-- W contrast via stent
C0881982|Kdny-Bl Flr PCNUS guid W contr via stnt
C0882001|Knee XR Merchants
C0882001|Knee X-ray Merchants
C0882001|View Merchants:Finding:Point in time:Knee:Document:XR
C0882001|View Merchants:Find:Pt:Knee:Doc:XR
C1114480|IAC MRI WO contr
C1114480|Internal auditory canal MRI WO contrast
C1114480|Multisection^WO contrast:Find:Pt:Internal auditory canal:Doc:MRI
C1114480|Multisection^WO contrast:Finding:Point in time:Internal auditory canal:Document:MRI
C1114491|Liver MRI WO contrast
C1114491|Liver MRI WO contr
C1114491|Multisection^WO contrast:Find:Pt:Liver:Doc:MRI
C1114491|Multisection^WO contrast:Finding:Point in time:Liver:Document:MRI
C1114493|Pelvis+Hip MRI WO contr
C1114493|Pelvis and Hip MRI WO contrast
C1114493|Multisection^WO contrast:Finding:Point in time:Pelvis+Hip:Document:MRI
C1114493|Multisection^WO contrast:Find:Pt:Pelvis+Hip:Doc:MRI
C1114537|View 1 portable:Finding:Point in time:Skull:Narrative:XR
C1114537|Skull X-ray Single view portable
C1114537|Skull XR 1V port
C1114537|View 1 portable:Find:Pt:Skull:Doc:XR
C1114537|View 1 portable:Finding:Point in time:Skull:Document:XR
C1114549|Chest XR W insp+exp
C1114549|Chest X-ray W inspiration and expiration
C1114549|Views^W inspiration & expiration:Finding:Point in time:Chest:Document:XR
C1114549|Views^W inspiration & expiration:Find:Pt:Chest:Doc:XR
C1114945|Pelvis+Hip XR
C1114945|Pelvis and Hip X-ray
C1114945|Views:Find:Pt:Pelvis+Hip:Doc:XR
C1114945|Views:Finding:Point in time:Pelvis+Hip:Document:XR
C1114591|Hip X-ray lateral frog
C1114591|Hip XR Lat Frog
C1114591|View lateral frog:Finding:Point in time:Hip:Document:XR
C1114591|View lateral frog:Find:Pt:Hip:Doc:XR
C1114643|Adrenal v-Bl XRA W contr IV
C1114643|Adrenal vein - bilateral Fluoroscopic angiogram W contrast IV
C1114643|Views^W contrast Intravenous:Finding:Point in time:Adrenal vein.bilateral:Document:XR.fluor.angio
C1114643|Views^W contrast IV:Find:Pt:Adrenal vein.bilateral:Doc:XR.fluor.angio
C1114643|VIEWS^W CONTRAST.XXX INTRAVENOUS:FINDING:POINT IN TIME:VEIN.ADRENAL.BILATERAL:NARRATIVE:XR.FLUOR.ANGIO
C1114653|C+T+L-spine MRI WO contr
C1114653|Spine Cervical and Thoracic and Lumbar MRI WO contrast
C1114653|Multisection^WO contrast:Finding:Point in time:Spine.cervical+Spine.thoracic+Spine.lumbar:Document:MRI
C1114653|Multisection^WO contrast:Find:Pt:Spine.cervical+Spine.thoracic+Spine.lumbar:Doc:MRI
C1114664|Renal ves MRI.Angio
C1114664|Renal vessels MRI angiogram
C1114664|Multisection:Finding:Point in time:Renal vessels:Document:MRI.angio
C1114664|Multisection:Find:Pt:Renal vessels:Doc:MRI.angio
C1114413|XXX CT RT guid W contr IV
C1114413|CT Guidance for radiation treatment of Unspecified body region-- W contrast IV
C1114413|Guidance for radiation treatment^W contrast IV:Find:Pt:XXX:Doc:CT
C1114413|Guidance for radiation treatment^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C1114419|Sinuses CT
C1114419|Multisection:Finding:Point in time:Head>Sinuses:Document:Computerized Tomography
C1114419|Multisection:Find:Pt:Head>Sinuses:Doc:CT
C1114429|Abd CT Bx guid
C1114429|CT Guidance for biopsy of Abdomen
C1114429|Guidance for biopsy:Find:Pt:Abdomen:Doc:CT
C1114429|Guidance for biopsy:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1114472|XXX Flr for Shunt
C1114472|Unspecified body region Fluoroscopy for shunt
C1114472|Views for shunt:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1114472|Views for shunt:Find:Pt:XXX:Doc:XR.fluor
C1543741|RI W Ga-67 IV
C1543741|Views^W Ga-67 IV:Find:Pt:^Patient:Doc:Radnuc
C1543741|Views^W Ga-67 Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543741|Scan W Ga-67 IV
C1543750|RI WB W I-131 mIBG IV
C1543750|Scan whole body W I-131 MIBG IV
C1543750|Views whole body^W I-131 MIBG IV:Find:Pt:^Patient:Doc:Radnuc
C1543750|Views whole body^W I-131 MIBG Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1543478|Should XR AP+Grashey+Ax
C1543478|Shoulder X-ray AP and Grashey and axillary
C1543478|Views AP & Grashey & axillary:Find:Pt:Shoulder:Doc:XR
C1543478|Views AP & Grashey & axillary:Finding:Point in time:Shoulder:Document:XR
C1543787|Hrt RI PF W ADE+Tl-201 IV
C1543787|Heart Scan perfusion W adenosine and W Tl-201 IV
C1543787|Views perfusion^W adenosine & W Tl-201 IV:Find:Pt:Heart:Doc:Radnuc
C1543787|Views perfusion^W adenosine & W Tl-201 Intravenous:Finding:Point in time:Heart:Document:Radnuc
C1543854|Bone RI W Tc99mHMPAO IV
C1543854|Bone Scan W Tc-99m HMPAO IV
C1543854|Views^W Tc-99m HMPAO IV:Find:Pt:Bone:Doc:Radnuc
C1543854|Views^W Tc-99m HMPAO Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543880|Views^W I-131 Intravenous:Finding:Point in time:Kidney.bilateral:Document:Radnuc
C1543880|Views^W I-131 IV:Find:Pt:Kidney.bilateral:Doc:Radnuc
C1543880|Kidney - bilateral Scan W I-131 IV
C1543880|Kdny-Bl RI W I-131 IV
C1543904|Bone RI 3 Phase WB W RNC IV
C1543904|Bone Scan 3 views phase whole body
C1543904|Views 3 phase whole body^W radionuclide Intravenous:Finding:Point in time:Bone:Document:Radnuc
C1543904|Views 3 phase whole body ^W radionuclide IV:Find:Pt:Bone:Doc:Radnuc
C1543501|Iliac artery US.doppler
C1543501|Iliac a DOP
C1543501|Multisection:Find:Pt:Iliac artery:Doc:US.doppler
C1543501|Multisection:Finding:Point in time:Iliac artery:Document:Ultrasound.doppler
C1543524|UE ves DOP
C1543524|Upper extremity vessels US.doppler
C1543524|Multisection:Finding:Point in time:Upper extremity vessels:Document:Ultrasound.doppler
C1543524|Multisection:Find:Pt:Upper extremity vessels:Doc:US.doppler
C1543155|Multisection^WO & W contrast IV:Find:Pt:Upper extremity:Doc:MRI
C1543155|UE MRI WO+W contr IV
C1543155|Multisection^WO & W contrast Intravenous:Finding:Point in time:Upper extremity:Document:MRI
C1543155|Upper extremity MRI WO and W contrast IV
C1543569|Ribs lower post-R XR
C1543569|Ribs lower posterior - right X-ray
C1543569|Views:Finding:Point in time:Ribs.lower.posterior.right:Document:XR
C1543569|Views:Find:Pt:Ribs.lower.posterior.right:Doc:XR
C1543166|Vein US limited
C1543166|Vein US Ltd
C1543166|Multisection limited:Finding:Point in time:Vein:Document:Ultrasound
C1543166|Multisection limited:Find:Pt:Vein:Doc:US
C1543194|Knee XR AP+Lat+R-Obl+L-Obl
C1543194|Knee X-ray AP and lateral and right oblique and left oblique
C1543194|Views AP & lateral & R-oblique & L-oblique:Finding:Point in time:Knee:Document:XR
C1543194|Views AP & lateral & R-oblique & L-oblique:Find:Pt:Knee:Doc:XR
C1543200|Hand XR PA+Obl
C1543200|Hand X-ray PA and oblique
C1543200|Views PA & oblique:Find:Pt:Hand:Doc:XR
C1543200|Views PA & oblique:Finding:Point in time:Hand:Document:XR
C1543593|Bones long X-ray survey limited
C1543593|Bones.long XR Survey Ltd
C1543593|Views survey limited:Find:Pt:Bones.long:Doc:XR
C1543593|Views survey limited:Finding:Point in time:Bones.long:Document:XR
C1543221|Ribs-R+Chest XR Lat+PA Chst
C1543221|Ribs - right and Chest X-ray lateral and PA chest
C1543221|Views lateral & PA chest:Find:Pt:Ribs.right+Chest:Doc:XR
C1543221|Views lateral & PA chest:Finding:Point in time:Ribs.right+Chest:Document:XR
C1543222|Ribs+Chest XR Lat+PA Chst
C1543222|Ribs and Chest X-ray lateral and PA chest
C1543222|Views lateral & PA chest:Finding:Point in time:Ribs+Chest:Document:XR
C1543222|Views lateral & PA chest:Find:Pt:Ribs+Chest:Doc:XR
C1525165|Lower extremity joint - right MRI limited WO contrast
C1525165|LE.joint-R MRI Ltd WO contr
C1525165|Multisection limited^WO contrast:Finding:Point in time:Lower extremity.joint.right:Document:MRI
C1525165|Multisection limited^WO contrast:Find:Pt:Lower extremity.joint.right:Doc:MRI
C1543266|Breast duct - left Mammogram W contrast intra multiple ducts
C1543266|Brst.duct-L Mam W contr intra Dcts
C1543266|Views^W contrast intra multiple ducts:Find:Pt:Breast.duct.left:Doc:Mam
C1543266|Views^W contrast intra multiple ducts:Finding:Point in time:Breast.duct.left:Document:Mam
C1543710|Hrt SPECT W DPY+RNC IV
C1543710|Heart SPECT W dipyridamole and W radionuclide IV
C1543710|Multisection^W dipyridamole & W radionuclide IV:Find:Pt:Heart:Doc:Radnuc.SPECT
C1543710|Multisection^W dipyridamole & W radionuclide Intravenous:Finding:Point in time:Heart:Document:Radnuc.SPECT
C1526789|Thoracic outlet - left MRI WO contrast
C1526789|TO-L MRI WO contr
C1526789|Multisection^WO contrast:Find:Pt:Thoracic outlet.left:Doc:MRI
C1526789|Multisection^WO contrast:Finding:Point in time:Thoracic outlet.left:Document:MRI
C1543379|LE MRI W contr IV
C1543379|Lower extremity MRI W contrast IV
C1543379|Multisection^W contrast IV:Find:Pt:Lower extremity:Doc:MRI
C1543379|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity:Document:MRI
C1543409|Abd XR R-Post Obl
C1543409|Abdomen X-ray right posterior oblique
C1543409|View R-posterior oblique:Find:Pt:Abdomen:Doc:XR
C1543409|View R-posterior oblique:Finding:Point in time:Abdomen:Document:XR
C2713302|Multisection:Finding:Point in time:Larynx:Narrative:MRI
C2713302|Larynx MRI
C2713302|Multisection:Finding:Point in time:Larynx:Document:MRI
C2713302|Multisection:Find:Pt:Larynx:Doc:MRI
C1525100|Kidney CT NT plac guid
C1525100|CT Guidance for placement of nephrostomy tube in Kidney
C1525100|Guidance for placement of nephrostomy tube:Finding:Point in time:Kidney:Document:Computerized Tomography
C1525100|Guidance for placement of nephrostomy tube:Find:Pt:Kidney:Doc:CT
C1524441|Abdomen CT limited
C1524441|Abd CT Ltd
C1524441|Multisection limited:Finding:Point in time:Abdomen:Document:Computerized Tomography
C1524441|Multisection limited:Find:Pt:Abdomen:Doc:CT
C1524239|L-spine CT Ltd WO contr
C1524239|Multisection limited^WO contrast:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C1524239|Multisection limited^WO contrast:Find:Pt:Spine.lumbar:Doc:CT
C1524239|Lumbar spine CT limited WO contrast
C1524241|T-spine MRI Ltd WO contr
C1524241|Multisection limited^WO contrast:Find:Pt:Spine.thoracic:Doc:MRI
C1524241|Multisection limited^WO contrast:Finding:Point in time:Spine.thoracic:Document:MRI
C1524241|Thoracic spine MRI limited WO contrast
C1524464|Hip MRI W contrast IS
C1524464|Hip MRI W contr IS
C1524464|Multisection^W contrast Intrasynovial:Finding:Point in time:Hip:Document:MRI
C1524464|Multisection^W contrast IS:Find:Pt:Hip:Doc:MRI
C1525292|Chest XR AP Upr port
C1525292|Chest X-ray AP upright portable
C1525292|View AP upright portable:Find:Pt:Chest:Doc:XR
C1525292|View AP upright portable:Finding:Point in time:Chest:Document:XR
C1525298|Hand - bilateral X-ray Brewerton
C1525298|Hand-Bl XR Brewerton
C1525298|View Brewerton:Finding:Point in time:Hand.bilateral:Document:XR
C1525298|View Brewerton:Find:Pt:Hand.bilateral:Doc:XR
C1525206|Multisection^W contrast IV:Find:Pt:Lower extremity>Vessels:Doc:CT.angio
C1525206|Lower extremity Vessels CT angiogram W contrast IV
C1525206|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity>Vessels:Document:Computerized Tomography.angio
C1525206|LE-ves CT.Angio W contr IV
C1525241|Temporal bone - left CT WO contrast
C1525241|Temporal bone-L CT WO contr
C1525241|Multisection^WO contrast:Finding:Point in time:Temporal bone.left:Document:Computerized Tomography
C1525241|Multisection^WO contrast:Find:Pt:Temporal bone.left:Doc:CT
C1525266|Multisection for calcium score:Finding:Point in time:Chest>Heart:Document:Computerized Tomography
C1525266|Multisection for calcium score:Find:Pt:Chest>Heart:Doc:CT
C1525266|Hrt CT for Calcium Score
C1525266|Heart CT for calcium scoring
C1525474|Humerus-Bl XR
C1525474|Humerus - bilateral X-ray
C1525474|Views:Finding:Point in time:Humerus.bilateral:Document:XR
C1525474|Views:Find:Pt:Humerus.bilateral:Doc:XR
C1525556|Should-L XR Grashey+Outlet
C1525556|Shoulder - left X-ray Grashey and outlet
C1525556|Views Grashey & outlet:Find:Pt:Shoulder.left:Doc:XR
C1525556|Views Grashey & outlet:Finding:Point in time:Shoulder.left:Document:XR
C1525564|Face XR Lat+Caldwell+Waters+SMV
C1525564|Facial bones X-ray lateral and Caldwell and Waters and submentovertex
C1525564|Views lateral & Caldwell & Waters & submentovertex:Finding:Point in time:Facial bones:Document:XR
C1525564|Views lateral & Caldwell & Waters & submentovertex:Find:Pt:Facial bones:Doc:XR
C1525618|Multisection:Finding:Point in time:Ankle+Foot:Narrative:MRI
C1525618|Ankle+Ft MRI
C1525618|Ankle and Foot MRI
C1525618|Multisection:Find:Pt:Ankle+Foot:Doc:MRI
C1525618|Multisection:Finding:Point in time:Ankle+Foot:Document:MRI
C1525635|Parotid gland MRI W contr IV
C1525635|Parotid gland MRI W contrast IV
C1525635|Multisection^W contrast Intravenous:Finding:Point in time:Parotid gland:Document:MRI
C1525635|Multisection^W contrast IV:Find:Pt:Parotid gland:Doc:MRI
C1525655|Temporomandibular joint - bilateral MRI WO and W contrast IV
C1525655|Multisection^WO & W contrast Intravenous:Finding:Point in time:Temporomandibular joint.bilateral:Document:MRI
C1525655|Multisection^WO & W contrast IV:Find:Pt:Temporomandibular joint.bilateral:Doc:MRI
C1525655|TMJ-Bl MRI WO+W contr IV
C1525667|TMJ-Bl MRI WO contr
C1525667|Temporomandibular joint - bilateral MRI WO contrast
C1525667|Multisection^WO contrast:Find:Pt:Temporomandibular joint.bilateral:Doc:MRI
C1525667|Multisection^WO contrast:Finding:Point in time:Temporomandibular joint.bilateral:Document:MRI
C1525681|Humerus bicipital groove X-ray
C1525681|Humerus bicipital groove XR
C1525681|Views:Find:Pt:Humerus.bicipital groove:Doc:XR
C1525681|Views:Finding:Point in time:Humerus.bicipital groove:Document:XR
C1525756|Brst MRI Dyn W contr IV
C1525756|Breast MRI dynamic W contrast IV
C1525756|Multisection dynamic^W contrast IV:Find:Pt:Breast:Doc:MRI
C1525756|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Breast:Document:MRI
C1525757|Deprecated Pituitary+ST CT Dyn W contr I
C1525757|Multisection dynamic^W contrast IV:Find:Pt:Head>Pituitary+Sella turcica:Doc:CT
C1525757|Multisection dynamic^W contrast Intravenous:Finding:Point in time:Head>Pituitary+Sella turcica:Document:Computerized Tomography
C1525757|Deprecated Pituitary and Sella turcica CT dynamic W contrast IV
C1524692|Wrist-R MRI W contr IS
C1524692|Multisection^W contrast IS:Find:Pt:Wrist.right:Doc:MRI
C1524692|Wrist - right MRI W contrast IS
C1524692|Multisection^W contrast Intrasynovial:Finding:Point in time:Wrist.right:Document:MRI
C1524698|Wrist-R CT W contr IV
C1524698|Wrist - right CT W contrast IV
C1524698|Multisection^W contrast Intravenous:Finding:Point in time:Wrist.right:Document:Computerized Tomography
C1524698|Multisection^W contrast IV:Find:Pt:Wrist.right:Doc:CT
C1525771|Wrist - left MRI WO contrast
C1525771|Wrist-L MRI WO contr
C1525771|Multisection^WO contrast:Find:Pt:Wrist.left:Doc:MRI
C1525771|Multisection^WO contrast:Finding:Point in time:Wrist.left:Document:MRI
C1525802|Multisection^W contrast Intravenous:Finding:Point in time:Head+Neck>Vessels:Document:Computerized Tomography.angio
C1525802|Multisection^W contrast IV:Find:Pt:Head+Neck>Vessels:Doc:CT.angio
C1525802|Head and Neck vessels CT angiogram W contrast IV
C1525802|Head+Neck Vess CT.Angio W contr IV
C1525816|Tib-Bl XR 10 Deg Cau Angle
C1525816|Tibia - bilateral X-ray 10 degree caudal angle
C1525816|View 10 degree caudal angle:Finding:Point in time:Tibia.bilateral:Document:XR
C1525816|View 10 degree caudal angle:Find:Pt:Tibia.bilateral:Doc:XR
C1525829|Toe fourth - left X-ray
C1525829|Toe 4th-L XR
C1525829|Views:Find:Pt:Toe.fourth.left:Doc:XR
C1525829|Views:Finding:Point in time:Toe.fourth.left:Document:XR
C1525836|Knee-Bl XR Holmblad stand
C1525836|Knee - bilateral X-ray Holmblad standing
C1525836|Views Holmblad^standing:Finding:Point in time:Knee.bilateral:Document:XR
C1525836|Views Holmblad^standing:Find:Pt:Knee.bilateral:Doc:XR
C1525949|Pelvis XR Outlet
C1525949|Pelvis X-ray outlet
C1525949|View outlet:Finding:Point in time:Pelvis:Document:XR
C1525949|View outlet:Find:Pt:Pelvis:Doc:XR
C1526120|Tib+Fib-R XR 2V
C1526120|Tibia - right and Fibula - right X-ray 2 views
C1526120|Views 2:Find:Pt:Tibia.right+Fibula.right:Doc:XR
C1526120|Views 2:Finding:Point in time:Tibia.right+Fibula.right:Document:XR
C1526123|Views^W contrast IS:Find:Pt:Temporomandibular joint.right:Doc:XR.fluor
C1526123|TMJ-R Flr W contr IS
C1526123|Temporomandibular joint - right Fluoroscopy W contrast IS
C1526123|Views^W contrast Intrasynovial:Finding:Point in time:Temporomandibular joint.right:Document:XR.fluor
C1526125|Toes - right X-ray 3 views
C1526125|Toes-R XR 3V
C1526125|Views 3:Find:Pt:Toes.right:Doc:XR
C1526125|Views 3:Finding:Point in time:Toes.right:Document:XR
C1525908|Deprecated Wrist-R XR 4V
C1525908|Views 4:Find:Pt:Wrist.right:Nar:XR
C1525908|Deprecated Wrist Right X-ray 4 views
C1525908|Views 4:Finding:Point in time:Wrist.right:Narrative:XR
C1525908|deprecated VIEWS 4:FINDING:POINT IN TIME:WRIST.RIGHT:NARRATIVE:XR
C1526060|Knee - right X-ray 5 views
C1526060|Knee-R XR 5V
C1526060|Views 5:Finding:Point in time:Knee.right:Document:XR
C1526060|Views 5:Find:Pt:Knee.right:Doc:XR
C1526068|Knee - right X-ray Rosenberg standing
C1526068|Knee-R XR Rosenberg stand
C1526068|View Rosenberg^standing:Finding:Point in time:Knee.right:Document:XR
C1526068|View Rosenberg^standing:Find:Pt:Knee.right:Doc:XR
C1526074|Knee-R XR
C1526074|Knee - right X-ray
C1526074|Views:Finding:Point in time:Knee.right:Document:XR
C1526074|Views:Find:Pt:Knee.right:Doc:XR
C1525126|Patella-R XR AP+Lat
C1525126|Patella - right X-ray AP and lateral
C1525126|Views AP & lateral:Find:Pt:Patella.right:Doc:XR
C1525126|Views AP & lateral:Finding:Point in time:Patella.right:Document:XR
C1525128|Popliteal a-R XRA W contr IA
C1525128|Popliteal artery - right Fluoroscopic angiogram W contrast IA
C1525128|Views^W contrast IA:Find:Pt:Popliteal artery.right:Doc:XR.fluor.angio
C1525128|Views^W contrast Intra-arterial:Finding:Point in time:Popliteal artery.right:Document:XR.fluor.angio
C1524276|Fluoroscopy Guidance for aspiration of Pleural space
C1524276|Pl space Flr Asp guid
C1524276|Guidance for aspiration:Finding:Point in time:Chest>Pleural space:Document:XR.fluor
C1524276|Guidance for aspiration:Find:Pt:Chest>Pleural space:Doc:XR.fluor
C1526202|Upper extremity X-ray 2 views
C1526202|UE XR 2V
C1526202|Views 2:Find:Pt:Upper extremity:Doc:XR
C1526202|Views 2:Finding:Point in time:Upper extremity:Document:XR
C1526220|Carotid artery.internal - right Fluoroscopic angiogram W contrast IA
C1526220|Carot a.Int-R XRA W contr IA
C1526220|Views^W contrast Intra-arterial:Finding:Point in time:Carotid artery.internal.right:Document:XR.fluor.angio
C1526220|Views^W contrast IA:Find:Pt:Carotid artery.internal.right:Doc:XR.fluor.angio
C1526243|Uterine a XRA W contr IA
C1526243|Uterine artery Fluoroscopic angiogram W contrast IA
C1526243|Views^W contrast IA:Find:Pt:Uterine artery:Doc:XR.fluor.angio
C1526243|Views^W contrast Intra-arterial:Finding:Point in time:Uterine artery:Document:XR.fluor.angio
C1524711|Head US limited
C1524711|Head US Ltd
C1524711|Multisection limited:Find:Pt:Head:Doc:US
C1524711|Multisection limited:Finding:Point in time:Head:Document:Ultrasound
C1526276|Mastoid US
C1526276|Multisection:Finding:Point in time:Mastoid:Document:Ultrasound
C1526276|Multisection:Find:Pt:Mastoid:Doc:US
C1526287|Visceral a US
C1526287|Visceral artery US
C1526287|Multisection:Finding:Point in time:Visceral artery:Document:Ultrasound
C1526287|Multisection:Find:Pt:Visceral artery:Doc:US
C1526290|Breast implant - right MRI
C1526290|Brst implant-R MRI
C1526290|Multisection:Finding:Point in time:Breast implant.right:Document:MRI
C1526290|Multisection:Find:Pt:Breast implant.right:Doc:MRI
C1526338|US Guidance for superficial aspiration.fine needle of Tissue
C1526338|Guidance for superficial aspiration.fine needle:Finding:Point in time:Tissue:Document:Ultrasound
C1526338|tiss US Sup FNA guid
C1526338|Guidance for superficial aspiration.fine needle:Find:Pt:Tissue:Doc:US
C1508082|Breast - bilateral Mammogram nipple profile
C1508082|Brst-Bl Mam Nipple Profile
C1508082|View nipple profile:Find:Pt:Breast.bilateral:Doc:Mam
C1508082|View nipple profile:Finding:Point in time:Breast.bilateral:Document:Mam
C1526315|Parotid gland-L Flr W contr intra SD
C1526315|Parotid gland - left Fluoroscopy W contrast intra salivary duct
C1526315|Views^W contrast intra salivary duct:Find:Pt:Parotid gland.left:Doc:XR.fluor
C1526315|Views^W contrast intra salivary duct:Finding:Point in time:Parotid gland.left:Document:XR.fluor
C1526316|Lacrimal duct - bilateral Fluoroscopy W contrast intra lacrimal duct
C1526316|Lacrimal duct-Bl Flr W contr intra LD
C1526316|Views^W contrast intra lacrimal duct:Find:Pt:Lacrimal duct.bilateral:Doc:XR.fluor
C1526316|Views^W contrast intra lacrimal duct:Finding:Point in time:Lacrimal duct.bilateral:Document:XR.fluor
C1524482|Ankle-L MRI W contr IV
C1524482|Ankle - left MRI W contrast IV
C1524482|Multisection^W contrast Intravenous:Finding:Point in time:Ankle.left:Document:MRI
C1524482|Multisection^W contrast IV:Find:Pt:Ankle.left:Doc:MRI
C1524498|Multisection^W contrast IV:Find:Pt:Calcaneus.right:Doc:CT
C1524498|Deprecated Heel-R CT W contr IV
C1524498|Multisection^W contrast Intravenous:Finding:Point in time:Calcaneus.right:Document:Computerized Tomography
C1524498|Deprecated Calcaneus - right CT W contrast IV
C1524893|Knee-L MRI WO contr
C1524893|Knee - left MRI WO contrast
C1524893|Multisection^WO contrast:Find:Pt:Knee.left:Doc:MRI
C1524893|Multisection^WO contrast:Finding:Point in time:Knee.left:Document:MRI
C1524517|Thigh MRI W contr IV
C1524517|Thigh MRI W contrast IV
C1524517|Multisection^W contrast IV:Find:Pt:Thigh:Doc:MRI
C1524517|Multisection^W contrast Intravenous:Finding:Point in time:Thigh:Document:MRI
C1524542|Upper arm MRI W contr IV
C1524542|Upper arm MRI W contrast IV
C1524542|Multisection^W contrast Intravenous:Finding:Point in time:Upper arm:Document:MRI
C1524542|Multisection^W contrast IV:Find:Pt:Upper arm:Doc:MRI
C1524543|Upper arm-L CT W contr IV
C1524543|Upper arm - left CT W contrast IV
C1524543|Multisection^W contrast Intravenous:Finding:Point in time:Upper arm.left:Document:Computerized Tomography
C1524543|Multisection^W contrast IV:Find:Pt:Upper arm.left:Doc:CT
C1524147|Scapula-L MRI WO contr
C1524147|Scapula - left MRI WO contrast
C1524147|Multisection^WO contrast:Find:Pt:Scapula.left:Doc:MRI
C1524147|Multisection^WO contrast:Finding:Point in time:Scapula.left:Document:MRI
C1524911|Scrotum+Test MRI WO contr
C1524911|Scrotum and Testicle MRI WO contrast
C1524911|Multisection^WO contrast:Find:Pt:Scrotum+Testicle:Doc:MRI
C1524911|Multisection^WO contrast:Finding:Point in time:Scrotum+Testicle:Document:MRI
C1524917|Lower leg - right MRI WO contrast
C1524917|Lower leg-R MRI WO contr
C1524917|Multisection^WO contrast:Find:Pt:Lower leg.right:Doc:MRI
C1524917|Multisection^WO contrast:Finding:Point in time:Lower leg.right:Document:MRI
C1524549|LE.joint-R MRI W contr IV
C1524549|Lower extremity joint - right MRI W contrast IV
C1524549|Multisection^W contrast IV:Find:Pt:Lower extremity.joint.right:Doc:MRI
C1524549|Multisection^W contrast Intravenous:Finding:Point in time:Lower extremity.joint.right:Document:MRI
C1524560|Knee-L MRI W contr IV
C1524560|Knee - left MRI W contrast IV
C1524560|Multisection^W contrast Intravenous:Finding:Point in time:Knee.left:Document:MRI
C1524560|Multisection^W contrast IV:Find:Pt:Knee.left:Doc:MRI
C1524196|Knee-Bl XR 1V
C1524196|Knee - bilateral X-ray Single view
C1524196|View 1:Finding:Point in time:Knee.bilateral:Document:XR
C1524196|View 1:Find:Pt:Knee.bilateral:Doc:XR
C1524939|Abdomen X-ray lateral
C1524939|Abd XR Lat
C1524939|View lateral:Find:Pt:Abdomen:Doc:XR
C1524939|View lateral:Finding:Point in time:Abdomen:Document:XR
C1524946|Foot - left X-ray lateral
C1524946|Ft-L XR Lat
C1524946|View lateral:Finding:Point in time:Foot.left:Document:XR
C1524946|View lateral:Find:Pt:Foot.left:Doc:XR
C1524281|IVC XRA Angpsty W contr IV
C1524281|Inferior vena cava Fluoroscopic angiogram Angioplasty W contrast IV
C1524281|Angioplasty^W contrast Intravenous:Finding:Point in time:Vena cava.inferior:Document:XR.fluor.angio
C1524281|Angioplasty^W contrast IV:Find:Pt:Vena cava.inferior:Doc:XR.fluor.angio
C1524606|Aorta abdominal MRI angiogram WO and W contrast IV
C1524606|Multisection^WO & W contrast IV:Find:Pt:Aorta.abdominal:Doc:MRI.angio
C1524606|Multisection^WO & W contrast Intravenous:Finding:Point in time:Aorta.abdominal:Document:MRI.angio
C1524606|Ab Ao MRI.Angio WO+W contr IV
C1524610|Breast MRI WO and W contrast IV
C1524610|Multisection^WO & W contrast IV:Find:Pt:Breast:Doc:MRI
C1524610|Brst MRI WO+W contr IV
C1524610|Multisection^WO & W contrast Intravenous:Finding:Point in time:Breast:Document:MRI
C1524987|Patella-L XR
C1524987|Patella - left X-ray
C1524987|Views:Find:Pt:Patella.left:Doc:XR
C1524987|Views:Finding:Point in time:Patella.left:Document:XR
C1524988|C-spine Flr
C1524988|Views:Find:Pt:Spine.cervical:Doc:XR.fluor
C1524988|Views:Finding:Point in time:Spine.cervical:Document:XR.fluor
C1524988|Cervical spine Fluoroscopy
C1524338|Ankle X-ray tomograph
C1524338|Ankle XRTomo
C1524338|Multisection:Find:Pt:Ankle:Doc:XR.tomo
C1524338|Multisection:Finding:Point in time:Ankle:Document:XR.tomo
C1526995|Ankle CT
C1526995|Multisection:Find:Pt:Ankle:Doc:CT
C1526995|Multisection:Finding:Point in time:Ankle:Document:Computerized Tomography
C1524653|Mandible X-ray 4 views
C1524653|Mandible XR 4V
C1524653|Views 4:Finding:Point in time:Mandible:Document:XR
C1524653|Views 4:Find:Pt:Mandible:Doc:XR
C1524654|Ribs - bilateral X-ray 4 views
C1524654|Ribs-Bl XR 4V
C1524654|Views 4:Finding:Point in time:Ribs.bilateral:Document:XR
C1524654|Views 4:Find:Pt:Ribs.bilateral:Doc:XR
C1524159|Deprecated Calcaneus X-ray 2 views
C1524159|Views 2:Finding:Point in time:Calcaneus:Document:XR
C1524159|Deprecated Heel XR 2V
C1524159|Views 2:Find:Pt:Calcaneus:Doc:XR
C1524162|Hip-L XR 2V
C1524162|Hip - left X-ray 2 views
C1524162|Views 2:Finding:Point in time:Hip.left:Document:XR
C1524162|Views 2:Find:Pt:Hip.left:Doc:XR
C1525011|Tib+Fib-L XR 2V
C1525011|Tibia - left and Fibula - left X-ray 2 views
C1525011|Views 2:Find:Pt:Tibia.left+Fibula.left:Doc:XR
C1525011|Views 2:Finding:Point in time:Tibia.left+Fibula.left:Document:XR
C1524351|IAC MRI
C1524351|Internal auditory canal MRI
C1524351|Multisection:Finding:Point in time:Internal auditory canal:Document:MRI
C1524351|Multisection:Find:Pt:Internal auditory canal:Doc:MRI
C1524380|Femur-Bl XRTomo
C1524380|Femur - bilateral X-ray tomograph
C1524380|Multisection:Find:Pt:Femur.bilateral:Doc:XR.tomo
C1524380|Multisection:Finding:Point in time:Femur.bilateral:Document:XR.tomo
C1524665|Multisection^WO & W contrast IV:Find:Pt:Femur.left:Doc:CT
C1524665|Femur - left CT WO and W contrast IV
C1524665|Multisection^WO & W contrast Intravenous:Finding:Point in time:Femur.left:Document:Computerized Tomography
C1524665|Femur-L CT WO+W contr IV
C1524746|Multisection^WO & W contrast IV:Find:Pt:Hip.bilateral:Doc:CT
C1524746|Hip - bilateral CT WO and W contrast IV
C1524746|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hip.bilateral:Document:Computerized Tomography
C1524746|Hip-Bl CT WO+W contr IV
C1524395|Hand-Bl CT
C1524395|Hand - bilateral CT
C1524395|Multisection:Find:Pt:Hand.bilateral:Doc:CT
C1524395|Multisection:Finding:Point in time:Hand.bilateral:Document:Computerized Tomography
C1524410|Hip-R CT
C1524410|Hip - right CT
C1524410|Multisection:Finding:Point in time:Hip.right:Document:Computerized Tomography
C1524410|Multisection:Find:Pt:Hip.right:Doc:CT
C1524793|Multisection^WO & W contrast IV:Find:Pt:Lower leg:Doc:CT
C1524793|Lower leg CT WO+W contr IV
C1524793|Lower leg CT WO and W contrast IV
C1524793|Multisection^WO & W contrast Intravenous:Finding:Point in time:Lower leg:Document:Computerized Tomography
C1524672|C-spine XR AP+Lat+Obl
C1524672|Views AP & lateral & oblique:Find:Pt:Spine.cervical:Doc:XR
C1524672|Views AP & lateral & oblique:Finding:Point in time:Spine.cervical:Document:XR
C1524672|Cervical spine X-ray AP and lateral and oblique
C1524677|Wrist - bilateral X-ray limited
C1524677|Wrist-Bl XR Ltd
C1524677|Views limited:Finding:Point in time:Wrist.bilateral:Document:XR
C1524677|Views limited:Find:Pt:Wrist.bilateral:Doc:XR
C1830206|Whole body CT
C1830206|Multisection:Finding:Point in time:Whole body:Document:Computerized Tomography
C1830206|Multisection:Find:Pt:Whole body:Doc:CT
C1715433|Kidney US Abscess drain guid
C1715433|US Guidance for drainage of abscess of Kidney
C1715433|Guidance for drainage of abscess:Finding:Point in time:Kidney:Document:Ultrasound
C1715433|Guidance for drainage of abscess:Find:Pt:Kidney:Doc:US
C1715439|Lower extremity vessels US.doppler
C1715439|LE ves DOP
C1715439|Multisection:Finding:Point in time:Lower extremity vessels:Document:Ultrasound.doppler
C1715439|Multisection:Find:Pt:Lower extremity vessels:Doc:US.doppler
C1715477|Fluoroscopy Guidance for fine needle aspiration of Kidney
C1715477|Kidney Flr FNA Asp
C1715477|Guidance for aspiration.fine needle:Finding:Point in time:Kidney:Document:XR.fluor
C1715477|Guidance for aspiration.fine needle:Find:Pt:Kidney:Doc:XR.fluor
C1717323|UE ves graft-Bl DOP Ltd
C1717323|Upper extremity vessel graft - bilateral US.doppler limited
C1717323|Multisection limited:Find:Pt:Upper extremity vessel graft.bilateral:Doc:US.doppler
C1717323|Multisection limited:Finding:Point in time:Upper extremity vessel graft.bilateral:Document:Ultrasound.doppler
C1644647|Femur-L XR port
C1644647|Femur - left X-ray portable
C1644647|Views portable:Find:Pt:Femur.left:Doc:XR
C1644647|Views portable:Finding:Point in time:Femur.left:Document:XR
C1645317|Knee - left X-ray 2 views and tunnel
C1645317|Knee-L XR 2V+Tunnel
C1645317|Views 2 & tunnel:Find:Pt:Knee.left:Doc:XR
C1645317|Views 2 & tunnel:Finding:Point in time:Knee.left:Document:XR
C1633482|Head CT W 133Xe IH
C1633482|Multisection^W Xe-133 Inhalation:Finding:Point in time:Head:Document:Computerized Tomography
C1633482|Head CT W Xe-133 IH
C1633482|Multisection^W Xe-133 IH:Find:Pt:Head:Doc:CT
C1714526|Foot - right X-ray 3 or 4 views
C1714526|Ft-R XR 3V or 4V
C1714526|Views 3 or 4:Finding:Point in time:Foot.right:Document:XR
C1714526|Views 3 or 4:Find:Pt:Foot.right:Doc:XR
C1714912|Axilla-R MRI WO+W contr IV
C1714912|Multisection^WO & W contrast IV:Find:Pt:Axilla.right:Doc:MRI
C1714912|Multisection^WO & W contrast Intravenous:Finding:Point in time:Axilla.right:Document:MRI
C1714912|Axilla - right MRI WO and W contrast IV
C1714923|Skull X-ray GE 5 views
C1714923|Skull XR GE 5V
C1714923|Views GE 5:Find:Pt:Skull:Doc:XR
C1714923|Views GE 5:Finding:Point in time:Skull:Document:XR
C1714785|Mammogram Guidance for needle biopsy of Breast - right
C1714785|Brst-R Mam Bx needle guid
C1714785|Guidance for biopsy.needle:Finding:Point in time:Breast.right:Document:Mam
C1714785|Guidance for biopsy.needle:Find:Pt:Breast.right:Doc:Mam
C1714945|Lower leg ves-R MRI.Angio
C1714945|Lower leg vessels - right MRI angiogram
C1714945|Multisection:Finding:Point in time:Lower leg vessels.right:Document:MRI.angio
C1714945|Multisection:Find:Pt:Lower leg vessels.right:Doc:MRI.angio
C1714947|XXX Flr DC change guide W contr IV
C1714947|Fluoroscopy Guidance for change of dialysis catheter in Unspecified body region-- W contrast IV
C1714947|Guidance for change of dialysis catheter^W contrast IV:Find:Pt:XXX:Doc:XR.fluor
C1714947|Guidance for change of dialysis catheter^W contrast Intravenous:Finding:Point in time:To be specified in another part of the message:Document:XR.fluor
C1717261|Skeletal Sys Axial RI BDM
C1717261|Skeletal system.axial Scan Bone density
C1717261|Bone density:Finding:Point in time:Skeletal system.axial:Document:Radnuc
C1717261|Bone density:Find:Pt:Skeletal system.axial:Doc:Radnuc
C1715016|Brain RI Flow W Tc99mGHA IV
C1715016|Brain Scan flow W Tc-99m glucoheptonate IV
C1715016|Views flow^W Tc-99m glucoheptonate IV:Find:Pt:Brain:Doc:Radnuc
C1715016|Views flow^W Tc-99m glucoheptonate Intravenous:Finding:Point in time:Brain:Document:Radnuc
C1715089|Vein-Bl XRA Thrombect guid W contr IV
C1715089|Fluoroscopic angiogram Guidance for thrombectomy of Vein - bilateral-- W contrast IV
C1715089|Guidance for thrombectomy^W contrast Intravenous:Finding:Point in time:Vein.bilateral:Document:XR.fluor.angio
C1715089|Guidance for thrombectomy^W contrast IV:Find:Pt:Vein.bilateral:Doc:XR.fluor.angio
C1715100|Kidney MRI WO contrast
C1715100|Kidney MRI WO contr
C1715100|Multisection^WO contrast:Finding:Point in time:Kidney:Document:MRI
C1715100|Multisection^WO contrast:Find:Pt:Kidney:Doc:MRI
C1715115|Liver+BDs+GB RI for Pat W Tc99mIV
C1715115|Liver and Biliary ducts and Gallbladder Scan for patency W Tc-99m IV
C1715115|Views for patency^W Tc-99m Intravenous:Finding:Point in time:Liver+Biliary ducts+Gallbladder:Document:Radnuc
C1715115|Views for patency^W Tc-99m IV:Find:Pt:Liver+Biliary ducts+Gallbladder:Doc:Radnuc
C1715118|Tibioperonl aa-R XRA Angpsty W contr IA
C1715118|Tibioperoneal arteries - right Fluoroscopic angiogram Angioplasty W contrast IA
C1715118|Angioplasty^W contrast Intra-arterial:Finding:Point in time:Tibioperoneal arteries.right:Document:XR.fluor.angio
C1715118|Angioplasty^W contrast IA:Find:Pt:Tibioperoneal arteries.right:Doc:XR.fluor.angio
C1645332|ST XR Lat+Towne
C1645332|Sella turcica X-ray lateral and Towne
C1645332|Views lateral & Towne:Find:Pt:Sella turcica:Doc:XR
C1645332|Views lateral & Towne:Finding:Point in time:Sella turcica:Document:XR
C1624108|Chest+Abd XR AP+Pa Chst
C1624108|Chest and Abdomen X-ray AP and PA chest
C1624108|Views AP & PA chest:Find:Pt:Chest+Abdomen:Doc:XR
C1624108|Views AP & PA chest:Finding:Point in time:Chest+Abdomen:Document:XR
C1631258|Chest+Abd CT WO+W contr IV
C1631258|Multisection^WO & W contrast IV:Find:Pt:Chest+Abdomen:Doc:CT
C1631258|Chest and Abdomen CT WO and W contrast IV
C1631258|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest+Abdomen:Document:Computerized Tomography
C1631786|Guidance for drainage of abscess:Finding:Point in time:Abdomen>Liver:Document:Computerized Tomography
C1631786|Guidance for drainage of abscess:Find:Pt:Abdomen>Liver:Doc:CT
C1631786|CT Guidance for drainage of abscess of Liver
C1631786|Liver CT Abscess drain guid
C1639940|Spine X-ray oblique single view
C1639940|Spine XR Obl 1V
C1639940|View oblique:Find:Pt:Spine:Doc:XR
C1639940|View oblique:Finding:Point in time:Spine:Document:XR
C1624699|XXX Flr <1h
C1624699|Unspecified body region Fluoroscopy Less than 1 hour
C1624699|View:Find:Lt 1H:XXX:Doc:XR.fluor
C1624699|View:Finding:Less than 1 hour:To be specified in another part of the message:Document:XR.fluor
C1625219|RI W In-111-T IV
C1625219|Scan W In-111 tiuxetan IV
C1625219|Views^W In-111 tiuxetan Intravenous:Finding:Point in time:^Patient:Document:Radnuc
C1625219|Views^W In-111 tiuxetan IV:Find:Pt:^Patient:Doc:Radnuc
C1954302|Upper extremity vein - right US
C1954302|UE v-R US
C1954302|Multisection:Find:Pt:Upper extremity vein.right:Doc:US
C1954302|Multisection:Finding:Point in time:Upper extremity vein.right:Document:Ultrasound
C1953986|Foot - bilateral X-ray GE 3 views
C1953986|Ft-Bl XR GE 3V
C1953986|Views GE 3:Finding:Point in time:Foot.bilateral:Document:XR
C1953986|Views GE 3:Find:Pt:Foot.bilateral:Doc:XR
C2734943|Lung PET
C2734943|Multisection:Find:Pt:Lung:Doc:Radnuc.PET
C2734943|Multisection:Finding:Point in time:Lung:Document:Radnuc.PET
C3169582|Guidance for percutaneous drainage:Find:Pt:XXX:Doc:US
C3169582|XXX US PC drain guid
C3169582|US Guidance for percutaneous drainage of Unspecified body region
C3169582|Guidance for percutaneous drainage:Finding:Point in time:To be specified in another part of the message:Document:Ultrasound
C3533567|Extr v-L US Laser ablation guid
C3533567|Guidance for laser ablation of vein(s):Find:Pt:Extremity vein.left:Doc:US
C3533567|US Guidance for laser ablation of vein(s) of Extremity vein - left
C3533567|Guidance for laser ablation of vein(s):Finding:Point in time:Extremity vein.left:Document:Ultrasound
C3533557|Guidance for replacement of percutaneous drainage tube:Finding:Point in time:Biliary ducts+Gallbladder:Document:XR.fluor
C3533557|Guidance for replacement of percutaneous drainage tube:Find:Pt:Biliary ducts+Gallbladder:Doc:XR.fluor
C3533557|BDs+GB Flr Replac of PC drain tube guid
C3533557|Fluoroscopy Guidance for replacement of percutaneous drainage tube in Biliary ducts and Gallbladder
C3262964|Knee-L XR 4V+AP stand
C3262964|Knee - left X-ray 4 views and AP standing
C3262964|Views 4 & AP^standing:Finding:Point in time:Knee.left:Document:XR
C3262964|Views 4 & AP^standing:Find:Pt:Knee.left:Doc:XR
C3262982|PA-Bl MRI.Angio W contr IA
C3262982|Pulmonary artery - bilateral MRI angiogram W contrast IA
C3262982|Multisection^W contrast Intra-arterial:Finding:Point in time:Pulmonary artery.bilateral:Document:MRI.angio
C3262982|Multisection^W contrast IA:Find:Pt:Pulmonary artery.bilateral:Doc:MRI.angio
C3263007|Upper extremity - bilateral MRI W contrast IV
C3263007|UE-Bl MRI W contr IV
C3263007|Multisection^W contrast Intravenous:Finding:Point in time:Upper extremity.bilateral:Document:MRI
C3263007|Multisection^W contrast IV:Find:Pt:Upper extremity.bilateral:Doc:MRI
C3263012|MRI Guidance for aspiration of cyst of Breast
C3263012|Brst MRI Cyst Asp guid
C3263012|Guidance for aspiration of cyst:Finding:Point in time:Breast:Document:MRI
C3263012|Guidance for aspiration of cyst:Find:Pt:Breast:Doc:MRI
C3263014|Finger MRI WO and W contrast IV
C3263014|Multisection^WO & W contrast Intravenous:Finding:Point in time:Finger:Document:MRI
C3263014|Multisection^WO & W contrast IV:Find:Pt:Finger:Doc:MRI
C3263014|Finger MRI WO+W contr IV
C3263053|Abd Flr PC Bx guid
C3263053|Fluoroscopy Guidance for percutaneous biopsy of Abdomen
C3263053|Guidance for percutaneous biopsy:Find:Pt:Abdomen:Doc:XR.fluor
C3263053|Guidance for percutaneous biopsy:Finding:Point in time:Abdomen:Document:XR.fluor
C3261469|Hand-L XR 1V
C3261469|Hand - left X-ray Single view
C3261469|View 1:Find:Pt:Hand.left:Doc:XR
C3261469|View 1:Finding:Point in time:Hand.left:Document:XR
C3261475|Radius+Ulna-R XR 1V
C3261475|Radius - right and Ulna - right X-ray Single view
C3261475|View 1:Finding:Point in time:Radius.right+Ulna.right:Document:XR
C3261475|View 1:Find:Pt:Radius.right+Ulna.right:Doc:XR
C3262894|Ribs - bilateral and Chest X-ray
C3262894|Views:Find:Pt:Ribs.bilateral+Chest:Doc:XR
C3262894|Views:Finding:Point in time:Ribs.bilateral+Chest:Document:XR
C3262894|Ribs-Bl+Chest XR
C3262902|Clavicle X-ray 45 degree cephalic angle
C3262902|Clavicle XR 45 Deg Ceph Angle
C3262902|View 45 degree cephalic angle:Find:Pt:Clavicle:Doc:XR
C3262902|View 45 degree cephalic angle:Finding:Point in time:Clavicle:Document:XR
C3262908|Multisection^WO & W contrast:Find:Pt:Abdomen>Renal vessels:Doc:CT.angio
C3262908|Deprecated Abdomen>Renal vessels CT angiogram WO and W contrast
C3262908|Deprecated Abd>Renal vls CT.Angio WO+W c
C3262908|Multisection^WO & W contrast:Finding:Point in time:Abdomen>Renal vessels:Document:Computerized Tomography.angio
C0203634|Nuclear medicine procedure
C0203634|Nuclear medicine
C0203634|Nuclear medicine procedure (procedure)
C0203634|Nuclear Medicine Procedures
C0203634|NM - Nuclear medicine
C0203634|Nuclear medicine procedure, NOS
C0203634|Radionuclide procedure, NOS
C0041618|Ultrasonography
C0041618|Imaging, Ultrasonic
C0041618|Diagnostic ultrasound
C0041618|ECHOTOMOGR
C0041618|ULTRASONOGR
C0041618|ECHOGR
C0041618|Medical Sonography
C0041618|Ultrasound imaging - action
C0041618|Ultrasound imaging
C0041618|sound measurement
C0041618|sonogram
C0041618|sonography
C0041618|Echography, NOS
C0041618|Echography
C0041618|GEN.US
C0041618|US
C0041618|Ultrasound procedure
C0041618|Ultrasound
C0041618|Imaging, Ultrasound
C0041618|Imagings, Ultrasound
C0041618|Ultrasound Imagings
C0041618|US - Ultrasound
C0041618|Ultrasonography (procedure)
C0041618|Ultrasound procedure (procedure)
C0041618|Ultrasound diagnostic procedure (procedure)
C0041618|Ultrasound scan (procedure)
C0041618|Ultrasound diagnostic procedure
C0041618|Ultrasound scan
C0041618|Ultrasonogram
C0041618|USS - Ultrasound scan
C0041618|ultrasound studies (procedure)
C0041618|ultrasound studies
C0041618|General ultrasound
C0041618|Diagnostic Ultrasound Procedures
C0041618|Ultrasonic imaging
C0041618|Unlisted ultrasound procedure (eg, diagnostic, interventional)
C0041618|UNLISTED US PROCEDURE
C0041618|Diagnostic ultrasound procedure
C0041618|Ultrasound, Diagnostic
C0041618|Diagnostic Ultrasounds
C0041618|Ultrasounds, Diagnostic
C0041618|Ultrasound scan NOS
C0041618|Sonography, Medical
C0041618|Echotomography
C0041618|Diagnostic ultrasonography
C0041618|Diagnostic sonar
C0041618|Ultrasound technique
C0041618|Diagnostic ultrasonography (procedure)
C0041618|Echography (procedure)
C0041618|Ultrasound imaging - action (qualifier value)
C0041618|Ultrasonography, NOS
C0041618|Diagnostic ultrasonography, NOS
C0041618|Ultrasound procedure, NOS
C0041618|Ultrasound scan, NOS
C0041618|ECHO EXAMINATION PROCEDURE
C0041618|Diagnosis (US)
C0041618|Diagnosis, Ultrasound
C0041618|Ultrasound Test
C0041618|Ultrasound, Medical
C0041618|ultrasound scanning
C0041618|ultrasound imaging/scanning
C0043299|Diagnostic radiologic examination
C0043299|RADIOL DIAG X RAY
C0043299|X Ray Radiology, Diagnostic
C0043299|DIAG X RAY
C0043299|Diagnostic X-Rays
C0043299|X-Rays, Diagnostic
C0043299|DIAG X RAY RADIOL
C0043299|ROENTGENOGR
C0043299|X RAY RADIOL DIAG
C0043299|X RAY DIAG
C0043299|X Ray, Diagnostic
C0043299|Diagnostic X Ray
C0043299|Radiology, Diagnostic X Ray
C0043299|Diagnostic X Ray Radiology
C0043299|Diagnostic radiography
C0043299|Diagnostic Radiology
C0043299|Radiology;diagnostic
C0043299|X-ray procedure
C0043299|X-Rays
C0043299|Diagnostic radiography (procedure)
C0043299|Diagnostic imaging procedure using X-rays (procedure)
C0043299|Diagnostic imaging procedure using X-rays
C0043299|Diagnostic radiology NOS
C0043299|Diagnostic radiology NOS (procedure)
C0043299|Diagnostic radiologic examination (procedure)
C0043299|Diagnostic Radiology (Diagnostic Imaging) Procedures
C0043299|Radiology, Diagnostic X-Ray
C0043299|Diagnostic X-Ray
C0043299|X-Ray, Diagnostic
C0043299|X-Ray Radiology, Diagnostic
C0043299|Diagnostic X-Ray Radiology
C0043299|Roentgenography
C0043299|Diagnostic radiologic examination, NOS
C0043299|Diagnostic radiography, NOS
C0043299|X-ray, NOS
C0043299|X Ray Diagnosis
C1742735|Breast, Mammography
C1740773|Bone/Joint Studies
C1689962|Radiologic Guidance
C1689962|Radiologic guidance procedure (procedure)
C1689962|Radiologic guidance procedure
C1522449|Radiotherapies
C1522449|Radiotherapy
C1522449|radiation therapy
C1522449|Radiation
C1522449|RT
C1522449|RADIOTHER
C1522449|radiation therapy (treatment)
C1522449|irradiation
C1522449|Therapeutic radiology
C1522449|Irradiate
C1522449|Irradiated
C1522449|Radiotherapy (regime/therapy)
C1522449|Radiation therapy (procedure)
C1522449|radiation therapy and/or radiation oncology
C1522449|radiation therapy and/or radiation oncology (treatment)
C1522449|Radiation therapy procedure or service
C1522449|radiation therapy procedure or service (treatment)
C1522449|Radiation Oncology Treatment
C1522449|Radiotherapy NOS
C1522449|RT - Radiotherapy
C1522449|Radiotherapy procedures
C1522449|Radiation oncology AND/OR radiotherapy (procedure)
C1522449|Radiation oncology AND/OR radiotherapy
C1522449|Radiation therapy procedure or service (procedure)
C1522449|therapy, radiation
C1522449|Radiation therapy procedure or service, NOS
C1522449|Radiation therapy, NOS
C1522449|Radiotherapy, NOS
C1522449|Cancer Radiotherapy
C1522449|Radiotherapeutics
C1522449|Therapeutic radiology procedure
C1522449|Therapeutic radiology for cancer treatment
C3870147|Pl space - L CT Abscess drain guid
C3870147|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space.left:Document:Computerized Tomography
C3870147|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space.left:Doc:CT
C3870147|CT Guidance for drainage of abscess of Pleural space - Left
C3870215|Guidance for placement of nephrostomy tube:Finding:Point in time:Kidney:Document:Ultrasound
C3870215|Guidance for placement of nephrostomy tube:Find:Pt:Kidney:Doc:US
C3870215|Kidney US NT plac guid
C3870215|US Guidance for placement of nephrostomy tube in Kidney
C3870149|Guidance for percutaneous biopsy:Find:Pt:Intervertebral disc:Doc:XR.fluor
C3870149|Guidance for percutaneous biopsy:Finding:Point in time:Intervertebral disc:Document:XR.fluor
C3870149|Fluoroscopy Guidance for percutaneous biopsy of Intervertebral disc
C3870149|I-disc Flr PC Bx guid
C3870151|Guidance for percutaneous aspiration:Finding:Point in time:Spine.cervical>Intervertebral disc:Document:Computerized Tomography
C3870151|C-spine interv disc CT PC Asp guid
C3870151|CT Guidance for percutaneous aspiration of Cervical spine Intervertebral disc
C3870151|Guidance for percutaneous aspiration:Find:Pt:Spine.cervical>Intervertebral disc:Doc:CT
C3870153|CT Guidance for drainage of abscess of Pleural space - Bilateral
C3870153|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space.bilateral:Doc:CT
C3870153|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space.bilateral:Document:Computerized Tomography
C3870153|Pl space-Bl CT Abscess drain guid
C3870218|Guidance for biopsy:Find:Pt:Bone marrow:Doc:XR.fluor
C3870218|Guidance for biopsy:Finding:Point in time:Bone marrow:Document:XR.fluor
C3870218|Fluoroscopy Guidance for biopsy of Bone marrow
C3870218|BM Flr Bx guid
C3870148|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space.left:Doc:XR.fluor
C3870148|Pl space - L Flr Abscess drain guid
C3870148|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space.left:Document:XR.fluor
C3870148|Fluoroscopy Guidance for drainage of abscess of Pleural space - Left
C3870216|Circle of Willis CT angiogram WO and W contrast IV
C3870216|Circle of Willis CT.Angio WO+W contr IV
C3870216|Multisection^WO & W contrast Intravenous:Finding:Point in time:Head+Neck>Circle of Willis:Document:Computerized Tomography.angio
C3870216|Multisection^WO & W contrast IV:Find:Pt:Head+Neck>Circle of Willis:Doc:CT.angio
C3870093|Views^W contrast EP:Find:Pt:Spine.thoracic.epidural space:Doc:XR.fluor.angio
C3870093|T-spine space XRA W contr EP
C3870093|Views^W contrast Epidural:Finding:Point in time:Spine.thoracic.epidural space:Document:XR.fluor.angio
C3870093|Spine thoracic epidural space Fluoroscopic angiogram W contrast EP
C3870152|Fluoroscopy Guidance for drainage of abscess of Pleural space - Bilateral
C3870152|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space.bilateral:Doc:XR.fluor
C3870152|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space.bilateral:Document:XR.fluor
C3870152|Pl space-Bl Flr Abscess drain guid
C3870055|Views^W contrast Vaginal:Finding:Point in time:Vaginal:Document:XR.fluor
C3870055|Vaginal Flr W contr VG
C3870055|Views^W contrast VG:Find:Pt:Vaginal:Doc:XR.fluor
C3870055|Vaginal Fluoroscopy W contrast VG
C3870217|Spine lumbar.epidural space Fluoroscopic angiogram W contrast EP
C3870217|Views^W contrast Epidural:Finding:Point in time:Spine.lumbar.epidural space:Document:XR.fluor.angio
C3870217|Views^W contrast EP:Find:Pt:Spine.lumbar.epidural space:Doc:XR.fluor.angio
C3870217|L-spine space XRA W contr EP
C3870150|Guidance for percutaneous aspiration:Finding:Point in time:Intervertebral disc:Document:XR.fluor
C3870150|Fluoroscopy Guidance for percutaneous aspiration of Intervertebral disc
C3870150|I-disc Flr PC Asp guid
C3870150|Guidance for percutaneous aspiration:Find:Pt:Intervertebral disc:Doc:XR.fluor
C3870091|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space.right:Document:XR.fluor
C3870091|Fluoroscopy Guidance for drainage of abscess of Pleural space - Right
C3870091|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space.right:Doc:XR.fluor
C3870091|Pl space - R Flr Abscess drain guid
C3870090|Guidance for drainage of abscess:Finding:Point in time:Chest>Pleural space.right:Document:Computerized Tomography
C3870090|CT Guidance for drainage of abscess of Pleural space - Right
C3870090|Guidance for drainage of abscess:Find:Pt:Chest>Pleural space.right:Doc:CT
C3870090|Pl space - R CT Abscess drain guid
C4036866|Hind+Mid ft-R XR 2V
C4036866|Views 2:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4036866|Views 2:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036866|Hindfoot - right and Midfoot - right X-ray 2 views
C4036855|Hind+Mid ft-R XR stand
C4036855|Views^standing:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036855|Views^standing:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4036855|Hindfoot - right and Midfoot - right X-ray standing
C4037011|Multisection for endograft:Finding:Point in time:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+Vessels.bilateral:Document:Computerized Tomography.angio
C4037011|Abdominal Aorta and Bilateral Vessels CT angiogram for endograft
C4037011|Abd Aorta+Ves-Bl CT.Angio for endograft
C4037011|Multisection for endograft:Find:Pt:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+Vessels.bilateral:Doc:CT.angio
C4037010|Multisection^W contrast IV:Find:Pt:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+Vessels.bilateral:Doc:CT.angio
C4037010|Deprecated Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+Vessels CT angiogram W contrast IV
C4037010|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+Vessels.bilateral:Document:Computerized Tomography.angio
C4037010|Deprecated Ab+Pl+Lx.b>A.ab+V CT.Angio W
C4036884|Hind+Mid ft DXA BDM
C4036884|Bone density:MAric:Pt:Hindfoot+Midfoot:Qn:XR.DXA
C4036884|Bone density:Mass Aeric:Point in time:Hindfoot+Midfoot:Quantitative:XR.DXA
C4036884|Hindfoot and Midfoot DXA Bone density
C4036880|Multisection^WO & W contrast IV:Find:Pt:Hindfoot+Midfoot:Doc:CT
C4036880|Hind+Mid ft CT WO+W contr IV
C4036880|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hindfoot+Midfoot:Document:Computerized Tomography
C4036880|Hindfoot and Midfoot CT WO and W contrast IV
C4036878|View 1:Find:Pt:Hindfoot+Midfoot:Doc:XR
C4036878|View 1:Finding:Point in time:Hindfoot+Midfoot:Document:XR
C4036878|Hind+Mid ft XR 1V
C4036878|Hindfoot and Midfoot X-ray Single view
C4037651|Hind+Mid ft-R CT WO+W contr IV
C4037651|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:Computerized Tomography
C4037651|Multisection^WO & W contrast IV:Find:Pt:Hindfoot.right+Midfoot.right:Doc:CT
C4037651|Hindfoot - right and Midfoot - right CT WO and W contrast IV
C4036859|Hind+Mid ft-Bl XR Ski Jump
C4036859|Views ski jump:Find:Pt:Hindfoot.bilateral+Midfoot.bilateral:Doc:XR
C4036859|Views ski jump:Finding:Point in time:Hindfoot.bilateral+Midfoot.bilateral:Document:XR
C4036859|Hindfoot - bilateral and Midfoot - bilateral X-ray ski jump
C4036856|Hind+Mid ft-L XR stand
C4036856|Views^standing:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4036856|Views^standing:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4036856|Hindfoot - left and Midfoot - left X-ray standing
C4036877|Hind+Mid ft XR
C4036877|Views:Find:Pt:Hindfoot+Midfoot:Doc:XR
C4036877|Views:Finding:Point in time:Hindfoot+Midfoot:Document:XR
C4036877|Hindfoot and Midfoot X-ray
C4037658|Views AP & lateral & oblique:Find:Pt:Hindfoot+Midfoot:Doc:XR
C4037658|Views AP & lateral & oblique:Finding:Point in time:Hindfoot+Midfoot:Document:XR
C4037658|Hind+Mid ft XR AP+Lat+Obl
C4037658|Hindfoot and Midfoot X-ray AP and lateral and oblique
C4037652|Hind+Mid ft-L CT WO+W contr IV
C4037652|Multisection^WO & W contrast Intravenous:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:Computerized Tomography
C4037652|Hindfoot - left and Midfoot - left CT WO and W contrast IV
C4037652|Multisection^WO & W contrast IV:Find:Pt:Hindfoot.left+Midfoot.left:Doc:CT
C4036871|Views:Find:Pt:Hindfoot.bilateral+Midfoot.bilateral:Doc:XR
C4036871|Hind+Mid ft-Bl XR
C4036871|Hindfoot - bilateral and Midfoot - bilateral X-ray
C4036871|Views:Finding:Point in time:Hindfoot.bilateral+Midfoot.bilateral:Document:XR
C4036867|Hind+Mid ft-L XR 2V
C4036867|Hindfoot - left and Midfoot - left X-ray 2 views
C4036867|Views 2:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4036867|Views 2:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4036865|Views AP & lateral:Find:Pt:Hindfoot.bilateral+Midfoot.bilateral:Doc:XR
C4036865|Views AP & lateral:Finding:Point in time:Hindfoot.bilateral+Midfoot.bilateral:Document:XR
C4036865|Hind+Mid ft-Bl XR AP+Lat
C4036865|Hindfoot - bilateral and Midfoot - bilateral X-ray AP and lateral
C4036766|Liver stiffness by US.transient elastography
C4036766|Liver stiffness:Pressure:Point in time:Liver:Quantitative:Ultrasound.transient elastography
C4036766|Liver stiffness US.TE
C4036766|Liver stiffness:Pres:Pt:Liver:Qn:US.transient elastography
C4036483|Multisection^WO & W contrast Intravenous:Finding:Point in time:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+RO vessels.bilateral:Document:Computerized Tomography.angio
C4036483|T+A.Ao+RO v-Bl CT.Angio WO+W contr IV
C4036483|Multisection^WO & W contrast IV:Find:Pt:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+RO vessels.bilateral:Doc:CT.angio
C4036483|Thoracic and Abdominal Aorta and Bilateral Runoff Vessels CT angiogram WO and W contrast IV
C4036886|Multisection for endograft:Find:Pt:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+Vessels.bilateral:Doc:CT.angio
C4036886|Thoracic and Abdominal Aorta and Bilateral Vessels CT angiogram for endograft
C4036886|T Ao+Abd Ao+Ves-Bl CT.Angio for endograf
C4036886|Multisection for endograft:Finding:Point in time:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+Vessels.bilateral:Document:Computerized Tomography.angio
C4036879|Hind+Mid ft CT WO contr
C4036879|Multisection^WO contrast:Finding:Point in time:Hindfoot+Midfoot:Document:Computerized Tomography
C4036879|Multisection^WO contrast:Find:Pt:Hindfoot+Midfoot:Doc:CT
C4036879|Hindfoot and Midfoot CT WO contrast
C4037657|Hind+Mid ft XR Broden
C4037657|Views Broden:Finding:Point in time:Hindfoot+Midfoot:Document:XR
C4037657|Views Broden:Find:Pt:Hindfoot+Midfoot:Doc:XR
C4037657|Hindfoot and Midfoot X-ray Broden
C4037650|Hind+Mid ft-L CT WO contr
C4037650|Hindfoot - left and Midfoot - left CT WO contrast
C4037650|Multisection^WO contrast:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:Computerized Tomography
C4037650|Multisection^WO contrast:Find:Pt:Hindfoot.left+Midfoot.left:Doc:CT
C4036862|Views Broden:Find:Pt:Hindfoot.bilateral+Midfoot.bilateral:Doc:XR
C4036862|Hindfoot - bilateral and Midfoot - bilateral X-ray Broden
C4036862|Views Broden:Finding:Point in time:Hindfoot.bilateral+Midfoot.bilateral:Document:XR
C4036862|Hind+Mid ft-Bl XR Broden
C4036858|Hind+Mid ft-L XR Ski Jump
C4036858|Views ski jump:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4036858|Views ski jump:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4036858|Hindfoot - left and Midfoot - left X-ray ski jump
C4036484|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+RO vessels.bilateral:Document:Computerized Tomography.angio
C4036484|Multisection^WO & W contrast IV:Find:Pt:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+RO vessels.bilateral:Doc:CT.angio
C4036484|Abdominal Aorta and Bilateral Runoff Vessels CT angiogram WO and W contrast IV
C4036484|Abd Aorta+ROves-Bl CT.Angio WO+WcontrIV
C4036876|Views 2:Finding:Point in time:Hindfoot+Midfoot:Document:XR
C4036876|Hind+Mid ft XR 2V
C4036876|Views 2:Find:Pt:Hindfoot+Midfoot:Doc:XR
C4036876|Hindfoot and Midfoot X-ray 2 views
C4037656|Views ski jump:Find:Pt:Hindfoot+Midfoot:Doc:XR
C4037656|Hind+Mid ft XR Ski Jump
C4037656|Views ski jump:Finding:Point in time:Hindfoot+Midfoot:Document:XR
C4037656|Hindfoot and Midfoot X-ray ski jump
C4036868|Views 2:Finding:Point in time:Hindfoot.bilateral+Midfoot.bilateral:Document:XR
C4036868|Views 2:Find:Pt:Hindfoot.bilateral+Midfoot.bilateral:Doc:XR
C4036868|Hindfoot - bilateral and Midfoot - bilateral X-ray 2 views
C4036868|Hind+Mid ft-Bl XR 2V
C4036863|Hind+Mid ft-R XR AP+Lat
C4036863|Hindfoot - right and Midfoot - right X-ray AP and lateral
C4036863|Views AP & lateral:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036863|Views AP & lateral:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4036861|Hind+Mid ft-L XR Broden
C4036861|Hindfoot - left and Midfoot - left X-ray Broden
C4036861|Views Broden:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4036861|Views Broden:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4036480|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+RO vessels.bilateral:Document:Computerized Tomography.angio
C4036480|Multisection^W contrast IV:Find:Pt:Abdomen+Pelvis+Lower extremity.bilateral>Aorta.abdominal+RO vessels.bilateral:Doc:CT.angio
C4036480|Abdominal Aorta and Bilateral Runoff Vessels CT angiogram W contrast IV
C4036480|Abd Aorta+RO ves-Bl CT.Angio W contr IV
C4036888|Multisection:Finding:Point in time:Hindfoot+Midfoot:Document:Computerized Tomography
C4036888|Multisection:Find:Pt:Hindfoot+Midfoot:Doc:CT
C4036888|Hind+Mid ft CT
C4036888|Hindfoot and Midfoot CT
C4037654|Hind+Mid ft-L CT W contr IV
C4037654|Multisection^W contrast Intravenous:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:Computerized Tomography
C4037654|Hindfoot - left and Midfoot - left CT W contrast IV
C4037654|Multisection^W contrast IV:Find:Pt:Hindfoot.left+Midfoot.left:Doc:CT
C4037653|Hind+Mid ft-R CT W contr IV
C4037653|Hindfoot - right and Midfoot - right CT W contrast IV
C4037653|Multisection^W contrast IV:Find:Pt:Hindfoot.right+Midfoot.right:Doc:CT
C4037653|Multisection^W contrast Intravenous:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:Computerized Tomography
C4037647|Hind+Mid ft-R XR 1V
C4037647|Hindfoot - right and Midfoot - right X-ray Single view
C4037647|View 1:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4037647|View 1:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036875|Hindfoot - bilateral and Midfoot - bilateral X-ray Harris
C4036875|View Harris:Finding:Point in time:Hindfoot.bilateral+Midfoot.bilateral:Document:XR
C4036875|View Harris:Find:Pt:Hindfoot.bilateral+Midfoot.bilateral:Doc:XR
C4036875|Hind+Mid ft-Bl XR Harris
C4036874|Hind+Mid ft-L XR Harris
C4036874|View Harris:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4036874|Hindfoot - left and Midfoot - left X-ray Harris
C4036874|View Harris:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4036873|Hind+Mid ft-R XR Harris
C4036873|View Harris:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036873|Hindfoot - right and Midfoot - right X-ray Harris
C4036873|View Harris:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4036872|Hind+Mid ft-Bl XR stand
C4036872|View^standing:Finding:Point in time:Hindfoot.bilateral+Midfoot.bilateral:Document:XR
C4036872|Hindfoot - bilateral and Midfoot - bilateral X-ray standing
C4036872|View^standing:Find:Pt:Hindfoot.bilateral+Midfoot.bilateral:Doc:XR
C4036864|Hind+Mid ft-L XR AP+Lat
C4036864|Views AP & lateral:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4036864|Views AP & lateral:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4036864|Hindfoot - left and Midfoot - left X-ray AP and lateral
C4036857|Hind+Mid ft-R XR Ski Jump
C4036857|Views ski jump:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036857|Views ski jump:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4036857|Hindfoot - right and Midfoot - right X-ray ski jump
C4036887|Multisection^W contrast IV:Find:Pt:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+Vessels.bilateral:Doc:CT.angio
C4036887|Deprecated Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+vessels CT angiogram W contrast IV
C4036887|Multisection^W contrast Intravenous:Finding:Point in time:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+Vessels.bilateral:Document:Computerized Tomography.angio
C4036887|Deprecated C+A+P+LxB>A.th+A CT.Angio W c
C4037655|Hind+Mid ft XR stand
C4037655|Views^standing:Find:Pt:Hindfoot+Midfoot:Doc:XR
C4037655|Views^standing:Finding:Point in time:Hindfoot+Midfoot:Document:XR
C4037655|Hindfoot and Midfoot X-ray standing
C4036870|Hind+Mid ft-L XR
C4036870|Hindfoot - left and Midfoot - left X-ray
C4036870|Views:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4036870|Views:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4036869|Hind+Mid ft-R XR
C4036869|Hindfoot - right and Midfoot - right X-ray
C4036869|Views:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036869|Views:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4036860|Hind+Mid ft-R XR Broden
C4036860|Views Broden:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:XR
C4036860|Hindfoot - right and Midfoot - right X-ray Broden
C4036860|Views Broden:Find:Pt:Hindfoot.right+Midfoot.right:Doc:XR
C4036883|Bone density:Tscore:Pt:Hindfoot+Midfoot:Qn:XR.DXA
C4036883|Bone density:T Score:Point in time:Hindfoot+Midfoot:Quantitative:XR.DXA
C4036883|Hind+Mid ft DXA T-score BDM
C4036883|Hindfoot and Midfoot DXA [T-score] Bone density
C4036882|Multisection:Find:Pt:Hindfoot+Midfoot:Doc:XR.tomo
C4036882|Hind+Mid ft XRTomo
C4036882|Multisection:Finding:Point in time:Hindfoot+Midfoot:Document:XR.tomo
C4036882|Hindfoot and Midfoot X-ray tomograph
C4036881|Multisection^W contrast Intravenous:Finding:Point in time:Hindfoot+Midfoot:Document:Computerized Tomography
C4036881|Hind+Mid ft CT W contr IV
C4036881|Multisection^W contrast IV:Find:Pt:Hindfoot+Midfoot:Doc:CT
C4036881|Hindfoot and Midfoot CT W contrast IV
C4037649|Hind+Mid ft-R CT WO contr
C4037649|Hindfoot - right and Midfoot - right CT WO contrast
C4037649|Multisection^WO contrast:Find:Pt:Hindfoot.right+Midfoot.right:Doc:CT
C4037649|Multisection^WO contrast:Finding:Point in time:Hindfoot.right+Midfoot.right:Document:Computerized Tomography
C4037648|Hind+Mid ft-L XR 1V
C4037648|View 1:Finding:Point in time:Hindfoot.left+Midfoot.left:Document:XR
C4037648|View 1:Find:Pt:Hindfoot.left+Midfoot.left:Doc:XR
C4037648|Hindfoot - left and Midfoot - left X-ray Single view
C4036479|Multisection^W contrast Intravenous:Finding:Point in time:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+RO vessels.bilateral:Document:Computerized Tomography.angio
C4036479|Thoracic and Abdominal Aorta and Bilateral Runoff Vessels CT angiogram W contrast IV
C4036479|T+A.Ao+RO v-Bl CT.Angio W contr IV
C4036479|Multisection^W contrast IV:Find:Pt:Chest+Abdomen+Pelvis+Lower extremity.bilateral>Aorta.thoracic+Aorta.abdominal+RO vessels.bilateral:Doc:CT.angio
C4070485|Colon and Rectum CT W contrast IV
C4070485|Colon+Rectum CT W contr IV
C4070485|Multisection^W contrast IV:Find:Pt:Abdomen+Pelvis>Colon+Rectum:Doc:CT
C4070485|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis>Colon+Rectum:Document:Computerized Tomography
C4070471|Multisection by reconstruction^WO contrast:Find:Pt:Head>Temporal bone:Doc:CT
C4070471|Multisection by reconstruction^WO contrast:Finding:Point in time:Head>Temporal bone:Document:Computerized Tomography
C4070471|Temporal bone CT by reconstruction WO contrast
C4070471|Temporal bone CT by reconstr WO contr
C4070709|Views GE 2:Finding:Point in time:Hip.right:Document:XR
C4070709|Hip - right X-ray GE 2 views
C4070709|Views GE 2:Find:Pt:Hip.right:Doc:XR
C4070709|Hip-R XR GE 2V
C4070707|Views GE 2:Find:Pt:Humerus:Doc:XR
C4070707|Humerus XR GE 2V
C4070707|Humerus X-ray GE 2 views
C4070707|Views GE 2:Finding:Point in time:Humerus:Document:XR
C4070461|Blad CT W contr IUB
C4070461|Multisection^W contrast intra bladder:Find:Pt:Pelvis>Urinary bladder:Doc:CT
C4070461|Multisection^W contrast intra bladder:Finding:Point in time:Pelvis>Urinary bladder:Document:Computerized Tomography
C4070461|Urinary bladder CT W contrast intra bladder
C4070456|Pelvis CT 3D post processing WO contrast
C4070456|Pelvis CT p 3D proc WO contr
C4070456|Multisection 3D post processing^WO contrast:Finding:Point in time:Pelvis:Document:Computerized Tomography
C4070456|Multisection 3D post processing^WO contrast:Find:Pt:Pelvis:Doc:CT
C4070260|Views GE 2:Finding:Point in time:Spine.cervical:Document:XR
C4070260|C-spine XR GE 2V
C4070260|Cervical spine X-ray GE 2 views
C4070260|Views GE 2:Find:Pt:Spine.cervical:Doc:XR
C4070259|Views GE 6:Find:Pt:Spine.cervical:Doc:XR
C4070259|Cervical spine X-ray GE 6 views
C4070259|C-spine XR GE 6V
C4070259|Views GE 6:Finding:Point in time:Spine.cervical:Document:XR
C4070483|Guidance for radiation treatment:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C4070483|XXX CT RT guid
C4070483|Guidance for radiation treatment:Find:Pt:XXX:Doc:CT
C4070483|CT Guidance for radiation treatment of Unspecified body region
C4070474|Multisection by reconstruction^WO contrast:Find:Pt:Spine.lumbar:Doc:CT
C4070474|Multisection by reconstruction^WO contrast:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C4070474|Lumbar spine CT by reconstruction WO contrast
C4070474|L-spine CT by reconstr WO contr
C4070473|Multisection by reconstruction^W contrast Intravenous:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C4070473|Thoracic spine CT by reconstruction W contrast IV
C4070473|Multisection by reconstruction^W contrast IV:Find:Pt:Spine.thoracic:Doc:CT
C4070473|T-spine CT by reconstr W contr IV
C4070468|Heart CT for calcium scoring WO contrast
C4070468|Multisection for calcium score^WO contrast:Find:Pt:Chest>Heart:Doc:CT
C4070468|Hrt CT for Calcium Score WO contr
C4070468|Multisection for calcium score^WO contrast:Finding:Point in time:Chest>Heart:Document:Computerized Tomography
C4071446|Hand XR 1V or 2V
C4071446|Views 1 or 2:Finding:Point in time:Hand:Document:XR
C4071446|Views 1 or 2:Find:Pt:Hand:Doc:XR
C4071446|Hand X-ray 1 or 2 views
C4070705|Views GE 4:Finding:Point in time:Knee:Document:XR
C4070705|Views GE 4:Find:Pt:Knee:Doc:XR
C4070705|Knee X-ray GE 4 views
C4070705|Knee XR GE 4V
C4070258|Ribs - bilateral X-ray GE 3 views
C4070258|Views GE 3:Finding:Point in time:Ribs.bilateral:Document:XR
C4070258|Views GE 3:Find:Pt:Ribs.bilateral:Doc:XR
C4070258|Ribs-Bl XR GE 3V
C4070252|Views GE 2:Finding:Point in time:Spine.lumbar+Sacrum:Document:XR
C4070252|L-spine+Sacrum XR GE 2V
C4070252|Spine Lumbar and Sacrum X-ray GE 2 views
C4070252|Views GE 2:Find:Pt:Spine.lumbar+Sacrum:Doc:XR
C4070465|L-spine CT.Dens WO contr
C4070465|Multisection^WO contrast:Find:Pt:Spine.lumbar:Doc:CT.densitometry
C4070465|Multisection^WO contrast:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography.densitometry
C4070465|Lumbar spine CT densitometry WO contrast
C4070460|Multisection:Finding:Point in time:Maxilla+Mandible>Teeth:Document:Computerized Tomography
C4070460|Teeth CT
C4070460|Multisection:Find:Pt:Maxilla+Mandible>Teeth:Doc:CT
C4070455|Multisection for screening:Find:Pt:Abdomen+Pelvis>Colon+Rectum:Doc:CT
C4070455|Colon+Rectum CT Screening
C4070455|Colon and Rectum CT for screening
C4070455|Multisection for screening:Finding:Point in time:Abdomen+Pelvis>Colon+Rectum:Document:Computerized Tomography
C4071408|Views GE 6:Finding:Point in time:Spine.lumbar+Sacrum:Document:XR
C4071408|Views GE 6:Find:Pt:Spine.lumbar+Sacrum:Doc:XR
C4071408|Spine Lumbar and Sacrum X-ray GE 6 views
C4071408|L-spine+Sacrum XR GE 6V
C4070486|Colon+Rectum CT Screening WO contr
C4070486|Multisection for screening^WO contrast:Find:Pt:Abdomen+Pelvis>Colon+Rectum:Doc:CT
C4070486|Colon and Rectum CT for screening WO contrast
C4070486|Multisection for screening^WO contrast:Finding:Point in time:Abdomen+Pelvis>Colon+Rectum:Document:Computerized Tomography
C4070479|Pelvis CT by reconstruction WO contrast
C4070479|Pelvis CT by reconstr WO contr
C4070479|Multisection by reconstruction^WO contrast:Finding:Point in time:Pelvis:Document:Computerized Tomography
C4070479|Multisection by reconstruction^WO contrast:Find:Pt:Pelvis:Doc:CT
C4070476|Multisection by reconstruction^WO contrast:Find:Pt:Spine.cervical:Doc:CT
C4070476|Cervical spine CT by reconstruction WO contrast
C4070476|Multisection by reconstruction^WO contrast:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C4070476|C-spine CT by reconstr WO contr
C4070470|Multisection^WO & W contrast IV:Find:Pt:Abdomen>Biliary ducts:Doc:CT
C4070470|Multisection^WO & W contrast Intravenous:Finding:Point in time:Abdomen>Biliary ducts:Document:Computerized Tomography
C4070470|Biliary ducts CT WO and W contrast IV
C4070470|BD CT WO+W contr IV
C4071445|Views GE 3:Find:Pt:Hand:Doc:XR
C4071445|Hand X-ray GE 3 views
C4071445|Views GE 3:Finding:Point in time:Hand:Document:XR
C4071445|Hand XR GE 3V
C4070706|Knee-Bl XR AP+Lat+Merchants stand
C4070706|Knee - bilateral X-ray AP and lateral and Merchants standing
C4070706|Views AP & lateral & Merchants^standing:Finding:Point in time:Knee.bilateral:Document:XR
C4070706|Views AP & lateral & Merchants^standing:Find:Pt:Knee.bilateral:Doc:XR
C4070458|Chest and Abdomen CT 3D post processing WO contrast
C4070458|Chest+Abd CT p 3D proc WO contr
C4070458|Multisection 3D post processing^WO contrast:Find:Pt:Chest+Abdomen:Doc:CT
C4070458|Multisection 3D post processing^WO contrast:Finding:Point in time:Chest+Abdomen:Document:Computerized Tomography
C4071448|Views GE 2:Find:Pt:Finger:Doc:XR
C4071448|Finger X-ray GE 2 views
C4071448|Finger XR GE 2V
C4071448|Views GE 2:Finding:Point in time:Finger:Document:XR
C4070572|Multisection for leg measurement^WO contrast:Find:Pt:Lower extremity.bilateral:Doc:CT.scanogram
C4070572|Multisection for leg measurement^WO contrast:Finding:Point in time:Lower extremity.bilateral:Document:Computerized Tomography.scanogram
C4070572|Lower extremity - bilateral Computed tomography scanogram for leg measurement WO contrast
C4070572|LE-Bl CT.scanogram leg meas WO contr
C4070484|Multisection^WO contrast:Finding:Point in time:Abdomen+Pelvis>Colon+Rectum:Document:Computerized Tomography
C4070484|Colon and Rectum CT WO contrast
C4070484|Colon+Rectum CT WO contr
C4070484|Multisection^WO contrast:Find:Pt:Abdomen+Pelvis>Colon+Rectum:Doc:CT
C4070255|Views GE 2:Find:Pt:Shoulder.left:Doc:XR
C4070255|Views GE 2:Finding:Point in time:Shoulder.left:Document:XR
C4070255|Shoulder - left X-ray GE 2 views
C4070255|Should-L XR GE 2V
C4070250|Toe X-ray GE 2 views
C4070250|Views GE 2:Find:Pt:Toe:Doc:XR
C4070250|Toe XR GE 2V
C4070250|Views GE 2:Finding:Point in time:Toe:Document:XR
C4070466|Multisection^W contrast IV:Find:Pt:Chest>Heart:Doc:CT
C4070466|Multisection^W contrast Intravenous:Finding:Point in time:Chest>Heart:Document:Computerized Tomography
C4070466|Hrt CT W contr IV
C4070466|Heart CT W contrast IV
C4070453|Multisection^W contrast IV:Find:Pt:Abdomen:Doc:CT
C4070453|Multisection^W contrast Intravenous:Finding:Point in time:Abdomen:Document:Computerized Tomography
C4070453|Abd CT W contr IV
C4070453|Abdomen CT W contrast IV
C4070488|Multisection^WO contrast:Find:Pt:Chest>Airway:Doc:CT
C4070488|Airway CT WO contrast
C4070488|Multisection^WO contrast:Finding:Point in time:Chest>Airway:Document:Computerized Tomography
C4070488|Airway CT WO contr
C4070482|Heart and Coronary arteries CT angiogram W contrast IV
C4070482|Hrt+CA CT.Angio W contr IV
C4070482|Multisection^W contrast IV:Find:Pt:Chest>Heart+Coronary arteries:Doc:CT.angio
C4070482|Multisection^W contrast Intravenous:Finding:Point in time:Chest>Heart+Coronary arteries:Document:Computerized Tomography.angio
C4070477|Multisection by reconstruction^W contrast IV:Find:Pt:Spine.cervical:Doc:CT
C4070477|Cervical spine CT by reconstruction W contrast IV
C4070477|C-spine CT by reconstr W contr IV
C4070477|Multisection by reconstruction^W contrast Intravenous:Finding:Point in time:Spine.cervical:Document:Computerized Tomography
C4070475|Lumbar spine CT by reconstruction W contrast IV
C4070475|Multisection by reconstruction^W contrast IV:Find:Pt:Spine.lumbar:Doc:CT
C4070475|L-spine CT by reconstr W contr IV
C4070475|Multisection by reconstruction^W contrast Intravenous:Finding:Point in time:Spine.lumbar:Document:Computerized Tomography
C4070472|Multisection by reconstruction^W contrast IV:Find:Pt:Head>Temporal bone:Doc:CT
C4070472|Multisection by reconstruction^W contrast Intravenous:Finding:Point in time:Head>Temporal bone:Document:Computerized Tomography
C4070472|Temporal bone CT by reconstruction W contrast IV
C4070472|Temporal bone CT by reconstr W contr IV
C4071444|Hip-Bl XR GE 4V
C4071444|Hip - bilateral X-ray GE 4 views
C4071444|Views GE 4:Finding:Point in time:Hip.bilateral:Document:XR
C4071444|Views GE 4:Find:Pt:Hip.bilateral:Doc:XR
C4070710|Hip-L XR GE 2V
C4070710|Views GE 2:Find:Pt:Hip.left:Doc:XR
C4070710|Hip - left X-ray GE 2 views
C4070710|Views GE 2:Finding:Point in time:Hip.left:Document:XR
C4070708|Views GE 2:Finding:Point in time:Hip:Document:XR
C4070708|Hip XR GE 2V
C4070708|Views GE 2:Find:Pt:Hip:Doc:XR
C4070708|Hip X-ray GE 2 views
C4070253|Views GE 2:Finding:Point in time:Shoulder:Document:XR
C4070253|Views GE 2:Find:Pt:Shoulder:Doc:XR
C4070253|Should XR GE 2V
C4070253|Shoulder X-ray GE 2 views
C4070462|Multisection 3D post processing:Finding:Point in time:To be specified in another part of the message:Document:Computerized Tomography
C4070462|XXX CT p 3D proc
C4070462|Unspecified body region CT 3D post processing
C4070462|Multisection 3D post processing:Find:Pt:XXX:Doc:CT
C4070261|Abd XR GE 3V
C4070261|Views GE 3:Find:Pt:Abdomen:Doc:XR
C4070261|Abdomen X-ray GE 3 views
C4070261|Views GE 3:Finding:Point in time:Abdomen:Document:XR
C4070490|Abd+Pelvis CT p 3D proc WO contr
C4070490|Multisection 3D post processing^WO contrast:Finding:Point in time:Abdomen+Pelvis:Document:Computerized Tomography
C4070490|Abdomen and Pelvis CT 3D post processing WO contrast
C4070490|Multisection 3D post processing^WO contrast:Find:Pt:Abdomen+Pelvis:Doc:CT
C4070487|Multisection for screening^W contrast Intravenous:Finding:Point in time:Chest:Document:Computerized Tomography
C4070487|Chest CT Screening W contr IV
C4070487|Chest CT for screening W contrast IV
C4070487|Multisection for screening^W contrast IV:Find:Pt:Chest:Doc:CT
C4070469|Multisection for screening^WO contrast:Find:Pt:Chest:Doc:CT
C4070469|Multisection for screening^WO contrast:Finding:Point in time:Chest:Document:Computerized Tomography
C4070469|Chest CT for screening WO contrast
C4070469|Chest CT Screening WO contr
C4070467|Hrt CT for congenital disease W contr IV
C4070467|Multisection for congenital disease^W contrast Intravenous:Finding:Point in time:Chest>Heart:Document:Computerized Tomography
C4070467|Heart CT for congenital disease W contrast IV
C4070467|Multisection for congenital disease^W contrast IV:Find:Pt:Chest>Heart:Doc:CT
C4070257|Views 2:Finding:Point in time:Ribs.unilateral+Chest:Document:XR
C4070257|Ribs-Ul+chest XR 2V
C4070257|Ribs - unilateral and Chest X-ray 2 views
C4070257|Views 2:Find:Pt:Ribs.unilateral+Chest:Doc:XR
C4070254|Shoulder - right X-ray GE 2 views
C4070254|Should-R XR GE 2V
C4070254|Views GE 2:Finding:Point in time:Shoulder.right:Document:XR
C4070254|Views GE 2:Find:Pt:Shoulder.right:Doc:XR
C4070249|Abdominal Aorta US for screening
C4070249|Abd Aorta US Screening
C4070249|Multisection for screening:Finding:Point in time:Abdomen>Aorta.abdominal:Document:Ultrasound
C4070249|Multisection for screening:Find:Pt:Abdomen>Aorta.abdominal:Doc:US
C4070459|Multisection 3D post processing^WO contrast:Finding:Point in time:Chest:Document:Computerized Tomography
C4070459|Chest CT 3D post processing WO contrast
C4070459|Multisection 3D post processing^WO contrast:Find:Pt:Chest:Doc:CT
C4070459|Chest CT p 3D proc WO contr
C4070457|Chest+Abd+Pelvis CT p 3D proc WO contr
C4070457|Chest and Abdomen and Pelvis CT 3D post processing WO contrast
C4070457|Multisection 3D post processing^WO contrast:Finding:Point in time:Chest+Abdomen+Pelvis:Document:Computerized Tomography
C4070457|Multisection 3D post processing^WO contrast:Find:Pt:Chest+Abdomen+Pelvis:Doc:CT
C4071754|Deprecated Spine CT.Dens WO contr
C4071754|Deprecated Spine CT densitometry WO contrast
C4071754|Multisection^WO contrast:Finding:Point in time:Spine:Document:Computerized Tomography.densitometry
C4071754|Multisection^WO contrast:Find:Pt:Spine:Doc:CT.densitometry
C4070478|Chest Pulmonary arteries CT angiogram for pulmonary embolus W contrast IV
C4070478|Chst Pulm art CT.Angio for PE W contr IV
C4070478|Multisection for pulmonary embolus^W contrast Intravenous:Finding:Point in time:Chest>Pulmonary arteries:Document:Computerized Tomography.angio
C4070478|Multisection for pulmonary embolus^W contrast IV:Find:Pt:Chest>Pulmonary arteries:Doc:CT.angio
C4070256|Views GE 2:Find:Pt:Sacrum+Coccyx:Doc:XR
C4070256|Sacrum and Coccyx X-ray GE 2 views
C4070256|Views GE 2:Finding:Point in time:Sacrum+Coccyx:Document:XR
C4070256|Sacrum+Coccyx XR GE 2V
C4070464|Thoracic spine CT by reconstruction WO contrast
C4070464|T-spine CT by reconstr WO contr
C4070464|Multisection by reconstruction^WO contrast:Find:Pt:Spine.thoracic:Doc:CT
C4070464|Multisection by reconstruction^WO contrast:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography
C4070463|Thoracic spine CT densitometry WO contrast
C4070463|Multisection^WO contrast:Find:Pt:Spine.thoracic:Doc:CT.densitometry
C4070463|T-spine CT.Dens WO contr
C4070463|Multisection^WO contrast:Finding:Point in time:Spine.thoracic:Document:Computerized Tomography.densitometry
C4070489|Abdomen CT 3D post processing WO contrast
C4070489|Multisection 3D post processing^WO contrast:Find:Pt:Abdomen:Doc:CT
C4070489|Multisection 3D post processing^WO contrast:Finding:Point in time:Abdomen:Document:Computerized Tomography
C4070489|Abd CT p 3D proc WO contr
C4070481|Kid+Uret+Blad CT p 3D proc WO+W contr IV
C4070481|Multisection 3D post processing^WO & W contrast Intravenous:Finding:Point in time:Abdomen+Pelvis>Kidney+Ureter+Urinary Bladder:Document:Computerized Tomography
C4070481|Kidney+Ureter+Urinary bladder CT 3D post processing WO and W contrast IV
C4070481|Multisection 3D post processing^WO & W contrast IV:Find:Pt:Abdomen+Pelvis>Kidney+Ureter+Urinary Bladder:Doc:CT
C4070480|Pelvis CT by reconstruction W contrast IV
C4070480|Multisection by reconstruction^W contrast IV:Find:Pt:Pelvis:Doc:CT
C4070480|Multisection by reconstruction^W contrast Intravenous:Finding:Point in time:Pelvis:Document:Computerized Tomography
C4070480|Pelvis CT by reconstr W contr IV
C4071447|Ft XR 3V stand
C4071447|Views 3^standing:Finding:Point in time:Foot:Document:XR
C4071447|Foot X-ray 3 views standing
C4071447|Views 3^standing:Find:Pt:Foot:Doc:XR
C4070251|Views GE 4:Finding:Point in time:Spine.lumbar+Sacrum:Document:XR
C4070251|Views GE 4:Find:Pt:Spine.lumbar+Sacrum:Doc:XR
C4070251|L-spine+Sacrum XR GE 4V
C4070251|Spine Lumbar and Sacrum X-ray GE 4 views
C4071449|Views GE 3:Find:Pt:Elbow:Doc:XR
C4071449|Elbow X-ray GE 3 views
C4071449|Elbow XR GE 3V
C4071449|Views GE 3:Finding:Point in time:Elbow:Document:XR
C0411971|X-ray soft tissue
C0411971|x-ray of soft tissue
C0411971|x-ray of soft tissue (procedure)
C0411971|Soft tissue X-ray NOS (procedure)
C0411971|Soft tissue X-ray NOS
C0411971|Soft tissue X-ray
C0411971|Diagnostic radiography of soft tissues (procedure)
C0411971|Diagnostic radiography of soft tissues
C0411971|Diagnostic radiography of soft tissues, NOS
C2017439|X-ray soft tissue calcifications
C2017439|x-ray of soft tissue: calcifications (procedure)
C2017439|x-ray of soft tissue: calcifications
C2017440|X-ray soft tissue gas
C2017440|x-ray of soft tissue: gas
C2017440|x-ray of soft tissue: gas (procedure)
C3161830|x-ray soft tissue calcifications arterial (procedure)
C3161830|x-ray soft tissue calcifications arterial
C0411990|Soft tissue X-ray nose (procedure)
C0411990|Soft tissue X-ray nose
C0559516|Trunk soft tissue X-ray
C0559516|Trunk soft tissue X-ray (procedure)
C0202678|Soft tissue X-ray of face, head AND neck (procedure)
C0202678|Soft tissue X-ray of face, head AND neck
C0202678|Soft tissue X-ray of face, head and neck, NOS
C0202678|Soft tissue x-ray of face, head, and neck
C0412041|Dynamic soft palate study
C0412041|Video soft palate
C0412041|Video soft palate (procedure)
C0203285|Radiography of soft tissue of ankle
C0203285|Radiography of soft tissue of ankle (procedure)
C0203269|Radiography of soft tissue of hip
C0203269|Radiography of soft tissue of hip (procedure)
C0373142|Radiologic examination; neck, soft tissue
C0373142|RADIOLOGIC EXAMINATION NECK SOFT TISSUE
C0373142|X-ray of soft tissue of neck
C0373142|Neck soft tissue X-ray
C0373142|Soft tissue X-ray neck NOS
C0373142|Neck soft tissue X-ray (procedure)
C0373142|Soft tissue X-ray neck NOS (procedure)
C0373142|X-RAY EXAM OF NECK
C0411976|Soft tissue X-ray limbs NOS (procedure)
C0411976|Soft tissue X-ray limbs (procedure)
C0411976|Soft tissue X-ray limbs
C0411976|Soft tissue X-ray limbs NOS
C0411987|Head soft tissue X-ray
C0411987|Head soft tissue X-ray (procedure)
C0203225|Radiography of soft tissue of shoulder
C0203225|Radiography of soft tissue of shoulder (procedure)
C0559518|Vascular soft tissue X-ray
C0559518|Vascular soft tissue X-ray (procedure)
C1536645|Imaging - soft tissue
C1536645|Tissue imaging - soft
C1536645|Soft tissue imaging
C1536645|Soft tissue imaging (& plain) (procedure)
C1536645|Soft tissue imaging - plain
C1536645|Soft tissue imaging (& plain)
C0203197|Radiography of pelvic soft tissue
C0203197|Radiography of pelvic soft tissue (procedure)
C0203233|Radiography of soft tissue of elbow
C0203233|Radiography of soft tissue of elbow (procedure)
C0203239|Radiography of soft tissue of forearm
C0203239|Radiography of soft tissue of forearm (procedure)
C0203248|Radiography of soft tissue of hand
C0203248|Hand soft tissue X-ray
C0203248|Radiography of soft tissue of hand (procedure)
C0203277|Radiography of soft tissue of knee
C0203277|Radiography of soft tissue of knee (procedure)
C0411975|Soft tissue X-ray lymph nodes
C0411975|Soft tissue X-ray lymph nodes (procedure)
C0411972|Postmortem radiology - soft tissue (procedure)
C0411972|Postmortem radiology - soft tissue
C0411972|Postmortem radiographic imaging of soft tissue (procedure)
C0411972|Postmortem radiographic imaging of soft tissue
C0034589|Dilution Technic, Radioisotope
C0034589|Dilution Technics, Radioisotope
C0034589|Dilution Technique, Radioisotope
C0034589|Dilution Techniques, Radioisotope
C0034589|Radioisotope Dilution Technics
C0034589|Radioisotope Dilution Technique
C0034589|Radioisotope Dilution Techniques
C0034589|Technic, Radioisotope Dilution
C0034589|Technics, Radioisotope Dilution
C0034589|Technique, Radioisotope Dilution
C0034589|Techniques, Radioisotope Dilution
C0034589|isotope dilution method
C0034589|Radioisotope Dilution Technic
C0004400|Autoradiography
C0004400|RADIOAUTOGR
C0004400|AUTORADIOGR
C0004400|radioautography
C0008797|Cinefluorographies
C0008797|Cineradiographies
C0008797|Cineradiography
C0008797|Radiocinematographies
C0008797|cinefluorography
C0008797|CINEFLUOROGR
C0008797|CINERADIOGR
C0008797|RADIOCINEMATOGR
C0008797|Cineradiography NOS
C0008797|Movement radiogr.
C0008797|(Cineradiography) or (movement radiography)
C0008797|(Cineradiography) or (movement radiography) (procedure)
C0008797|Cineradiography NOS (procedure)
C0008797|Movement radiography
C0008797|Cineradiography (procedure)
C0008797|Radiocinematography
C0008797|Movement radiography (procedure)
C0008797|Cineradiography, NOS
C0008797|videofluorography
C0034575|Radiography, Dental
C0034575|dental radiography
C0034575|DENT RADIOGR
C0034575|RADIOGR DENT
C0034575|X-ray teeth
C0034575|x-ray of teeth
C0034575|x-ray of teeth (procedure)
C0034575|X-ray dental
C0034575|Dental X-ray (procedure)
C0034575|Dental X-ray
C0034575|Plain X-ray teeth NOS (procedure)
C0034575|Plain X-ray teeth NOS
C0034575|Plain X-ray teeth
C0034575|Radiography of teeth
C0034575|Radiography of teeth (procedure)
C0034575|Radiography of teeth, NOS
C0034575|X-ray;dental
C0016356|Fluoroscopies
C0016356|Fluoroscopy
C0016356|Fluoroscopic imaging - action
C0016356|Fluoroscopic imaging
C0016356|fluoroscopy (procedure)
C0016356|Fluoroscopy NOS
C0016356|Fluoroscopy NOS (procedure)
C0016356|Fluoroscopic imaging procedure (procedure)
C0016356|Fluoroscopy technique
C0016356|Fluoroscopic imaging - action (qualifier value)
C0016356|Fluoroscopy, NOS
C0024671|Mammographies
C0024671|Mammography
C0024671|Mammogram
C0024671|MAMMOGR
C0024671|mammogram (procedure)
C0024671|Mam
C0024671|Mammography (procedure)
C0024671|Radiographic examination of breast
C0024671|Mammography, NOS
C0024671|Radiographic examination of breast, NOS
C0024671|Mammogram, NOS
C0026015|Microradiography
C0026015|Microradiographies
C0026015|MICRORADIOGR
C0000853|Absorptiometry, Photon
C0000853|photon absorptiometry
C0040395|Tomographies
C0040395|Tomography
C0040395|TOMOGR
C0040395|Tomographic imaging procedure
C0040395|Tomography (procedure)
C0040395|Tomographic imaging
C0040395|Tomography - NOS
C0040395|Tomography - NOS (procedure)
C0040395|Tomographic imaging, plain radiologic - action (qualifier value)
C0040395|Tomograms
C0040395|Diagnostic tomography
C0040395|Diagnostic tomographic examination
C0040395|Diagnostic laminographic examination
C0040395|Diagnostic tomography (procedure)
C0040395|Tomogram
C0040395|Tomographic imaging - action (qualifier value)
C0040395|Tomographic imaging - action
C0040395|Tomographic imaging procedure (procedure)
C0040395|Tomographic imaging, plain radiologic - action
C0040395|Diagnostic tomography, NOS
C0040395|Diagnostic laminographic examination, NOS
C0040395|Diagnostic tomographic examination, NOS
C0597348|radiocardiography
C0597511|stereoradiography
C0001780|Age Determination by Skeleton
C0002978|Angiographies
C0002978|Angiography
C0002978|ANGIOGR
C0002978|angiography (procedure)
C0002978|Angiogram
C0002978|Angiogram NOS
C0002978|Angiograph
C0002978|Diagnostic angiogram
C0002978|Diagnostic angiography
C0002978|Angiography, NOS
C0002978|Angiogram, NOS
C0003885|Arthrographies
C0003885|Arthrography
C0003885|Arthrogram
C0003885|ARTHROGR
C0003885|Contrast arthrogram
C0003885|Arthrography NOS (procedure)
C0003885|Arthrography NOS
C0003885|Arthrograph
C0003885|Joint X-ray study
C0003885|Arthrography (procedure)
C0003885|Arthrography, NOS
C0003885|Arthrogram, NOS
C0013828|Electrokymographies
C0013828|Electrokymography
C0013828|Kymographies, Radiographic
C0013828|Radiographic Kymographies
C0013828|Roentgenkymographies
C0013828|RADIOGR KYMOGR
C0013828|KYMOGR RADIOGR
C0013828|ROENTGENKYMOGR
C0013828|ELECTROKYMOGR
C0013828|Kymography, Radiographic
C0013828|Radiographic Kymography
C0013828|Roentgenkymography
C0020709|Hysterosalpingographies
C0020709|Hysterosalpingography
C0020709|Hysterosalpingogram
C0020709|HYSTEROSALPINGOGR
C0020709|HSG (hysterosalpingogram)
C0020709|hysterosalpingography (procedure)
C0020709|X-ray hysterosalpingography
C0020709|Hysterosalpingogram (procedure)
C0020709|Hysterosalpingography NOS (procedure)
C0020709|Hysterosalpingography NOS
C0020709|Salp - Hysterosalpingogram
C0020709|HSG - Hysterosalpingogram
C0020709|Hysterosalpingography, NOS
C0020709|Hysterosalpingography (procedure) [Ambiguous]
C0024290|Lymphographies
C0024290|Lymphography
C0024290|LYMPHOGR
C0027904|Neuroradiography
C0027904|Neuroradiographies
C0027904|NEURORADIOGR
C0032323|Air Radiographies
C0032323|Contrast Radiographies, Negative
C0032323|Insufflation Radiographies
C0032323|Negative Contrast Radiographies
C0032323|Pneumoradiographies
C0032323|Pneumoradiography
C0032323|Radiographies, Air
C0032323|Radiographies, Insufflation
C0032323|Radiographies, Negative Contrast
C0032323|INSUFFLATION RADIOGR
C0032323|RADIOGR AIR
C0032323|CONTRAST RADIOGR NEGATIVE
C0032323|AIR RADIOGR
C0032323|RADIOGR INSUFFLATION
C0032323|RADIOGR NEGATIVE CONTRAST
C0032323|PNEUMORADIOGR
C0032323|NEGATIVE CONTRAST RADIOGR
C0032323|Radiography, Insufflation
C0032323|Negative Contrast Radiography
C0032323|Radiography, Air
C0032323|Radiography, Negative Contrast
C0032323|Air Radiography
C0032323|Contrast Radiography, Negative
C0032323|Insufflation Radiography
C0034564|Enhancement, Radiographic Image
C0034564|Enhancements, Radiographic Image
C0034564|Image Enhancements, Radiographic
C0034564|Radiographic Image Enhancement
C0034564|Radiographic Image Enhancements
C0034564|RADIOGR IMAGE ENHANCEMENT
C0034564|IMAGE ENHANCEMENT RADIOGR
C0034564|Image Enhancement, Radiographic
C0034568|Magnifications, Radiographic
C0034568|Radiographic Magnification
C0034568|Radiographic Magnifications
C0034568|RADIOGR MAGNIFICATION
C0034568|MAGNIFICATION RADIOGR
C0034568|Magnification, Radiographic
C0034573|Radiography, Abdominal
C0034573|Abdominal Radiographies
C0034573|Radiographies, Abdominal
C0034573|Abdominal X-Ray
C0034573|RADIOGR ABDOMINAL
C0034573|ABDOMINAL RADIOGR
C0034573|x-ray of abdomen (procedure)
C0034573|x-ray of abdomen
C0034573|X-ray;abdomen
C0034573|Abdominal X-ray (procedure)
C0034573|Radiologic examination, abdomen
C0034573|Abdomen--Radiography
C0034573|Abdominal X-ray NOS
C0034573|Abdominal Radiography
C0034573|AXR - Abdominal X-ray
C0034573|Diagnostic radiography of abdomen (procedure)
C0034573|Diagnostic radiography of abdomen
C0034573|Radiologic examination of abdomen
C0034573|Radiologic procedure on abdomen
C0034573|Radiologic examination of abdomen, NOS
C0034573|X-ray of abdomen, NOS
C0034573|Radiologic procedure on abdomen, NOS
C0034573|X-ray of the abdomen
C3665494|Radiographies, Thoracic
C3665494|Radiography, Thoracic
C3665494|Thoracic Radiographies
C3665494|Thoracic Radiography
C3665494|THORACIC RADIOGR
C3665494|RADIOGR THORACIC
C3665494|Radiologic examination of chest
C3665494|X-ray thoracic cage NOS (procedure)
C3665494|Radiographic procedure on chest (procedure)
C3665494|X-ray thoracic cage NOS
C3665494|Thoracic cage X-ray
C3665494|Thoracic cage X-ray (procedure)
C3665494|Radiographic procedure on chest
C3665494|CXR - Chest X-ray
C3665494|Chest x-ray
C3665494|Radiography of chest
C3665494|Thorax X-ray
C0040404|Tomography, X-Ray
C0040404|RADIOGR TOMOGR
C0040404|TOMOGR X RAY
C0040404|TOMOGR RADIOGR
C0040404|TOMOGR XRAY
C0040404|ZONOGR
C0040404|X RAY TOMOGR
C0040404|TOMOGR TRANSM
C0040404|XRAY TOMOGR
C0040404|TRANSM TOMOGRAPHY
C0040404|X-ray tomography (procedure)
C0040404|X-ray tomography
C0040404|X Ray Tomography
C0040404|Tomography, X Ray
C0040404|Tomography, Radiographic
C0040404|Tomography, Xray
C0040404|Xray Tomography
C0040404|Transmission Tomography
C0040404|Radiographic Tomography
C0040404|Tomography, Transmission
C0040404|Zonography
C0040404|Zonography (procedure)
C0042070|Urography
C0042070|UROGR
C0042070|Urogram
C0043350|Xeroradiographies
C0043350|Xeroradiography
C0043350|XERORADIOGR
C0043350|xerography
C0043350|xeroradiography (procedure)
C0043350|Xeroradiography, NOS
C0043350|Xerography, NOS
C1962945|Radiography
C1962945|Radiology
C1962945|RADIOGR
C1962945|Radiographic imaging procedure
C1962945|Medical Imaging, X-Ray
C1962945|Conventional X-Ray
C1962945|X-Ray Imaging
C1962945|XR
C1962945|Roentgenography
C1962945|X-ray
C1962945|radiographic imaging procedure (procedure)
C0034565|Radiographic Image Interpretation, Computer-Assisted
C0034565|RADIOGR IMAGE INTERP COMPUTER ASSISTED
C0034565|RADIOGR IMAGE INTERP
C0034565|COMPUTER ASSISTED RADIOGR IMAGE INTERP
C0034565|Computer Assisted Radiographic Image Interpretation
C0034565|Radiographic Image Interpretation, Computer Assisted
C0034565|Computer-Assisted Radiographic Image Interpretation
C0034578|Radiography, Interventional
C0034578|RADIOGR INTERVENTIONAL
C0034578|INTERVENTIONAL RADIOGR
C0034578|Interventional Radiography
C1956099|Sex Determination by Skeleton
C2183262|diagnostic service sources radiology labs X-ray (procedure)
C2183262|x-ray department
C2183262|Diagnostic service sources - radiology labs X-ray
C2183262|diagnostic service sources radiology labs x-ray
C2585137|Parallel beam scanography (procedure)
C2585137|Parallel beam scanography
C0411842|Postmortem radiology NOS (procedure)
C0411842|Postmortem radiology (procedure)
C0411842|Postmortem radiology NOS
C0411842|Postmortem radiology
C0411842|Postmortem radiographic imaging
C0411842|Postmortem radiographic imaging (procedure)
C0411831|Stereographic radiogr.
C0411831|Stereographic radiography
C0411831|Stereographic radiography (procedure)
C3178874|Radiostereometric Analysis
C3178874|Analysis, Radiostereometric
C3178874|Analyses, Radiostereometric
C3178874|Stereophotogrammetry, Roentgen
C3178874|Radiostereometric Analyses
C3178874|radiostereometric analysis (procedure)
C3178874|Roentgen Stereophotogrammetry
C3178874|Radiostereometry
C3272922|Total Body Radiography
C0473880|Esophageal radiological intervention
C0473880|Oesophageal radiological intervention
C0473880|Oesophageal intervention
C0473880|Esophageal intervention
C0473880|Esophageal intervention (procedure)
C0202616|Radiologic examination, osseous survey; complete (axial and appendicular skeleton)
C0202616|RADIOLOGIC EXAMINATION OSSEOUS SURVEY COMPL
C0202616|Radiologic examination, osseous survey, complete
C0202616|Skeletal survey
C0202616|Skeletal series x-ray
C0202616|complete osseous survey (procedure)
C0202616|complete osseous survey
C0202616|X-RAYS BONE SURVEY COMPLETE
C0202616|X-ray: skeletal survey NOS (procedure)
C0202616|Skeletal X-ray
C0202616|Skeletal X-ray (procedure)
C0202616|X-ray: skeletal survey NOS
C0202616|Skeletal X-ray (& general survey) (procedure)
C0202616|X-ray: general skeletal survey
C0202616|Skeletal X-ray (& general survey)
C0202616|X-ray of whole skeleton
C0202616|Radiography for bone survey
C0202616|Complete skeletal series
C0202616|Skeletal series
C0202616|Radiographic skeletal survey
C0202616|Skeletal survey X-ray
C0202616|Radiologic examination, osseous survey, complete (procedure)
C0202616|Skeletal X-ray, NOS
C0202616|Skeletal series, NOS
C0202616|Skeletal survey, NOS
C0579019|Transesophageal aortography
C0579019|Transoesophageal aortography
C0579019|Transesophageal aortography (procedure)
C0400529|Endoscopic retrograde pancreatography and collection of pancreatic juice
C0400529|Endoscopic retrograde pancreatography and collection of pancreatic juice (procedure)
C1261034|Unilateral imaging of coronary artery with recording (situation)
C1261034|Unilateral imaging of coronary artery with recording
C1261034|Coronary angiography, unilateral selective injection includes angiogram and recording (procedure)
C1261034|Coronary angiography, unilateral selective injection includes angiogram and recording
C0013518|ECHOCARDIOGR CONTRAST
C0013518|CONTRAST ECHOCARDIOGR
C0013518|Contrast echocardiography (procedure)
C0013518|Contrast echocardiography
C0013518|Contrast echocardiography procedure
C0013518|Echocardiography, Contrast
C0203067|Radiologic examination of pharynx and cervical esophagus
C0203067|Radiologic examination of pharynx and cervical oesophagus
C0203067|Radiologic examination of pharynx and cervical esophagus (procedure)
C1285406|Radiologic guidance for diagnostic procedure (procedure)
C1285406|Radiologic guidance for diagnostic procedure
C0581644|Plain film by body site (procedure)
C0581644|Plain film by body site
C0581644|Plain film of body region
C0581644|Plain film of body region (procedure)
C0438940|Percutaneous transluminal vertebral artery balloon angioplasty
C0438940|percutaneous transluminal angioplasty of vertebral artery
C0438940|percutaneous transluminal angioplasty of vertebral artery (treatment)
C0438940|Percutaneous transluminal vertebral artery balloon angioplasty (procedure)
C0438940|PTA of head and neck arteries, vertebral
C0411822|Stereotactic/stereoscopic test - soft tissue (procedure)
C0411822|Stereotactic/stereoscopic test - soft tissue
C0202848|Radiographic procedure on cardiovascular system (procedure)
C0202848|Radiographic procedure on cardiovascular system
C0202848|Radiologic procedure on cardiovascular system
C2732671|Radiologic intervention on respiratory tract (procedure)
C2732671|Radiologic intervention on respiratory tract
C2732671|Respiratory tract intervention
C2732671|Respiratory tract intervention (procedure)
C2732671|Respiratory tract radiological intervention
C0456899|X-ray guided biopsy
C0456899|X-ray guided biopsy (procedure)
C0344093|Interventional Radiology Procedure
C0344093|Interventional radiologic procedures
C0344093|Interventional radiology
C0344093|Interventional radiology (procedure)
C1285361|Musculoskeletal system diagnostic imaging procedure (procedure)
C1285361|Musculoskeletal system diagnostic imaging procedure
C2733119|Radiologic intervention on gastrointestinal tract (procedure)
C2733119|Radiologic intervention on gastrointestinal tract
C2733119|Gastrointestinal tract radiological intervention
C2733119|Gastrointestinal tract intervention
C2733119|Gastrointestinal tract intervention (procedure)
C0581425|CT of regions (procedure)
C0581425|Computed tomography of regions (procedure)
C0581425|Computed tomography of regions
C0581425|CT of regions
C0202640|fluoroscopy and radiography (procedure)
C0202640|fluoroscopy and radiography
C0202640|Fluoroscopy and radiography NOS
C0202640|Fluoroscopy and radiography NOS (procedure)
C0202640|Diagnostic radiologic examination with fluoroscopy
C0202640|Fluoroscopic monitoring with radiography
C0202640|Fluoroscopy of regions
C0202640|Diagnostic radiologic examination with fluoroscopy (procedure)
C0202640|Fluoroscopy of regions (procedure)
C0684210|Diagnostic imaging and nuclear medicine procedures
C0684210|Diagnostic imaging and nuclear medicine procedures (procedure)
C0684210|Diagnostic imaging and nuclear medicine procedures (navigational concept)
C0039985|Chest X-ray
C0039985|chest X ray
C0039985|chest radiography
C0039985|CXR
C0039985|chest xray
C0039985|x-ray of chest (procedure)
C0039985|x-ray of chest
C0039985|X-ray;chest
C0039985|Radiography of chest
C0039985|Radiography of chest (procedure)
C0039985|Radiologic examination of chest
C0039985|Chest exclusion X-ray
C0039985|CXR - Chest X-ray
C0039985|Radiologic examination, chest
C0039985|Radiologic examination
C0039985|Chest--Radiography
C0039985|Plain chest X-ray
C0039985|X-ray NOS chest
C0039985|Plain chest X-ray (procedure)
C0039985|Radiography of chest, NOS
C0039985|Radiologic examination of chest, NOS
C0039985|Chest x-ray, NOS
C0039985|thoracic radiography
C0039985|X-ray of chest NOS
C0202888|Percutaneous transluminal balloon angioplasty of renal artery
C0202888|Percutaneous transluminal renal artery balloon angioplasty
C0202888|Percutaneous transluminal renal artery balloon angioplasty (procedure)
C0436374|Radiology - general (context-dependent category)
C0436374|Radiology - general NOS (context-dependent category)
C0436374|Radiology - general NOS
C0436374|Radiology - general NOS (procedure)
C0436374|Radiology - general
C0436374|Radiology - general (procedure)
C0436374|Radiology - general NOS (situation)
C0436374|Radiology - general (situation)
C0848630|Radiographic imaging of bone (procedure)
C0848630|Radiographic imaging of bone
C0848630|X-ray of bone
C0848630|Plain X-ray of bone
C0848630|X-ray of bone (procedure)
C0848630|Plain X-ray;bone(s)
C0848630|X-ray;bone(s)
C0848630|X-ray of bones
C0848630|Plain bone X-ray NOS
C0848630|Plain bone X-ray NOS (procedure)
C0848630|plain X-ray of the bone(s)
C0848630|bone xray
C0542435|Contrast radiography NOS (procedure)
C0542435|Contrast radiography NOS
C0542435|Diagnostic radiography with contrast media
C0542435|diagnostic radiography with contrast media (procedure)
C0542435|Diagnostic radiologic examination with contrast media
C0542435|Contrast radiography
C0542435|Contrast radiology
C0542435|Contrast radiology excluding angiography
C0542435|Diagnostic radiography with contrast media, NOS
C0542435|Diagnostic radiologic examination with contrast media, NOS
C1976630|Miscellaneous systems
C0005898|Body Regions
C0005898|Body Region
C0005898|Region, Body
C0005898|Regions, Body
C0005898|Anatomic Region
C0005898|ANTREG
C0005898|Body region structure
C0005898|Topographic region
C0005898|Body region structure (body structure)
C0005898|Topographic region, NOS
C0005898|Anatomic region, NOS
C0005898|Body region, NOS
C0015965|Fetus
C0015965|Fetal
C0015965|fetuses
C0015965|^Fetus
C0015965|Fetus (person)
C0370003|Sample
C0370003|Specimen
C0370003|Specimen (specimen)
C0370003|Research Specimen
C1987595|Exhaled gas &#x7C; Radnuc
C0460002|body system
C0460002|Body system -RETIRED-
C0460002|Body systems
C0460002|Body system (body structure)
C0460002|BODSYS
C0460002|Body system structure
C0460002|Organ system
C0460002|Body system structure (body structure)
C0460002|Body apparatus, NOS
C0460002|Body system, NOS
C3887560|Devices
C3887560|Radiology Devices
C0175730|TUBE
C0175730|Tube, device
C0175730|Tube, device (physical object)
C0175730|Tube, NOS
C0175730|biomedical tube device
C0030705|Patient
C0030705|Patients
C0030705|PT
C0030705|*^patient
C0030705|^Patient
C0030705|LAY USER/PATIENT
C0030705|Patient (person)
C3668859|Radiologic examination
C3668859|Radiologic examination of the Gastrointestinal Tract
C4027283|x-ray of shunt (procedure)
C4027283|x-ray of shunt
C3861026|x-ray foreign body
C3861026|x-ray of foreign body
C3861026|x-ray of foreign body (procedure)
C4027281|x-ray of unilateral ribs with chest, three or more views and PA chest views (procedure)
C4027281|x-ray of unilateral ribs with chest, three or more views and PA chest views
C4027281|x-ray unilateral ribs + chest 3+ views + posteroanterior chest
C4027963|portable x-ray of unilateral ribs with chest three or more views and PA chest views
C4027963|portable x-ray of unilateral ribs with chest three or more views and posteroanterior chest views
C4027963|portable x-ray of unilateral ribs with chest three or more views and PA chest views (procedure)
C4027272|x-ray with manual stress (procedure)
C4027272|x-ray with manual stress
C4029665|x-ray comparison view
C4029665|comparison view x-ray (procedure)
C4029665|comparison view x-ray
C4027868|radiographic imaging upper gastrointestinal tract (procedure)
C4027868|radiographic imaging upper gastrointestinal tract
C0011926|Diagnostic radiography with measurements
C0011926|Diagnostic radiography with measurements (procedure)
C0202586|Diagnostic radiography, survey
C0202586|Diagnostic radiography, survey (procedure)
C0202586|Diagnostic radiography, survey, NOS
C0203661|Multi-plane radionuclide tomography
C0203661|Multi-plane radionuclide tomography (procedure)
C0203661|Multi-plane radionuclide tomography, NOS
C0337380|Endoscopic retrograde pancreatography
C0337380|x-ray gastrointestinal EPR
C0337380|endoscopic retrograde pancreatography (procedure)
C0337380|Endosc retro pancreatog
C0337380|Diagnostic endoscopic retrograde examination of pancreatic duct NOS (procedure)
C0337380|Diagnostic endoscopic retrograde examination of pancreatic duct NOS
C0337380|ERP
C0337380|ERP - Endoscopic retrograde pancreatography
C0337380|Diagnostic endoscopic retrograde examination of pancreatic duct
C0337380|Endoscopic retrograde pancreatography [ERP]
C0202576|Diagnostic radiography, stereo
C0202576|Diagnostic radiography, stereo (procedure)
C0202577|Diagnostic radiography, stereotactic localization
C0202577|Diagnostic radiography, stereotactic localisation
C0202577|Diagnostic radiography, stereotactic localization (procedure)
C0202585|Diagnostic radiography for foreign body detection and localization
C0202585|Diagnostic radiography for foreign body detection and localisation
C0202585|Diagnostic radiography for foreign body detection and localization (procedure)
C0202613|Fistulogram
C0202613|Fistulogram (procedure)
C0202613|Diagnostic radiography of fistula or sinus tract, positive contrast
C0202613|Diagnostic radiography of fistula or sinus tract, positive contrast (procedure)
C1306645|Radiograph
C1306645|Radiogram
C1306645|X-ray
C1306645|x-ray (procedure)
C1306645|Plain film (procedure)
C1306645|Plain radiography (procedure)
C1306645|Plain film
C1306645|Plain radiography
C1306645|Plain film diagnostic procedure (procedure)
C1306645|Plain film diagnostic procedure
C1306645|X-rays
C1306645|Radiographs
C1306645|X-ray NOS
C1306645|Roentgenography
C1306645|Roentgenogram
C1306645|Skiagram
C1306645|Plain x-ray
C0040405|CAT Scans, X-Ray
C0040405|Computed Tomography, Xray
C0040405|Computed X-Ray Tomography
C0040405|CT X Rays
C0040405|Scan, X-Ray CAT
C0040405|Scans, X-Ray CAT
C0040405|Tomographies, Computed X-Ray
C0040405|Tomography, Computed X-Ray
C0040405|Tomography, X-Ray Computed
C0040405|X Ray, CT
C0040405|X Rays, CT
C0040405|X-Ray CAT Scan
C0040405|X-Ray CAT Scans
C0040405|X-Ray Computed Tomography
C0040405|X-Ray Computerized Tomography
C0040405|Xray Computed Tomography
C0040405|CAT scan
C0040405|computed axial tomography
C0040405|CT
C0040405|Computerized Tomography
C0040405|Computerized axial tomography scan - NOS (procedure)
C0040405|CT XRAY
C0040405|CT scan
C0040405|EMI scan
C0040405|computerized tomography (procedure)
C0040405|CT (computerized tomography)
C0040405|X Ray Computer Assisted Tomography
C0040405|X-Ray CT Scans
C0040405|Tomography, X Ray Computerized
C0040405|Scans, X-Ray CT
C0040405|Transmission Computed Tomography
C0040405|Tomography, X Ray Computer Assisted
C0040405|Computed Tomography, X Ray
C0040405|CT Scans, X-Ray
C0040405|X-Ray CT Scan
C0040405|CT Scan, X Ray
C0040405|Scan, X-Ray CT
C0040405|Computed Tomography, Transmission
C0040405|TOMOGRAPHY TRANSM COMPUTED
C0040405|Computerised tomogram
C0040405|CTT
C0040405|computed tomography
C0040405|computed tomography (procedure)
C0040405|Computed tomography procedure
C0040405|CAT Scans
C0040405|CT Scans
C0040405|Computerized axial tomography scan - NOS
C0040405|CAT scan - NOS
C0040405|Computed tomography scan - NOS
C0040405|CAT scan - NOS (procedure)
C0040405|Computed tomography scan - NOS (procedure)
C0040405|Computerised axial tomography scan - NOS
C0040405|tomography
C0040405|computerized axial tomography
C0040405|Computerized transverse axial tomography
C0040405|Computerized transverse axial tomogram
C0040405|Computerised axial tomogram
C0040405|Computerised axial tomography
C0040405|CTT scan
C0040405|CAT
C0040405|Computer-assisted transaxial tomography
C0040405|Computerized axial tomogram
C0040405|Computerised tomography
C0040405|Computerised transverse axial tomogram
C0040405|Computerised transverse axial tomography
C0040405|Computerized tomogram
C0040405|X-Ray Computer Assisted Tomography
C0040405|X Ray Tomography, Computed
C0040405|CAT Scan, X Ray
C0040405|Computerized Tomography, X-Ray
C0040405|X-Ray Tomography, Computed
C0040405|Computed X Ray Tomography
C0040405|Tomography, X-Ray Computerized
C0040405|X Ray Computerized Tomography
C0040405|CT Scan, X-Ray
C0040405|CT X Ray
C0040405|Tomodensitometry
C0040405|Tomography, X-Ray Computer Assisted
C0040405|CAT Scan, X-Ray
C0040405|Tomography, Transmission Computed
C0040405|Tomography, X Ray Computed
C0040405|Tomography, Xray Computed
C0040405|Computerized Tomography, X Ray
C0040405|Computed Tomography, X-Ray
C0040405|Computerized transaxial tomography
C0040405|CAT - Computerised axial tomography
C0040405|CAT - Computerized axial tomography
C0040405|CT - Computerised tomography
C0040405|CT - Computerized tomography
C0040405|Computerised tomograph scan
C0040405|Computerized tomograph scan
C0040405|Computerised transaxial tomography
C0040405|Computerized axial tomography (procedure)
C0040405|tomography, computed
C0040405|Computerized axial tomography, NOS
C0040405|Computerized transaxial tomography without IV contrast
C0040405|Computerized tomography without IV contrast
C0040405|CT scan without IV contrast
C0040405|CAT scan, NOS
C0040405|Computerized transaxial tomography, NOS
C0040405|C.A.T. scan NOS
C0524310|Intra-arterial digital subtraction angiography
C0524310|Intra-arterial DSA
C0524310|Intra-arterial digital subtraction angiography (procedure)
C0524311|Intravenous DSA
C0524311|Intravenous digital subtraction angiography
C0524311|Intravenous digital subtraction angiography (procedure)
C0412204|Pneumocystogram
C0412204|Pneumocystogram (procedure)
C0412209|Tenogram
C0412209|Tenogram (procedure)
C0412006|Whole body X-ray of stillborn infant
C0412006|Whole body X-ray of stillborn infant (procedure)
C0412004|X-ray of pathological specimen (procedure)
C0412004|X-ray of pathological specimen
C0581651|Specific plain X-ray investigations
C0581651|Specific plain X-ray investigations (procedure)
C0581652|Plain X-ray imaging - action
C0581652|Plain X-ray imaging
C0581652|Plain X-ray techniques
C0581652|Plain radiography technique
C0581652|Plain X-ray technique
C0581652|Plain X-ray imaging - action (qualifier value)
C0581652|Plain X-ray techniques (procedure)
C0581652|Plain film technique
C0473893|Computerised diagnostic radiology (procedure)
C0473893|Computerised diagnostic radiology NOS
C0473893|Computerised diagnostic radiology
C0473893|Computerised diagnostic radiology NOS (procedure)
C0473893|Computerized diagnostic radiology NOS
C0473893|Computerized diagnostic radiology NOS (procedure)
C0473893|Computerized diagnostic radiology
C0473893|Computerized diagnostic radiology (procedure)
C0202630|Diagnostic radiologic examination with special study
C0202630|Diagnostic radiography with special study (procedure)
C0202630|Diagnostic radiography with special study
C0202630|Diagnostic radiography with special study, NOS
C0202630|Diagnostic radiologic examination with special study, NOS
C1266814|Radiographic imaging procedure by site (procedure)
C1266814|Topography specific radiographic procedure
C1266814|Radiographic imaging procedure by site
C1266814|Topography specific radiographic procedure (procedure)
C1266814|Topography specific radiologic procedure
C0412221|Cardiac shunt study
C0412221|Cardiac shunt study (procedure)
C0032279|Pneumoencephalographies
C0032279|Pneumoencephalography
C0032279|Air Encephalography
C0032279|PNEUMOENCEPHALOGR
C0032279|pneumoencephalography (procedure)
C0032279|X-ray pneumoencephalography
C0032279|Pneumoencephalogram
C0032279|Pneumencephalography
C0032279|Encephalography (Air)
C0032279|Pneumoventriculogram
C0202584|Diagnostic radiography during operative procedure
C0202584|Diagnostic radiography during operative procedure (procedure)
C0193504|Endosc retro cholangio
C0193504|Endoscopic retrograde cholangiography
C0193504|ERC
C0193504|Diagnostic endoscopic retrograde examination of bile duct NOS
C0193504|Diagnostic endoscopic retrograde examination of bile duct NOS (procedure)
C0193504|ERC - Endoscopic retrograde cholangiography
C0193504|Endoscopic retrograde cholangiography (procedure)
C0193504|Diagnostic endoscopic retrograde examination of bile duct
C0193504|Diagnostic endoscopic retrograde examination of bile duct (procedure)
C0193504|ERC, NOS
C0193504|Endoscopic retrograde cholangiography [ERC]
C0401385|Cystoscopy and retrograde pyelography
C0401385|Cystoscopy and retrograde pyelography (procedure)
C0193505|Endoscopic retrograde cholangiopancreatography (ERCP); with biopsy, single or multiple
C0193505|Endoscopic retrograde cholangiopancreatography (ERCP) with biopsy
C0193505|ERCP W/BIOPSY SINGLE/MULTIPLE
C0193505|Endoscopic retrograde cholangiopancreatography with biopsy
C0193505|ERCP with biopsy
C0193505|ERCP with biopsy (procedure)
C0193505|Endoscopic retrograde cholangiopancreatography with biopsy (procedure)
C0193505|ENDO CHOLANGIOPANCREATOGRAPH
C0193527|Laparoscopy with guided transhepatic cholangiography
C0193527|Laparoscopy with guided transhepatic cholangiography (procedure)
C0401387|Ascending ureterogram
C0401387|Blow up ureteropyelogram
C0401387|Cystoscopy and bulb catheter ureteropyelography
C0401387|Cystoscopy and bulb catheter ureteropyelography (procedure)
C0203114|Antegrade pyelogram
C0203114|antegrade pyelogram (procedure)
C0203114|Nephrostogram
C0203114|Loopogram
C0203114|Antegrade urography
C0203114|Nephrostography
C0203114|Nephrostomography
C0203114|Percutaneous pyelogram by direct puncture
C0203114|Tube nephrostogram
C0203114|Antegrade urogram
C0203114|Nephrostogram (procedure)
C0203114|Antegrade urography (procedure)
C0203114|Urinary tract loopogram
C0203114|Fluoroscopic antegrade pyelography (procedure)
C0203114|Fluoroscopic antegrade pyelography
C0203114|Fluoroscopic nephrostography (procedure)
C0203114|Fluoroscopic nephrostography
C0006282|Bronchographies
C0006282|Bronchography
C0006282|Bronchogram
C0006282|BRONCHOGR
C0006282|bronchography (procedure)
C0006282|Contrast bronchogram (procedure)
C0006282|Contrast bronchogram
C0006282|Contrast bronchogram, NOS
C0205917|Renographies
C0205917|RENOGR
C0205917|Renography
C1519363|Small Bowel Follow Through Procedure
C0203057|Upper GI Series
C0203057|Retired procedure (procedure) [P5-50110]
C0203057|Retired procedure [P5-50110]
C0203057|upper gastrointestinal series
C0203057|Barium study of esophagus stomach and duodenum
C0203057|Barium study of oesophagus stomach and duodenum
C0203057|Upper gastrointestinal tract series
C0203057|Upper gastrointestinal tract series (procedure)
C0203057|Barium-Swallow X-ray
C0203057|Upper GI
C0203057|Upper Gastrointestinal Tract Radiography
C0203126|Cystogram
C0203126|Cystography
C0203126|Cystography (procedure)
C0203126|Cystography NOS
C0203126|Cystogram (procedure)
C0203126|Cystography NOS (procedure)
C0203126|Contrast radiography of bladder
C0203126|Cystography, NOS
C0203126|Contrast radiography of bladder, NOS
C0203126|Cystography (procedure) [Ambiguous]
C0203126|Fluoroscopic cystography (procedure)
C0203126|Fluoroscopic cystography
C1519939|Vaginography
C1318509|Oesophagram
C1318509|esophagogram
C1318509|esophagogram (procedure)
C1318509|contrast esophagram
C1318509|esophagram
C1318509|Contrast radiography of esophagus
C1318509|Contrast radiography of oesophagus
C1318509|Contrast radiography of esophagus (procedure)
C1318509|Contrast Esophagraphy
C1318509|Esophagography
C0438653|Portable X-ray (context-dependent category)
C0438653|Portable X-ray (situation)
C0438653|Portable X-ray
C0438653|Portable X-ray (procedure)
C0412765|X-ray photon absorptiometry
C0412765|X-ray photon absorptiometry (procedure)
C1998274|Radiopharmaceutical imaging (procedure)
C1998274|Radiopharmaceutical imaging
C0026995|Myelographies
C0026995|Myelography
C0026995|Myelogram
C0026995|MYELOGR
C0026995|myelography (procedure)
C0026995|Contrast myelogram
C0026995|Myelogram (procedure)
C0026995|Spinal myelogram
C0026995|Spinal myelograph
C0026995|Myelograph spinal
C0026995|Myelogram, NOS
C0026995|Myelography, NOS
C0026995|Myelogram (procedure) [Ambiguous]
C0026995|Myelogram [Ambiguous]
C0203103|Nephrotomography
C0203103|Tomography - kidneys (procedure)
C0203103|Tomography - kidneys
C0203103|Nephrotomogram
C0203103|Nephrotomogram (procedure)
C0203103|Tomography of kidney
C0203103|Nephrotomogram, NOS
C0203103|Nephrotomography, NOS
C0203103|Tomography of kidney, NOS
C0203108|Intravenous pyelogram
C0203108|intravenous pyelogram (procedure)
C0203108|X-ray renal intravenous pyelogram (IVP)
C0203108|Pyelogram;intravenous
C0203108|Intravenous pyelography
C0203108|Intravenous urogram (procedure)
C0203108|Retired procedure (procedure) [P5-60030]
C0203108|Intravenous urogram
C0203108|Retired procedure [P5-60030]
C0203108|IVP
C0203108|IVU
C0203108|Pyelogram intravenous
C0203108|Excretory urography
C0203108|Pyelogram
C0203108|Intravenous urography without KUB
C0203108|Intravenous pyelogram without KUB
C0203108|IVP - Intravenous pyelogram
C0203108|IVU - Intravenous urogram
C0203108|Intravenous urography
C0203108|Intravenous pyelogram, NOS
C0203108|Intravenous urography, NOS
C0008307|Cholangiographies
C0008307|Cholangiography
C0008307|Cholangiogram
C0008307|CHOLANGIOGR
C0008307|Biliary contrast radiography
C0008307|Biliary contrast radiography NOS
C0008307|Biliary contrast radiog
C0008307|Biliary contrast radiography NOS (procedure)
C0008307|Cholangiogram (procedure)
C0008307|Contrast radiography of bile ducts
C0008307|Biliary contrast radiography (procedure)
C0008307|Cholangiogram, NOS
C0008307|Contrast radiography of bile ducts, NOS
C1860232|X-RAY SENSITIVITY
C1860232|XRS
C2362745|(Radiology &/or physics in medicine) or (radiology) or (X-rays) (procedure)
C2362745|(Radiology &/or physics in medicine) or (radiology) or (X-rays)
C0412201|Chest wall sinogram
C0412201|Fistulogram of chest wall
C0412201|Fistulogram of chest wall (procedure)
C0412201|Sinogram of chest wall
C0412201|Chest wall fistulography
C0412201|Chest wall fistulography (procedure)
C0411329|Percutaneous imaging guided diagnostic aspiration
C0411329|Percutaneous imaging guided diagnostic aspiration (procedure)
C0203130|X-ray male external genitalia
C0203130|X-ray male external genitalia (procedure)
C0203130|Radiography of male genital organs (procedure)
C0203130|Radiography of male genital organs
C0203130|Radiography of male genital organs, NOS
C0554738|X-ray;leg
C0554738|Leg X-ray (procedure)
C0554738|Radiography of lower limb
C0554738|Lower limb X-ray
C0554738|Leg X-ray
C0554738|X-ray of lower limb
C0554738|Radiography of lower limb (procedure)
C0554738|X-ray NOS lower limb
C0554738|Radiography of lower limb, NOS
C0554738|X-ray of lower limb, NOS
C0554738|Leg X-ray procedure
C0554738|X-ray of the leg
C0203221|X-ray shoulder
C0203221|Radiography of shoulder
C0203221|x-ray of shoulder
C0203221|x-ray of shoulder (procedure)
C0203221|X-ray;shoulder
C0203221|Shoulder X-ray
C0203221|Shoulder X-ray (procedure)
C0203221|Glenoid X-ray
C0203221|Radiography of shoulder (procedure)
C0203221|Radiography of shoulder, NOS
C0203221|X-ray of the shoulder
C0411826|Stereotactic/stereoscopic test - mediastinum
C0411826|Stereotactic/stereoscopic test - mediastinum (procedure)
C0203768|Radioisotope scan of pancreas
C0203768|Radioisotope scan of pancreas (procedure)
C0200170|Ophthalmoscopy with medical evaluation, extended, with fluorescein angiography (procedure)
C0200170|Ophthalmoscopy with medical evaluation, extended, with fluorescein angiography
C0203054|X-ray gastrointestinal
C0203054|GI x-ray
C0203054|x-ray of gastrointestinal tract
C0203054|x-ray of gastrointestinal tract (procedure)
C0203054|X-ray;digestive tract
C0203054|Radiographic procedure on gastrointestinal tract
C0203054|Radiologic procedure on gastrointestinal tract
C0203054|Radiographic procedure on gastrointestinal tract (procedure)
C0203054|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Gastrointestinal Tract
C0203054|Gastrointestinal tract X-ray NOS
C0203054|Digestive tract X-ray
C0203054|GI tract X-ray NOS
C0203054|X-ray gastrointestinal tract
C0203054|X-ray NOS gastrointestinal tract
C0203054|Digestive tract X-ray NOS
C0203054|Radiography of gastrointestinal tract
C0203054|Gastrointestinal tract x-ray
C0203054|Radiography of gastrointestinal tract (procedure)
C0203054|Radiography of digestive tract, NOS
C0203054|Gastrointestinal tract x-ray, NOS
C0203054|X-ray of the digestive tract
C0203677|Transmission bone density study
C0203677|Transmission bone density study (procedure)
C0203677|Transmission bone imaging
C0203677|Transmission bone density study, NOS
C0203677|Transmission bone imaging, NOS
C0411827|Stereotactic/stereoscopic test - heart
C0411827|Stereotactic/stereoscopic test - heart (procedure)
C0411825|Stereotactic/stereoscopic test - lungs
C0411825|Stereotactic/stereoscopic test - lungs (procedure)
C0202677|Radiography of face, head AND/OR neck (procedure)
C0202677|Radiography of face, head AND/OR neck
C0202677|Radiography of face, head and neck, NOS
C0202757|Radiologic examination of neck
C0202757|Radiographic procedure on neck
C0202757|Diagnostic radiography of neck (procedure)
C0202757|Diagnostic radiography of neck
C0202757|Radiographic procedure on neck (procedure)
C1285408|Radiologic imaging, special views and positions (procedure)
C1285408|Radiologic imaging, special views and positions
C0202740|Radiography of uvula
C0202740|Radiography of uvula (procedure)
C0202740|Noncontrast x-ray of uvula
C0203015|Radiologic guidance for percutaneous drainage of abscess
C0203015|Radiologic guidance for percutaneous drainage of abscess (procedure)
C0202742|Radiography of nasolacrimal duct
C0202742|Radiography of nasolacrimal duct (procedure)
C0202742|Noncontrast x-ray of nasolacrimal duct
C0203236|X-ray radius and ulna
C0203236|x-ray of radius and ulna
C0203236|x-ray of radius and ulna (procedure)
C0203236|Radiography of forearm
C0203236|X-ray of forearm
C0203236|Radius and ulna X-ray
C0203236|Radius and ulna X-ray (procedure)
C0203236|Forearm X-ray
C0203236|Radiography of forearm (procedure)
C0203236|Radius and/or ulna X-ray (procedure)
C0203236|Radius and/or ulna X-ray
C0203236|Radius and ulna X-ray [Ambiguous]
C0203236|X-ray of the forearm
C0203236|X-ray of the radius/ulna
C0203236|X-ray;forearm
C0203236|X-ray;radius/ulna
C0203038|X-ray of gravid uterus
C0203038|Radiography of gravid uterus
C0203038|X-ray of gravid uterus (procedure)
C0203038|Radiography of gravid uterus (procedure)
C0203038|Radiography of gravid uterus (procedure) [Ambiguous]
C0202633|Radiologic supervision and interpretation of procedure (procedure)
C0202633|Radiologic supervision and interpretation of procedure
C0202633|Radiologic supervision and interpretation of procedure, NOS
C0412671|Digital slit-beam radiograph of leg length
C0412671|Digital slit-beam radiograph of leg length (procedure)
C0202811|Tracheography
C0202811|Tracheography (procedure)
C0202811|Tracheography, NOS
C0204135|Radiographic dental examination for personal identification
C0204135|Radiographic dental examination for personal identification (procedure)
C0203412|ultrasonic guidance for renal pelvis aspiration
C0203412|ultrasonic guidance for renal pelvis aspiration (procedure)
C0203036|Female genital organs X-ray
C0203036|X-ray NOS female genital organs
C0203036|X-ray of female genital organs
C0203036|Radiography of female genital organs (procedure)
C0203036|Radiography of female genital organs
C0203036|Radiography of female genital organs, NOS
C0203036|X-ray of female genital organs, NOS
C0202772|Radiography of adenoids
C0202772|Radiography of adenoids (procedure)
C0202772|Noncontrast x-ray of adenoid
C0203229|Diagnostic radiography of scapula
C0203229|x-ray of scapula (procedure)
C0203229|x-ray of scapula
C0203229|Scapula X-ray (procedure)
C0203229|Scapula X-ray
C0203229|Diagnostic radiography of scapula (procedure)
C0203229|Radiologic examination of scapula
C0203229|Diagnostic radiography of scapula, NOS
C0203229|Radiologic examination of scapula, NOS
C0411917|Diagnostic radiography of finger
C0411917|x-ray of finger (procedure)
C0411917|x-ray of finger
C0411917|Fingers X-ray (procedure)
C0411917|Fingers X-ray
C0411917|X-ray of fingers
C0411917|X-ray fingers
C0411917|Diagnostic radiography of finger (procedure)
C0411917|Diagnostic radiography of finger, NOS
C0411917|X-ray of fingers (procedure)
C0202849|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Heart
C0202849|Diagnostic radiography of heart
C0202849|Radiography of heart (procedure)
C0202849|Radiography of heart
C0202849|Radiography of heart, NOS
C0202849|Diagnostic radiography of heart, NOS
C0554740|pelvic x-ray (procedure)
C0554740|pelvic x-ray
C0554740|Pelvis X-ray
C0554740|X-ray;pelvis
C0554740|X-ray of pelvis
C0554740|Radiologic examination, pelvis
C0554740|Pelvis X-ray (procedure)
C0554740|X-ray of the pelvis
C0412753|Serial radiography of lungs (procedure)
C0412753|Serial radiography of lungs
C0034579|Orthopantomographies
C0034579|Panoramic Radiographies
C0034579|Pantomographies
C0034579|Radiographies, Panoramic
C0034579|Radiography, Panoramic
C0034579|ORTHOPANTOGRAM
C0034579|Panoramic Radiography
C0034579|PANORAMIC RADIOGR
C0034579|PANTOMOGR
C0034579|RADIOGR PANORAMIC
C0034579|ORTHOPANTOMOGR
C0034579|X-ray facial orthopantogram
C0034579|orthopantogram (procedure)
C0034579|X-ray teeth panoramic
C0034579|x-ray of teeth: panoramic (procedure)
C0034579|x-ray of teeth: panoramic
C0034579|Orthopantogram (eg, panoramic x-ray)
C0034579|Panoramic dental X-ray
C0034579|Pantomography dental
C0034579|Orthopantomography
C0034579|Pantomography
C0034579|Dental panoramic X-ray
C0034579|OPG - Orthopantomogram
C0034579|OPT - Orthopantomogram
C0034579|Orthopantograph
C0034579|Panoral X-ray
C0034579|PANORAMIC X-RAY OF JAWS
C0456846|Percutaneous computer tomography guided aspiration
C0456846|Percutaneous computer tomography guided aspiration (procedure)
C0203012|Radiologic guidance for percutaneous specimen collection
C0203012|Radiologic guidance for percutaneous specimen collection (procedure)
C0203215|Radiography of humerus
C0203215|x-ray of humerus (procedure)
C0203215|x-ray of humerus
C0203215|Humerus X-ray
C0203215|Humerus X-ray (procedure)
C0203215|Upper arm X-ray
C0203215|Radiography of humerus (procedure)
C0203215|Radiography of humerus, NOS
C0203215|X-ray of the humerus
C0203215|X-ray;humerus
C1299998|Plain film of head
C1299998|Plain film of head (procedure)
C0411832|Stereo-tactic/scopic investig.
C0411832|Stereotactic/stereoscopic investigation
C0411832|Stereotactic/stereoscopic investigation (procedure)
C0032743|Positron-Emission Tomography
C0032743|positron emission tomography
C0032743|PETT
C0032743|POSITRON EMISS TOMOGR
C0032743|TOMOGR POSITRON EMISS
C0032743|Positron emission tomographic imaging - action
C0032743|Positron emission tomographic imaging
C0032743|PET scan
C0032743|PET
C0032743|positron emission tomography (procedure)
C0032743|Positron emission tomogram
C0032743|Imaging, PET
C0032743|PET imaging
C0032743|PET Scans
C0032743|proton magnetic resonance spectroscopic imaging
C0032743|positron emission tomography scan
C0032743|Tomography, Positron-Emission
C0032743|PET - Positron emission tomography
C0032743|Positron emission tomographic imaging - action (qualifier value)
C0032743|Positron emission tomography, NOS
C0032743|PET scan, NOS
C0032743|Scan, PET
C0032743|Scans, PET
C0032743|Tomography, Positron Emission
C0032743|Medical Imaging, Positron Emission Tomography
C0032743|Positron emission tomography (PET)
C0202712|Radiography of supraorbital area
C0202712|Radiography of supraorbital area (procedure)
C0401265|Lithotripsy, extracorporeal shock wave
C0401265|ultrasonic fragmentation of urinary stones
C0401265|ultrasonic fragmentation of urinary stones (treatment)
C0401265|Ultrason fragment-stone
C0401265|LITHOTRIPSY XTRCORP SHOCK WAVE
C0401265|Extracorporeal shockwave lithotripsy for renal calculus NOS (procedure)
C0401265|Extracorporeal shockwave lithotripsy for renal calculus NOS
C0401265|Ultrasonic fragmentation of urinary stones (procedure)
C0401265|Extracorporeal shockwave lithotripsy of the kidney
C0401265|ESWL of kidney
C0401265|ESWL - Extracorporeal shockwave lithotripsy for renal calculus
C0401265|Extracorporeal fragmentation of renal calculus
C0401265|Extracorporeal shockwave lithotripsy for renal calculus
C0401265|Extracorporeal shockwave lithotripsy for renal calculus (procedure)
C0401265|Extracorporeal shockwave lithotripsy of the kidney (procedure)
C0401265|Ultrasonic fragmentation of urinary stone
C0401265|Ultrasonic fragmentation of urinary stone, NOS
C0401265|FRAGMENTING OF KIDNEY STONE
C0401265|Shattered urinary stones
C0456907|Plain X-ray guidance
C0456907|Plain X-ray guidance (procedure)
C0203139|Radiography of spine, NOS
C0203139|X-ray of spine, NOS
C0203139|Spinal x-ray, NOS
C0203139|Plain X-ray spine
C0203139|X-ray of spine
C0203139|Plain X-ray spine NOS
C0203139|Spine X-ray
C0203139|Vertebral column X-ray
C0203139|Back X-ray
C0203139|Vert. column X-ray
C0203139|X-ray of region of spine (procedure)
C0203139|X-ray of region of spine
C0203139|Plain X-ray spine NOS (procedure)
C0203139|X-ray NOS spine
C0203139|Spinal X-ray
C0203139|Radiography of spine
C0203139|Radiography of spine (procedure)
C0203139|Spinal x-ray NOS
C0203139|X-ray of the back
C0203139|X-ray of the spine
C0203139|X-ray;back
C0203139|X-ray;spine
C0203100|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Urinary Tract
C0203100|Radiographic procedure on genitourinary system (procedure)
C0203100|Radiographic procedure on genitourinary system
C0203100|Radiologic procedure on genitourinary system
C0519641|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Head and Neck
C1611783|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Vascular System
C0519643|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Upper Extremities
C0203138|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Spine and Pelvis
C0203138|Radiographic procedure on spine AND/OR pelvis (procedure)
C0203138|Radiographic procedure on spine AND/OR pelvis
C0203138|Radiologic procedure on spine AND/OR pelvis
C0412755|Other diagnostic radiology and related techniques
C0412755|Other diagnostic radiology NOS (procedure)
C0412755|Other diagnostic radiology NOS
C0412755|Other Diagnostic Radiology (Diagnostic Imaging) Related Procedures
C0519644|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Lower Extremities
C0519642|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Chest
C0519645|Diagnostic Radiology (Diagnostic Imaging) Procedures of the Abdomen
C0203025|Gynecological and Obstetrical Diagnostic Radiology (Diagnostic Imaging) Procedures
C0412112|Radiologic examination, small intestine, includes multiple serial films
C0412112|Small bowel series
C0412112|Radiologic examination, small intestine, includes multiple serial images
C0412112|RADEX SMALL INTESTINE W/MULTIPLE SERIAL IMAGES
C0412112|Radiography of digestive tract, small bowel series
C0412112|Diagnostic radiography of small bowel, serial films
C0412112|Radiologic examination of small bowel, serial films
C0412112|Small bowel series (procedure)
C0412112|X-RAY EXAM OF SMALL BOWEL
C0412112|Small intestine barium study
C0438647|Radiology/physics in medicine (procedure)
C0438647|Radiology/physics in medicine
C0438647|Physics in medicine
C0203184|Diagnostic radiography of sacrum
C0203184|x-ray of sacrum (procedure)
C0203184|x-ray of sacrum
C0203184|Sacral spine X-ray
C0203184|X-ray of sacral spine
C0203184|Sacrum X-ray
C0203184|Diagnostic radiography of sacrum (procedure)
C0203184|Diagnostic radiography of sacrum, NOS
C0203251|Diagnostic radiography of all fingers
C0203251|Diagnostic radiography of all fingers (procedure)
C0202763|x-ray of larynx
C0202763|x-ray of larynx (procedure)
C0202763|Diagnostic radiography of larynx
C0202763|Radiography of larynx
C0202763|Larynx X-ray
C0202763|Diagnostic radiography of larynx (procedure)
C0202763|Diagnostic roentgenographic imaging procedure on larynx
C0043348|Xeromammography
C0043348|XERORADIOGR BREAST
C0043348|BREAST XERORADIOGR
C0043348|XEROMAMMOGR
C0043348|Breast xerography
C0043348|Breast Xeroradiography
C0043348|Xeroradiography, Breast
C0043348|Xerography of breast
C0043348|Xeromammogram
C0043348|Xeromammography (procedure)
C0202575|Diagnostic radiography, oblique, special
C0202575|Diagnostic radiography, oblique, special (procedure)
C0202581|Diagnostic radiography, supine and erect studies
C0202581|Diagnostic radiography, supine and erect studies (procedure)
C0202587|Diagnostic radiography, special views
C0202587|Diagnostic radiography, special views (procedure)
C0202570|Diagnostic radiography, bilateral
C0202570|Diagnostic radiography, bilateral (procedure)
C0202578|Diagnostic radiography, combined posteroanterior and lateral (procedure)
C0202578|Diagnostic radiography, combined PA and lateral (procedure)
C0202578|Diagnostic radiography, combined posteroanterior and lateral
C0202578|Diagnostic radiography, combined PA and lateral
C0202592|Diagnostic radiography with oral contrast
C0202592|Diagnostic radiography with contrast media by ingestion
C0202592|Diagnostic radiography with oral contrast (procedure)
C0203102|X-ray of kidney, ureter & bladder
C0203102|KUB X-ray
C0203102|Radiography of kidney-ureter-bladder
C0203102|Kidneys, ureter, bladder X-ray
C0203102|Radiography of kidney-ureter-bladder (procedure)
C0203102|X-ray of the kidney/ureter/bladder
C0203102|X-ray;kidney/ureter/bladder
C0203064|Radiologic examination; esophagus
C0203064|x-ray of esophagus
C0203064|x-ray of esophagus (procedure)
C0203064|CONTRAST X-RAY ESOPHAGUS
C0203064|X-ray;oesophagus
C0203064|RADEX ESOPHAGUS
C0203064|Radiography of esophagus (procedure)
C0203064|Radiography of esophagus
C0203064|Radiography of oesophagus
C0203064|Radiologic examination of esophagus
C0203064|Radiologic examination of oesophagus
C0203064|Radiography of esophagus, NOS
C0203064|Radiologic examination of esophagus, NOS
C0203064|X-ray;esophagus
C0203064|X-ray of the esophagus
C0203064|X-ray of the oesophagus
C0203244|X-ray hand(s)
C0203244|Radiography of hand
C0203244|x-ray of hand
C0203244|x-ray of hand (procedure)
C0203244|X-ray;hand
C0203244|Hand X-ray (procedure)
C0203244|Hand X-ray
C0203244|Radiography of hand (procedure)
C0203244|Radiography of hand, NOS
C0203244|X-ray of the hand
C0203211|Upper limb X-ray
C0203211|X-ray NOS upper limb
C0203211|X-ray of upper limb
C0203211|Radiography of upper limb
C0203211|Radiography of upper limb (procedure)
C0203211|Radiography of upper limb, NOS
C0203211|X-ray of upper limb, NOS
C0203211|Radiographic procedure on upper extremity
C0411863|Radiography of mandible
C0411863|x-ray of mandible (procedure)
C0411863|x-ray of mandible
C0411863|Mandible X-ray (procedure)
C0411863|Mandible X-ray
C0411863|Lower jaw X-ray
C0411863|Radiography of mandible (procedure)
C0203170|Lumbar spine X-ray (procedure)
C0203170|Lumbar spine X-ray
C0203170|x-ray of lumbar spine
C0203170|x-ray of lumbar spine (procedure)
C0203170|x-ray lumbar spine
C0203170|Diagnostic radiography of lumbar spine
C0203170|Diagnostic radiography of lumbar spine (procedure)
C0203170|X-ray of the lumbar spine
C0203170|X-ray;spine;lumbar
C0203186|Diagnostic radiography of sacroiliac joints
C0203186|x-ray of sacroiliac joint
C0203186|x-ray of sacroiliac joint (procedure)
C0203186|X-ray of sacroiliac joints
C0203186|Sacroiliac joint X-ray
C0203186|Sacroiliac joint X-ray (procedure)
C0203186|Diagnostic radiography of sacroiliac joints (procedure)
C0411900|Clavicle X-ray
C0411900|x-ray of clavicle (procedure)
C0411900|x-ray of clavicle
C0411900|Clavicle X-ray (procedure)
C0411900|X-ray of the clavicle
C0411900|X-ray;clavicle
C0202722|Diagnostic radiography of temporomandibular joint
C0202722|Temporomandibular joint X-ray
C0202722|Temporomandibular joint X-ray (procedure)
C0202722|x-ray of temporomandibular joint (procedure)
C0202722|x-ray of temporomandibular joint
C0202722|x-ray temporomandibular joint
C0202722|TMJ X-ray
C0202722|Diagnostic radiography of temporomandibular joint (procedure)
C0202722|Diagnostic radiography of temporomandibular joint, NOS
C0202722|X-ray of the temporomandibular joint
C0202722|X-ray;temporomandibular joint
C0202746|Diagnostic radiography of orbits
C0202746|X-ray of orbits
C0202746|Orbits X-ray (procedure)
C0202746|Orbits X-ray
C0202746|x-ray of orbit
C0202746|x-ray face orbits
C0202746|x-ray of orbit (procedure)
C0202746|Diagnostic radiography of orbits (procedure)
C0202746|Radiography of orbit
C0202746|Diagnostic radiography of orbits, NOS
C0202746|Radiography of orbit, NOS
C0411950|Diagnostic radiography of coccyx
C0411950|Diagnostic radiography of coccyx (procedure)
C0203190|Diagnostic radiography of sacrococcygeal joint
C0203190|Diagnostic radiography of sacrococcygeal joint (procedure)
C0203188|Radiography of sacrococcygeal spine
C0203188|Diagnostic radiography of sacrum and coccyx
C0203188|Radiography of sacrococcygeal spine (procedure)
C0203066|Diagnostic radiography of cervical esophagus
C0203066|Diagnostic radiography of cervical oesophagus
C0203066|Diagnostic radiography of cervical esophagus (procedure)
C0412001|Diagnostic radiography of pharynx
C0412001|x-ray of pharynx
C0412001|x-ray of pharynx (procedure)
C0412001|Diagnostic roentgenographic imaging procedure on pharynx (procedure)
C0412001|Nasopharynx X-ray with water soluble contrast
C0412001|Pharynx X-ray
C0412001|Pharynx X-ray (procedure)
C0412001|Pharyngogram
C0412001|Diagnostic roentgenographic imaging procedure on pharynx
C0412001|Diagnostic radiography of pharynx (procedure)
C1963529|Neck X-ray
C1963529|x-ray of neck (procedure)
C1963529|x-ray of neck
C1963529|X-ray;neck
C1963529|X-ray of the neck
C0202732|X-ray face sinus
C0202732|Radiography of nasal sinuses
C0202732|X-ray;sinus
C0202732|X-ray of paranasal sinuses
C0202732|Plain X-ray facial sinuses (procedure)
C0202732|Plain X-ray facial sinuses
C0202732|x-ray of sinus (procedure)
C0202732|x-ray of sinus
C0202732|x-ray of paranasal sinus
C0202732|Diagnostic radiography of paranasal sinuses
C0202732|Sinuses X-ray
C0202732|Radiography of nasal sinuses (procedure)
C0202732|Radiography of nasal sinuses, NOS
C0202732|sinus X-ray
C0202727|Diagnostic radiography of mastoids
C0202727|Diagnostic radiography of mastoids (procedure)
C0085532|Angiographies, Coronary
C0085532|Coronary Angiographies
C0085532|Coronary Angiography
C0085532|Coronary arteriography
C0085532|ANGIOGR CORONARY
C0085532|CORONARY ANGIOGR
C0085532|coronary angiography (procedure)
C0085532|Arteriogram coronary
C0085532|Angiography;coronary
C0085532|Diagnostic Coronary Angiography
C0085532|Coronary angiogram
C0085532|Angiogram coronary
C0085532|Angiograph coronary
C0085532|Coronary angiograph
C0085532|Angiography, Coronary
C0085532|Coronary arteriogram
C0085532|Angiography of coronary arteries
C0085532|Coronary angiography, NOS
C0085532|Angiography of coronary arteries, NOS
C0085532|Coronary arteriography, NOS
C0085532|Coronary angiogram, NOS
C0085532|Coronary arteriography NOS
C0085532|Angiogram;coronary
C0017191|Gastrointestinal Transit
C0017191|Gastrointestinal Transits
C0017191|Transit, Gastrointestinal
C0017191|Transits, Gastrointestinal
C0017191|GI TRANSIT
C0017191|Gastrointestinal transit procedure
C0017191|Gastrointestinal transit study
C0017191|Gastrointestinal transit study (procedure)
C0008327|Cholecystographies
C0008327|Cholecystography
C0008327|CHOLECYSTOGR
C0008327|Cholecystogram
C0008327|CG - Cholecystogram
C0008327|Cholecystogram (procedure)
C0034185|pyelography
C0034185|PYELOGR
C0202590|Unilateral diagnostic radiographic imaging with contrast media
C0202590|Diagnostic radiography with contrast media, unilateral
C0202590|Diagnostic radiography with contrast media, unilateral (procedure)
C0202590|Unilateral diagnostic radiographic imaging with contrast media (situation)
C0202591|Diagnostic radiography with contrast media, bilateral
C0202591|Diagnostic radiography with contrast media, bilateral (procedure)
C0202593|Roentgenography, negative contrast (procedure)
C0202593|Roentgenography, negative contrast
C0202593|Roentgenography, negative contrast, NOS
C0202596|Diagnostic radiography with contrast media by injection, unilateral
C0202596|Unilateral diagnostic radiographic imaging with injection of contrast media (situation)
C0202596|Unilateral diagnostic radiographic imaging with injection of contrast media
C0202596|Diagnostic radiography with contrast media by injection, unilateral (procedure)
C0202597|Diagnostic radiography with contrast media by injection, bilateral
C0202597|Diagnostic radiography with contrast media by injection, bilateral (procedure)
C0202603|Diagnostic radiography double contrast (procedure)
C0202603|Diagnostic radiography double contrast
C0202603|Diagnostic radiography with contrast media by injection, positive and negative contrast (procedure)
C0202603|Diagnostic radiography with contrast media by injection, positive and negative contrast
C0202603|Diagnostic radiography double contrast, NOS
C0202603|Diagnostic radiography with contrast media by injection, positive and negative contrast, NOS
C0202603|Diagnostic radiography double contrast (procedure) [Ambiguous]
C0043304|SPECTROMETRY PROTON IND X RAY EMISS
C0043304|PROTON IND X RAY EMISS SPECTROMETRY
C0043304|Proton Induced X Ray Emission Spectrometry
C0043304|Spectrometry, Proton Induced X Ray Emission
C0043304|Proton-Induced X-Ray Emission Spectrometry
C0043304|Spectrometry, Proton-Induced X-Ray Emission
C0205954|Emission Spectroscopy, X-Ray
C0205954|Emission Spectroscopy, Xray
C0205954|Spectroscopy, X-Ray Emission
C0205954|Spectroscopy, Xray Emission
C0205954|X Ray Emission Spectroscopy
C0205954|X Ray Fluorescence Spectroscopy
C0205954|Fluorescence Spectroscopy, X-Ray
C0205954|Spectroscopy, X-Ray Fluorescence
C0205954|X-Ray Fluorescence Spectroscopies
C0205954|X-Ray Fluorescence Spectroscopy
C0205954|Xray Emission Spectroscopy
C0205954|X-Ray Emission Spectroscopy
C0206755|Crystallography, X-Ray
C0206755|Crystallographies, X Ray
C0206755|X Ray Crystallographies
C0206755|X ray crystallography
C0206755|CRYSTALLOGR XRAY
C0206755|XRAY CRYSTALLOGR
C0206755|X RAY CRYSTALLOGR
C0206755|CRYSTALLOGR X RAY
C0206755|X-ray crystallography
C0206755|Crystallography, Xray
C0206755|Crystallography, X Ray
C0206755|Xray Crystallography
C0206755|X-ray crystallography (procedure)
C0206755|Crystallography, X-Ray Diffraction
C0206755|Crystallography, X-Ray/Neutron
C0206755|Single Crystal Diffraction
C0024867|Mass Chest X Ray
C0024867|Mass Chest X-Ray
C0024867|Mass Chest X-Rays
C0024867|Mass Chest Xrays
C0024867|X-Ray, Mass Chest
C0024867|X-Rays, Mass Chest
C0024867|Xray, Mass Chest
C0024867|Xrays, Mass Chest
C0024867|Mass Chest Xray
C0411941|Calcaneum X-ray (procedure)
C0411941|Calcaneum X-ray
C0411941|Diagnostic radiography of calcaneus
C0411941|Heel X-Ray
C0411941|Os calcis X-ray
C0411941|Diagnostic radiography of calcaneus (procedure)
C0411941|X-ray of the heel
C0411941|X-ray;heel
C0202582|Diagnostic radiography, flexion and/or extension studies
C0202582|Diagnostic radiography, flexion and/or extension studies (procedure)
C0037804|Emission Spectrometry, X-Ray
C0037804|Emission Spectrometry, Xray
C0037804|Spectrometry, X Ray Emission
C0037804|Spectrometry, X-Ray Emission
C0037804|X Ray Emission Spectrometry
C0037804|Xray Emission Spectrometry
C0037804|PARTICLE IND X RAY EMISS SPECTROMETRY
C0037804|SPECTROMETRY PARTICLE IND X RAY EMISS
C0037804|X-ray fluorescence spectrometry
C0037804|X-ray fluorescence spectrometry (procedure)
C0037804|X-ray fluorescence spectromet. (procedure)
C0037804|X-ray fluorescence spectromet.
C0037804|Spectrometry, X-Ray Fluorescence
C0037804|Spectrometry, Xray Emission
C0037804|Particle Induced X Ray Emission Spectrometry
C0037804|X-Ray Emission Spectrometry
C0037804|Spectrometry, Particle-Induced X-Ray Emission
C0037804|Spectrometry, Particle Induced X Ray Emission
C0037804|Particle-Induced X-Ray Emission Spectrometry
C0037804|Fluorescence Spectrometry, X-Ray
C0037804|Spectrometry, X Ray Fluorescence
C0037804|X Ray Fluorescence Spectrometry
C0184695|Hospital admission, for laboratory work-up, radiography, etc.
C0184695|Hospital admission, for laboratory work-up, radiography, etc. (procedure)
C0200745|Electron microscopy study, scanning, examination and report
C0200745|Electron microscopy study, scanning, examination and report (procedure)
C0201818|Calculus analysis, quantitative, X-ray diffraction
C0201818|Calculus analysis, quantitative, X-ray diffraction (procedure)
C0202568|Diagnostic radiography, right
C0202568|Diagnostic radiography, right (procedure)
C0202569|Diagnostic radiography, left
C0202569|Diagnostic radiography, left (procedure)
C0202571|Diagnostic radiography, lateral
C0202571|Diagnostic radiography, lateral (procedure)
C0202572|Diagnostic radiography, anteroposterior (AP) (procedure)
C0202572|Diagnostic radiography, anteroposterior (procedure)
C0202572|Diagnostic radiography, anteroposterior
C0202572|Diagnostic radiography, anteroposterior (AP)
C0202573|Diagnostic radiography, posteroanterior (procedure)
C0202573|Diagnostic radiography, posteroanterior (PA) (procedure)
C0202573|Diagnostic radiography, posteroanterior
C0202573|Diagnostic radiography, posteroanterior (PA)
C0202574|Diagnostic radiography, oblique, standard
C0202574|Diagnostic radiography, oblique, standard (procedure)
C0202579|Diagnostic radiography, combined AP and lateral (procedure)
C0202579|Diagnostic radiography, combined anteroposterior and lateral
C0202579|Diagnostic radiography, combined anteroposterior and lateral (procedure)
C0202579|Diagnostic radiography, combined AP and lateral
C0202580|Diagnostic radiography, lateral decubitus studies
C0202580|Diagnostic radiography, lateral decubitus studies (procedure)
C0202583|Diagnostic radiography, minifilm
C0202583|Diagnostic radiography, minifilm (procedure)
C0008310|Cholangiopancreatographies, Endoscopic Retrograde
C0008310|Cholangiopancreatography, Endoscopic Retrograde
C0008310|Endoscopic Retrograde Cholangiopancreatographies
C0008310|Endoscopic Retrograde Cholangiopancreatography
C0008310|Retrograde Cholangiopancreatographies, Endoscopic
C0008310|Endoscopic retrograde choledochopancreatography
C0008310|CHOLANGIOPANCREATOGR ENDOSCOPIC RETROGRADE
C0008310|ENDOSCOPIC RETROGRADE CHOLANGIOPANCREATOGR
C0008310|RETROGRADE CHOLANGIOPANCREATOGR ENDOSCOPIC
C0008310|ERCP (endoscopic retrograde cholangiopancreatography)
C0008310|Endoscopic retrograde cholangiopancreatography -RETIRED-
C0008310|Endosc retro cholangiopa
C0008310|endoscopic retrograde cholangiopancreatography (procedure)
C0008310|endoscopic retrograde cholangiopancreatography (treatment)
C0008310|ERCP
C0008310|Diagnostic endoscopic retrograde examination of bile duct and pancreatic duct NOS
C0008310|Diagnostic endoscopic retrograde examination of bile duct and pancreatic duct
C0008310|ERCP - Endoscopic retrograde cholangiopancreatography
C0008310|Diagnostic endoscopic retrograde examination of bile duct and pancreatic duct NOS (procedure)
C0008310|Endoscopic retrograde cholangiopancreatography (ERCP)
C0008310|Retrograde Cholangiopancreatography, Endoscopic
C0008310|Endoscopic catheterization of pancreatic duct and bile duct systems
C0008310|Diagnostic endoscopic retrograde examination of bile duct and pancreatic duct (procedure)
C0008310|Endoscopic catheterisation of pancreatic duct and bile duct systems
C0008310|Endoscopic catheterization of pancreatic duct and bile duct systems (procedure)
C0008310|Endoscopic retrograde cholangiopancreatography, NOS
C0008310|ERCP, NOS
C0008310|Endoscopic retrograde cholangiopancreatography (procedure) [Ambiguous]
C0008310|Endoscopic retrograde cholangiopancreatography [ERCP]
C0203238|Skel xray-elbow/forearm
C0203238|Skeletal X-ray of elbow and forearm
C0203238|Skeletal X-ray of elbow and forearm (procedure)
C0203286|Skel xray-ankle & foot
C0203286|Skeletal X-ray of ankle and foot
C0203286|Skeletal X-ray of ankle and foot (procedure)
C0845973|X-ray study of eye
C0202777|Radiologic examination, teeth; complete, full mouth
C0202777|Full-mouth x-ray
C0202777|Full mouth x-ray of teeth (procedure)
C0202777|Full mouth x-ray of teeth
C0202777|RADIOLOGIC EXAM TEETH COMPLETE FULL MOUTH
C0202777|X-ray of teeth, full mouth
C0202777|Retired procedure [P5-11006]
C0202777|Retired procedure (procedure) [P5-11006]
C0202777|Full-mouth x-ray of teeth
C0002971|Angiocardiographies
C0002971|Angiocardiography
C0002971|ANGIOCARDIOGR
C0002971|Angiocardiography NOS
C0002971|Cardiac angiography
C0002971|Cardiac angiography (procedure)
C0002971|Cardioangiography
C0002971|Angiocardiography (procedure)
C0002971|Angiography of heart
C0002971|Angiocardiography, NOS
C0002971|Angiography of heart, NOS
C0002971|Angiocardiography, not otherwise specified
C0024219|Lymphangiographies
C0024219|Lymphangiogram
C0024219|LYMPHANGIOGR
C0024219|Lymphography
C0024219|lymphangiography
C0024219|lymphangiography (procedure)
C0024219|Lymphangiography NOS (procedure)
C0024219|Lymphatic system contrast procedure
C0024219|Lymphatic system contrast procedure (procedure)
C0024219|Contrast radiology of lymphatic tissue NOS
C0024219|Lymphangiography NOS
C0024219|Contrast radiology of lymphatic tissue NOS (procedure)
C0024219|Lymphatic system contrast procedure (disorder)
C0024219|Lymphangiograph
C0024219|Contrast radiology of lymphatic tissue
C0024219|Lymphogram
C0024219|Lymphangiogram (procedure)
C0024219|Lymphangiogram, NOS
C0024219|Lymphangiography, NOS
C0599271|heavy particle radiography
C0029562|Brain/skull contrst xray
C0029562|Other contrast radiogram of brain and skull
C0177719|Head tomography NEC
C0177719|Other tomography of head
C0177721|Contrast laryngogram
C0177722|Head soft tiss x-ray NEC
C0177722|Other soft tissue x-ray of face, head, and neck
C0029572|Dental x-ray NEC
C0029572|Other dental x-ray
C0177726|Facial bone x-ray NEC
C0177726|Other x-ray of facial bones
C0029875|Skull x-ray NEC
C0029875|Other x-ray of skull
C0177727|Cervical spine x-ray NEC
C0177727|Other x-ray of cervical spine
C0177728|Thoracic spine x-ray NEC
C0177728|Other x-ray of thoracic spine
C0177729|Lumbosac spine x-ray NEC
C0177729|Other x-ray of lumbosacral spine
C0177730|Spinal x-ray NEC
C0177730|Other x-ray of spine
C0029561|Contrast bronchogram NEC
C0029561|Other contrast bronchogram
C0177732|Contr mammary ductogram
C0177732|Contrast radiogram of mammary ducts
C0029664|Mammography NEC
C0029664|Other mammography
C0177733|Thorax sft tiss xray NEC
C0177733|Other soft tissue x-ray of chest wall
C0177735|Thoracic tomography NEC
C0177735|Other tomography of thorax
C0177737|Chest x-ray NEC
C0177737|Other chest x-ray
C0177737|Other x-ray of thorax
C0177739|Perc hepat Cholangiogram
C0177739|Percutaneous hepatic cholangiogram
C0029538|Cholangiogram NEC
C0029538|Other cholangiogram
C0177740|Biliary tract x-ray NEC
C0177740|Other biliary tract x-ray
C0177742|Intestinal x-ray NEC
C0177742|Other x-ray of intestine
C0009926|Contrast pancreatogram
C0177743|Digestive tract xray NEC
C0177743|Other digestive tract x-ray
C0177745|Nephrotomogram NEC
C0177745|Other nephrotomogram
C0177746|Percutaneous pyelogram
C0177747|Cystogram NEC
C0177747|Other cystogram
C0846489|Ileal conduitogram
C0846489|Fluoroscopic loopogram
C0846489|Fluoroscopic ileal conduitography (procedure)
C0846489|Fluoroscopic ileal conduitography
C0177749|Urinary system x-ray NEC
C0177749|Other x-ray of the urinary system
C0177750|Gas hysterosalpingogram
C0177750|Gas contrast hysterosalpingogram
C0177751|Dye hysterosalpingogram
C0177751|Opaque dye contrast hysterosalpingogram
C0177752|Tube & uterus x-ray NEC
C0177752|Other x-ray of fallopian tubes and uterus
C0177753|Female genital x-ray NEC
C0177753|Other x-ray of female genital organs
C0177756|Prostat/sem ves xray NEC
C0177756|Other x-ray of prostate and seminal vesicles
C0177757|Contrast epididymogram
C0177758|Contrast vasogram
C0177759|Epididymis/vas x-ray NEC
C0177759|Other x-ray of epididymis and vas deferens
C0177760|Male genital x-ray NEC
C0177760|Other x-ray of male genital organs
C0177762|Abdominal tomography NEC
C0177762|Other abdomen tomography
C0177763|Abdominal wall x-ray NEC
C0177763|Other soft tissue x-ray of abdominal wall
C0177764|Pelvic dye contrast xray
C0177764|Pelvic opaque dye contrast radiography
C0177766|Periton pneumogram NEC
C0177766|Other peritoneal pneumogram
C0177767|Retroperiton pneumogram
C0177767|Retroperitoneal pneumogram
C0177768|Retroperitoneal xray NEC
C0177768|Other retroperitoneal x-ray
C0029874|Abdominal x-ray NEC
C0029874|Other x-ray of abdomen
C0177770|Skl xray-shoulder/up arm
C0177770|Skeletal x-ray of shoulder and upper arm
C0177771|Skel xray-pelvis/hip NEC
C0177771|Other skeletal x-ray of pelvis and hip
C0177772|Skel xray-thigh/knee/leg
C0177772|Skeletal x-ray of thigh, knee, and lower leg
C0177774|Other skeletal x-ray
C0202999|Upper limb lymphangiogrm
C0202999|Arm lymphangiogram (procedure)
C0202999|Arm lymphangiogram
C0202999|Lymphangiography upper limb
C0202999|Lymphangiogram of upper extremity (procedure)
C0202999|Lymphangiogram of upper extremity
C0202999|Lymphangiogram of upper extremity, NOS
C0202999|Lymphangiogram of upper limb
C0177776|Up limb sft tis xray NEC
C0177776|Other soft tissue x-ray of upper limb
C0177778|Lo limb sft tis xray NEC
C0177778|Other soft tissue x-ray of lower limb
C0597417|roentgen videodensitometry
C0030796|Pelvimetries
C0030796|Pelvimetry
C0030796|Pelvimetry (procedure)
C0034592|Radioisotope Renographies
C0034592|Radioisotope Renography
C0034592|Renographies, Radioisotope
C0034592|Renography, Radioisotope
C0034592|radionuclide renography
C0034592|RADIOISOTOPE RENOGR
C0202686|Radiologic examination, sella turcica
C0202686|X-ray skull sella turcica
C0202686|Radiologic examination of sella turcica
C0202686|x-ray of sella turcica (procedure)
C0202686|x-ray of sella turcica
C0202686|X-RAY EXAM PITUITARY SADDLE
C0202686|RADIOLOGIC EXAMINATION SELLA TURCICA
C0202686|Diagnostic radiography of sella turcica
C0202686|Coned pituitary fossa X-ray
C0202686|Pituitary fossa X-ray
C0202686|Sella turcica X-ray
C0202686|Radiologic examination of sella turcica (procedure)
C0202725|Arthrogram of temporomandibular joint (procedure)
C0202725|Tm contrast arthrogram
C0202725|Temporomandibular joint arthrogram (procedure)
C0202725|Temporomandibular joint arthrogram
C0202725|Arthrogram of temporomandibular joint
C0202725|Temporomandibular contrast arthrogram
C0202735|Contrast radiography of nasal sinuses
C0202735|Contrast x-ray of sinus
C0202735|Contrast radiography of nasal sinuses (procedure)
C0202735|Contrast radiography of paranasal sinuses
C0202735|Contr.radiog.paranasal sinuses
C0202735|Contrast radiography of paranasal sinuses (procedure)
C0202735|Contrast radiogram of sinus
C0202745|Contrast dacryocystogram
C0202745|Contrast dacryocystogram (procedure)
C0202750|Contrast x-ray of orbit
C0202750|Contrast radiography orbit (procedure)
C0202750|Contrast radiography of orbit (procedure)
C0202750|Contrast radiography orbit
C0202750|Contrast radiography of orbit
C0202750|Contrast radiography of orbit, NOS
C0202750|Contrast radiogram of orbit
C0202806|Endotracheal bronchogram
C0202806|Endotracheal bronchography (procedure)
C0202806|Endotracheal bronchography
C0202806|Endotracheal bronchography, NOS
C0202806|Endotracheal bronchogram, NOS
C0202812|Mediastinal pneumogram
C0202812|Pneumomediastinography
C0202812|Mediastinal pneumogram (procedure)
C0202819|Radiologic examination of ribs, sternum and clavicle
C0202819|Rib/sternum/clavic x-ray
C0202819|X-ray of ribs, sternum and clavicle
C0202819|Radiologic examination of ribs, sternum AND clavicle (procedure)
C0202819|X-ray of ribs, sternum, and clavicle
C0202823|CT of chest (procedure)
C0202823|CT of thoracic region (procedure)
C0202823|Computed tomography of chest (procedure)
C0202823|Computed tomography of chest
C0202823|chest CT
C0202823|CAT scan of thorax
C0202823|CT of chest
C0202823|chest CT scan
C0202823|C.A.T. scan of thorax
C0202823|CT scan chest
C0202823|CT of thorax
C0202823|Retired procedure (procedure) [P5-20700]
C0202823|Retired procedure [P5-20700]
C0202823|Computerised tomogram thorax
C0202823|Computed tomography of thoracic region (procedure)
C0202823|CT of thoracic region
C0202823|Computed tomography of thoracic region
C0202823|Thorax CAT
C0202823|Computerized tomogram thorax
C0202823|Computerized axial tomography of thorax
C0202823|Tomography with use of computer, x-rays, and camera of thorax
C0202823|CT scan;chest
C0202823|CT scan of the chest
C0202842|Abdominal wall sinogram
C0202842|Fistulogram of abdominal wall
C0202842|Sinogram of abdominal wall
C0202842|Fistulogram of abdominal wall (procedure)
C0202843|Retroperiton fistulogram
C0202843|Retroperitoneal fistulogram
C0202843|Sinogram of retroperitoneum
C0202843|Retroperitoneal fistulogram (procedure)
C0202989|Cervical lymphangiogram
C0202989|Cervical lymphangiogram (procedure)
C0202990|Intrathor lymphangiogram
C0202990|Intrathoracic lymphangiogram (procedure)
C0202990|Thoracic lymphangiogram (procedure)
C0202990|Thoracic lymphangiogram
C0202990|Intrathoracic lymphangiogram
C0202990|Lymphangiography thorax
C0203040|percutaneous hysterogram
C0203040|percutaneous hysterogram (procedure)
C0203065|Barium swallow
C0203065|barium swallow (procedure)
C0203065|Barium swallow NOS
C0203065|Barium swallow NOS (procedure)
C0203065|an upper GI series - barium swallow
C0203065|BA - Barium swallow
C0203065|BS - Barium swallow
C0203065|Barium swallow (procedure) [Ambiguous]
C0203110|Retrograde pyelogram
C0203110|X-ray renal retrograde pyelogram
C0203110|retrograde pyelogram (procedure)
C0203110|Pyelogram retrograde
C0203110|Pyelogram;retrograde
C0203110|Retrograde urography
C0203110|RPG - Retrograde pyelogram
C0203110|Retrograde urogram
C0203110|Retrograde pyelography
C0203110|Retrograde ureteropyelography
C0203110|Retrograde pyelogram, NOS
C0203243|Skel xray-wrist & hand
C0203243|Skeletal X-ray of wrist and hand
C0203243|Skeletal X-ray of wrist and hand (procedure)
C0031545|Phlebographies
C0031545|Phlebography
C0031545|Venographies
C0031545|venography
C0031545|PHLEBOGR
C0031545|VENOGR
C0031545|venography (procedure)
C0031545|Venogram
C0031545|Venography - procedure
C0031545|Venography - procedure (procedure)
C0031545|Venograph
C0031545|Phlebogram
C0031545|Phlebography, NOS
C0031545|Phlebogram, NOS
C0031545|Venogram, NOS
C0031545|Venography, NOS
C0202991|Abdominal lymphangiogram
C0202991|Abdominal lymphangiogram (procedure)
C0202991|Lymphangiography abdomen
C0202991|Abdominal lymphangiogram, NOS
C0202741|Radiologic examination, salivary gland for calculus
C0202741|RADIOLOGIC EXAMINATION SALIVARY GLAND CALCULUS
C0202741|Retired procedure [P5-10375]
C0202741|Retired procedure (procedure) [P5-10375]
C0202741|X-RAY EXAM OF SALIVARY GLAND
C0202741|Noncontrast x-ray of salivary gland
C0864368|Intrauterine cephalometry by x-ray
C0202845|Pelvic gas contrast xray
C0202845|Gas contrast radiography of pelvis
C0202845|Pelvic pneumography
C0202845|Gas contrast radiography of pelvis (procedure)
C0202845|Pelvic gas contrast radiography
C0202845|Pelvic pneumoperitoneum
C0200746|Electron microscopy study, scanning, with X-ray analysis, examination and report
C0200746|Electron microscopy study, scanning, with X-ray analysis, examination and report (procedure)
C0553584|[V]Radiological examination NEC (context-dependent category)
C0553584|Encounter due to routine chest X-ray
C0553584|[V]Routine chest X-ray
C0553584|[V]Radiological examination NEC (situation)
C0553584|[V]Radiological examination NEC
C0553584|Routine chest x-ray
C0177755|Contr semin vesiculogram
C0177755|Contrast seminal vesiculogram
C0177779|Other C.A.T. scan
C0177779|Other CT scan
C0177779|CT scan - other
C0177779|Other computerized axial tomography
C0202784|Routine chest X-ray
C0202784|Standard chest X-ray NOS (procedure)
C0202784|Standard chest X-ray
C0202784|Standard chest X-ray NOS
C0202784|Standard chest X-ray (procedure)
C0202784|Routine chest X-ray (procedure)
C0202784|Chest X-ray - routine
C0202784|Routine chest x-ray, so described
C0412620|CT of abdomen (procedure)
C0412620|CT of abdominal organs (procedure)
C0412620|Computed tomography of abdomen (procedure)
C0412620|Computed tomography of abdomen
C0412620|CT of abdomen
C0412620|CT scan of abdomen
C0412620|abdominal CT scan
C0412620|C.A.T. scan of abdomen
C0412620|CT scan abdomen
C0412620|Computed tomography of abdominal organs (procedure)
C0412620|Computed tomography of abdominal organs
C0412620|CT of abdominal organs
C0412620|Computed tomography, abdomen
C0412620|CT scan - abdominal
C0412620|Computerized axial tomography of abdomen
C0412620|CT scan;abdomen
C0412620|CT scan of the abdomen
C0412623|abdominal CT kidney
C0412623|abdominal computed tomography kidney
C0412623|C.A.T. scan of kidney
C0412623|Kidney CT
C0412623|computed tomography of kidney
C0412623|CT scan of kidney
C0412623|CT scan of kidney (procedure)
C0412623|CT of kidney
C0412623|Computerized axial tomography of kidney
C0412623|CAT scan of kidney
C0412623|CT of kidneys
C0412623|Computerised axial tomography of kidney
C0412623|Computerized axial tomography of kidney (procedure)
C0412623|CT scan;kidney
C0412623|CT scan of the kidney
C0003844|Arteriographies
C0003844|ARTERIOGR
C0003844|arteriography
C0003844|Arteriography (procedure)
C0003844|Arteriography using contrast material
C0202748|Radiologic examination; optic foramina
C0202748|Diagnostic radiography of optic foramina
C0202748|X-ray of optic foramina
C0202748|x-ray of optic foramen
C0202748|x-ray of optic foramen (procedure)
C0202748|x-ray skull optic foramen
C0202748|Radiologic examination of optic foramina
C0202748|Optic foramina X-ray
C0202748|Diagnostic radiography of optic foramina (procedure)
C0202748|X-RAY EXAM OF EYE SOCKETS
C0202748|RADEX OPTIC FORAMINA
C0203082|intravenous cholangiography
C0203082|intravenous cholangiography (procedure)
C0203082|X-ray IV. cholangiography (IVC)
C0203082|Intraven cholangiogram
C0203082|Intravenous cholangiogram
C0203082|Intravenous cholangiogram (procedure)
C0203082|IVC - Intravenous cholangiogram
C0203082|Infusion cholangiogram
C0203145|C-spine x-ray
C0203145|x-ray of cervical spine
C0203145|x-ray of cervical spine (procedure)
C0203145|Radiography of cervical spine
C0203145|Cervical spine X-ray (procedure)
C0203145|Cervical spine X-ray
C0203145|Radiography of cervical spine (procedure)
C0203145|Radiography of cervical spine, NOS
C0203145|X-ray of cervical spine, NOS
C0203145|X-ray of the cervical spine
C0203145|X-ray;spine;cervical
C0203156|x-ray of thoracic spine (procedure)
C0203156|x-ray of thoracic spine
C0203156|T-spine x-ray
C0203156|Thoracic spine X-ray
C0203156|Thoracic spine X-ray (procedure)
C0203156|Radiography of thoracic spine
C0203156|Dorsal spine X-ray
C0203156|Radiography of thoracic spine (procedure)
C0203156|Radiography of thoracic spine, NOS
C0203156|X-ray of thoracic spine, NOS
C0203156|X-ray of the thoracic spine
C0203156|X-ray;spine;thoracic
C0203293|X-ray toes
C0203293|Diagnostic radiography of toes
C0203293|X-ray of toe
C0203293|X-ray of toes
C0203293|Toe X-ray (procedure)
C0203293|Toe X-ray
C0203293|x-ray of toes (procedure)
C0203293|Toes X-ray
C0203293|Diagnostic radiography of toes (procedure)
C0203293|Diagnostic radiography of toes, NOS
C0203293|X-ray;toe(s)
C0203293|X-ray of the toes
C0203075|Barium enema
C0203075|Barium Enema Injection
C0203075|lower GI series
C0203075|Lower GI series (procedure)
C0203075|Lower gastrointestinal series
C0203075|Lower gastrointestinal series (procedure)
C0203075|X-ray barium enema
C0203075|barium enema (procedure)
C0203075|Radiologic examination of colon with barium
C0203075|BA - Barium enema
C0203075|BE - Barium enema
C0203075|Lower gastrointestinal tract contrast procedure
C0203075|Lower gastrointestinal tract contrast procedure (procedure)
C0203075|Barium enema, NOS
C0203075|Barium enema (procedure) [Ambiguous]
C0203125|Retrogr cystourethrogram
C0203125|Retrograde urethrocystography
C0203125|Retrograde cystourethrogram
C0203125|Retrograde cystourethrogram (procedure)
C0203083|Intraoperative cholangiogram
C0203083|Intraoper cholangiogram
C0203083|Operative cholangiogram (procedure)
C0203083|Operative cholangiogram
C0203083|Cholangiography during surgery
C0203083|On table cholangiogram
C0203083|Peroperative cholangiogram
C0203083|Operative cholangiography
C0203083|Intraoperative cholangiogram (procedure)
C0202681|X-ray of skull
C0202681|X-ray skull
C0202681|x-ray of skull (procedure)
C0202681|X-ray;skull
C0202681|Plain X-ray skull NOS
C0202681|Plain X-ray skull
C0202681|Plain X-ray skull NOS (procedure)
C0202681|Skull X-ray
C0202681|X-ray NOS skull
C0202681|Diagnostic radiography of skull
C0202681|SXR - Skull X-ray
C0202681|Diagnostic radiography of skull (procedure)
C0202681|X-ray of the skull
C0599913|X ray visualization
C0202730|X-ray face nasal bones
C0202730|Diagnostic radiography of nasal bones
C0202730|X-ray of nasal bones
C0202730|X-ray (& plain)nose &/or malar
C0202730|X-ray (& plain)nose &/or malar (procedure)
C0202730|Nose X-ray
C0202730|Plain X-ray nasal/malar
C0202730|Nasal bone X-ray
C0202730|x-ray of nasal bones (procedure)
C0202730|X-ray of nose
C0202730|Radiography of nose
C0202730|Nasal bones X-ray
C0202730|Diagnostic radiography of nasal bones (procedure)
C0202730|X-ray of the nose
C0202730|X-ray;nose
C0202774|Nasophary contrast x-ray
C0202774|Contrast radiography of nasopharynx (procedure)
C0202774|Contrast radiography of nasopharynx
C0202774|Nasopharyngogram
C0202774|Contrast radiogram of nasopharynx
C0411916|Bone age studies
C0411916|X-RAYS FOR BONE AGE
C0411916|Radiography for bone age studies (procedure)
C0411916|bone age studies (procedure)
C0411916|Imaging for bone age assessment
C0411916|Radiography for bone age studies
C0411916|Bone age studies by X-ray
C0411916|Bone age X-ray
C0202709|x-ray of facial bones (procedure)
C0202709|x-ray of facial bones
C0202709|Diagnostic radiography of facial bones
C0202709|Facial bones X-ray
C0202709|Facial bones X-ray (procedure)
C0202709|x-ray of facial bone
C0202709|Diagnostic radiography of facial bones (procedure)
C0202709|Radiography of facial bones
C0202709|Radiography of facial bones, NOS
C0202709|X-ray of the facial bones
C0202709|X-ray;facial bone(s)
C0202830|Soft tissue X-ray chest wall
C0202830|Soft tissue X-ray chest wall (procedure)
C0202830|Soft tissue X-ray chest NOS
C0202830|Soft tissue X-ray chest NOS (procedure)
C0202830|Soft tissue X-ray chest
C0202830|Soft tissue X-ray chest (procedure)
C0202830|cxr thoracic wall soft tissue
C0202830|chest x-ray of thoracic wall soft tissue (procedure)
C0202830|chest x-ray of thoracic wall soft tissue
C0202830|Soft tissue X-ray of chest wall
C0202830|Soft tissue X-ray of chest wall (procedure)
C0202830|Soft tissue x-ray of thorax
C0202846|Radiography of retroperitoneum (procedure)
C0202846|Radiography of retroperitoneum
C0202846|Retroperitoneal X-ray
C0202846|Radiography of retroperitoneum, NOS
C0202846|Retroperitoneal X-ray, NOS
C0203002|Lower limb lymphangiogrm
C0203002|Leg lymphangiogram
C0203002|Leg lymphangiogram (procedure)
C0203002|Lymphangiography lower limb
C0203002|Lymphangiogram of lower extremity
C0203002|Lymphangiography of lower extremity (procedure)
C0203002|Lymphangiography of lower extremity
C0203002|Lymphangiography of lower extremity, NOS
C0203002|Lymphangiogram of lower extremity, NOS
C0203002|Lymphangiogram of lower limb
C0203101|X-ray;urinary tract
C0203101|X-ray NOS urinary system
C0203101|Urinary system X-ray NOS
C0203101|Urinary system X-ray
C0203101|Renal tract X-ray
C0203101|Urinary tract X-ray
C0203101|Radiography of urinary system (procedure)
C0203101|Radiography of urinary system
C0203101|Radiography of urinary system, NOS
C0203101|Urinary system x-ray, NOS
C0203101|X-ray of urinary system
C0203101|X-ray of the urinary tract
C0203192|Radiography of pelvic bones
C0203192|Radiography of pelvic bones (procedure)
C0581654|Skel xray-upper limb NOS
C0581654|Upper skeletal extremity X-ray
C0581654|Arm skeleton X-ray
C0581654|Skeletal X-ray of upper limb (procedure)
C0581654|Skeletal X-ray of upper limb
C0581654|Skeletal X-ray of upper limb, NOS
C0581654|Skeletal x-ray of upper limb, not otherwise specified
C0581655|Skel xray-lower limb NOS
C0581655|Lower skeletal extremity X-ray
C0581655|Leg skeleton X-ray
C0581655|Skeletal X-ray of lower limb (procedure)
C0581655|Skeletal X-ray of lower limb
C0581655|Skeletal X-ray of lower limb, NOS
C0581655|Skeletal x-ray of lower limb, not otherwise specified
C0186190|hip arthroscopy
C0186190|hip arthroscopy (treatment)
C0186190|arthroscopy of hip (procedure)
C0186190|arthroscopy of hip
C0186190|Arthroscopy, hip
C0186190|Diagnostic arthroscopy of hip joint
C0186190|Diagnostic arthroscopy of hip joint (procedure)
C0186190|Arthroscopy of hip, NOS
C0188624|ankle arthroscopy (treatment)
C0188624|ankle arthroscopy
C0188624|arthroscopy of ankle
C0188624|arthroscopy of ankle (procedure)
C0188624|Arthroscopy;ankle
C0188624|Arthroscopy, ankle
C0188624|Diagnostic arthroscopy of ankle joint
C0188624|Diagnostic arthroscopy of ankle joint (procedure)
C0188624|Arthroscopy of ankle, NOS
C0188624|arthroscopy of the ankle
C0864361|X-ray examination for fracture
C0202691|CT of structures of the head (procedure)
C0202691|head CT scan
C0202691|C.A.T. scan of head
C0202691|CT scan of head
C0202691|CT of head
C0202691|CT of head (procedure)
C0202691|Computed tomography of head (procedure)
C0202691|Head CT
C0202691|Computed tomography of structures of the head (procedure)
C0202691|Computed tomography of structures of the head
C0202691|CT of structures of the head
C0202691|Computed tomography of head
C0202691|CT scan of head (procedure)
C0202691|Computerized axial tomography of head
C0202691|CAT scan of head
C0202691|Computerized tomography of head
C0202691|Computerised axial tomography of head
C0202691|Computerised tomography of head
C0202691|CT scan;head
C0202691|CT scan of the head
C0203179|X-ray lumbosacral spine
C0203179|x-ray of lumbosacral spine
C0203179|LS spine x-ray
C0203179|x-ray of lumbosacral spine (procedure)
C0203179|Lumbosacral spine X-ray (procedure)
C0203179|Lumbosacral spine X-ray
C0203179|Radiography of lumbosacral spine
C0203179|X-ray of lumbosacral spine, NOS
C0203179|Radiography of lumbosacral spine, NOS
C0203179|X-ray of the lumbosacral spine
C0203179|X-ray;spine;lumbosacral
C0177738|Biliary tract X-ray
C0177738|Biliary tract X-ray (procedure)
C0177754|X-ray of male genital organs
C0177723|Other x-ray of face, head, and neck
C0177741|Other x-ray of digestive system
C1659593|Sialographies
C1659593|Sialography
C1659593|Sialogram
C1659593|SIALOGR
C1659593|Radiography of salivary gland
C1659593|X-ray sialography
C1659593|sialography (procedure)
C1659593|X-ray of salivary gland
C1659593|Radiography of salivary gland (procedure)
C1659593|Salivary gland X-ray (procedure)
C1659593|Contrast sialogram (procedure)
C1659593|Salivary gland X-ray
C1659593|Contrast sialogram
C1659593|Salivary glands--Radiography
C1659593|Dental saliography
C1659593|Radiography of salivary gland (procedure) [Ambiguous]
C1659593|salivary gland xray
C1659593|Xray;salivary gland
C2029656|head MRA without contrast followed by contrast
C2029656|magnetic resonance angiography of head without contrast followed by contrast
C2029656|magnetic resonance angiography of head without contrast followed by contrast (procedure)
C0918141|Magnetic resonance angiography, head; without contrast material(s)
C0918141|MRA HEAD W/O CONTRST MATERIAL
C0918141|MRA of head without contrast
C0918141|magnetic resonance angiography of head without contrast material
C0918141|MR angiography of the head without contrast material
C0918141|MR angiography of the head without contrast material (procedure)
C0918141|MR ANGIOGRAPHY HEAD W/O DYE
C0918143|Mr angiograph head w/o&w/dye
C0918143|Magnetic resonance angiography, head; without contrast material(s), followed by contrast material(s) and further sequences
C0918143|MRA HEAD W/O & W/CONTRAST MATERIAL
C0918143|MRA of head without contrast, followed by contrast and further sequences
C1997063|Plain X-ray guided wire localization of breast lesion (procedure)
C1997063|Plain X-ray guided wire localization of breast lesion
C1997063|X-ray guided wire localization of breast lesion
C1997063|Plain X-ray guided wire localisation of breast lesion
C1997063|X-ray guided wire localisation of breast lesion
C2315956|X-ray of thorax using mobile image intensifier (procedure)
C2315956|X-ray of thorax using mobile image intensifier
C2317240|X-ray of thoracic spine using mobile image intensifier (procedure)
C2317240|X-ray of thoracic spine using mobile image intensifier
C2584965|Mammogram in compression view (procedure)
C2584965|Mammogram in compression view
C2073430|X-ray chest bronchi
C2073430|x-ray of chest: bronchus (procedure)
C2073430|x-ray of chest: bronchus
C2073429|X-ray chest bronchioles
C2073429|x-ray of chest: bronchioles
C2073429|x-ray of chest: bronchioles (procedure)
C2073499|X-ray chest esophagus
C2073499|x-ray of chest: esophagus
C2073499|x-ray of chest: esophagus (procedure)
C2073658|X-ray chest pulmonary veins
C2073658|x-ray of chest: appearance of pulmonary veins (procedure)
C2073658|x-ray of chest: appearance of pulmonary veins
C2073515|X-ray chest hila
C2073515|x-ray of chest: appearance of hilum (procedure)
C2073515|x-ray of chest: appearance of hilum
C2073657|X-ray chest pulmonary vasculature
C2073657|x-ray of chest: pulmonary vasculature (procedure)
C2073657|x-ray of chest: pulmonary vasculature
C2073511|X-ray chest heart
C2073511|x-ray of chest: appearance of heart
C2073511|x-ray of chest: appearance of heart (procedure)
C2073488|X-ray chest diaphragm
C2073488|x-ray of chest: diaphragm (procedure)
C2073488|x-ray of chest: diaphragm
C2073582|X-ray chest mediastinum
C2073582|x-ray of chest: mediastinum
C2073582|x-ray of chest: mediastinum (procedure)
C2919783|X-ray of thoracic and lumbar spine (procedure)
C2919783|X-ray of thoracic and lumbar spine
C2919783|x-ray spine thoracic and lumbar
C2073600|X-ray chest pacemaker present
C2073600|x-ray of chest: pacemaker present
C2073600|x-ray of chest: pacemaker present (procedure)
C2073466|X-ray chest cardioverter-defibrillator present
C2073466|a chest x-ray showed a cardioverter-defibrillator present
C2073466|x-ray of chest: cardioverter-defibrillator present
C2073466|x-ray of chest: cardioverter-defibrillator present (procedure)
C2073710|review prior CXR film
C2073710|review previous chest x-ray
C2073710|review previous chest x-ray (procedure)
C2073713|x-ray of chest with computer analysis and physician review
C2073713|x-ray of chest with computer analysis and physician review (procedure)
C2318073|chest x-ray portable
C2318073|portable x-ray of chest (procedure)
C2318073|portable x-ray of chest
C2073592|X-ray chest no evidence of osteoarticular abnormalities seen
C2073592|no radiographic evidence of osteoarticular abnormalities is seen
C2073592|x-ray of chest: no evidence of osteoarticular abnormalities seen (procedure)
C2073592|x-ray of chest: no evidence of osteoarticular abnormalities seen
C2073709|x-ray of chest, views
C2073709|x-ray of chest, views (procedure)
C0581647|X-ray chest lungs
C0581647|X-ray of lungs (procedure)
C0581647|CXR lungs
C0581647|X-ray of lungs
C0581647|Lung X-ray
C0581647|Lung X-ray (procedure)
C0581647|X-ray of lung NOS
C2073601|X-ray chest pleura and thoracic wall
C2073601|x-ray of chest: pleura and thoracic wall
C2073601|x-ray of chest: pleura and thoracic wall (procedure)
C2073638|X-ray chest pulmonary arteries
C2073638|x-ray of chest: appearance of pulmonary arteries
C2073638|x-ray of chest: appearance of pulmonary arteries (procedure)
C3164095|Radiofrequency biopsy of breast using X-ray guidance
C3164095|Radiofrequency biopsy of breast using X-ray guidance (procedure)
C0202785|diagnostic chest x-ray, lateral view (procedure)
C0202785|cxr diagnostic lateral view
C0202785|diagnostic chest x-ray, lateral view
C0202785|Diagnostic radiography of chest, lateral
C0202785|Diagnostic radiography of chest, lateral (procedure)
C0202788|Diagnostic radiography of chest, posteroanterior
C0202788|Diagnostic radiography of chest, PA (procedure)
C0202788|Diagnostic radiography of chest, posteroanterior (procedure)
C0202788|cxr diagnostic pa view
C0202788|diagnostic chest x-ray, PA view
C0202788|diagnostic chest x-ray, PA view (procedure)
C0202788|Diagnostic radiography of chest, PA
C0202793|Diagnostic radiography of chest, combined PA and lateral (procedure)
C0202793|Diagnostic radiography of chest, combined posteroanterior and lateral (procedure)
C0202793|Diagnostic radiography of chest, combined posteroanterior and lateral
C0202793|diagnostic chest x-ray, PA and lateral views
C0202793|cxr diagnostic pa and lateral views
C0202793|diagnostic chest x-ray, PA and lateral views (procedure)
C0202793|Diagnostic radiography of chest, combined PA and lateral
C0202786|diagnostic chest x-ray, stereo
C0202786|cxr diagnostic stereo
C0202786|diagnostic chest x-ray, stereo (procedure)
C0202786|Diagnostic radiography of chest, stereo
C0202786|Diagnostic radiography of chest, stereo (procedure)
C0202790|Diagnostic radiography of chest, oblique, standard
C0202790|Diagnostic radiography of chest, oblique, standard (procedure)
C0202789|cxr diagnostic minifilm
C0202789|diagnostic chest x-ray, minifilm (procedure)
C0202789|diagnostic chest x-ray, minifilm
C0202789|Diagnostic radiography of chest, minifilm
C0202789|Diagnostic radiography of chest, minifilm (procedure)
C0420046|Screening chest X-ray (procedure)
C0420046|Screening chest X-ray
C0420046|CXR - screening
C1964255|chest x-ray of thoracic wall (procedure)
C1964255|chest x-ray of thoracic wall
C1964255|cxr thoracic wall
C1964255|Radiography of chest wall (procedure)
C1964255|X-ray of chest wall
C1964255|Radiography of chest wall
C1964255|Radiography of chest wall, NOS
C1964255|X-ray of chest wall, NOS
C0202787|Radiologic examination, chest; stereo, frontal
C0202787|chest X-ray stereo, frontal
C0202787|RADIOLOGIC EXAMINATION CHEST STERO FRONTAL
C0202787|CHEST X-RAY STEREO FRONTAL
C0202787|X-ray of chest, stereo, front
C0202787|Retired procedure (procedure) [P5-20032]
C0202787|Retired procedure [P5-20032]
C0202787|CXR with stereo frontal views (procedure)
C0202787|CXR with stereo frontal views
C0202821|Radiologic examination; sternum, minimum of two views
C0202821|Radiologic examination; sternum, minimum of 2 views
C0202821|X-RAY EXAM BREASTBONE 2/>VWS
C0202821|Retired procedure [P5-20672]
C0202821|Retired procedure (procedure) [P5-20672]
C0202821|X-ray of sternum, minimum of 2 views
C0202821|RADEX STERNUM MINIMUM 2 VIEWS
C0202791|Radiologic examination, chest; single view, frontal
C0202791|RADIOLOGIC EXAMINATION CHEST SINGLE VIEW FRONTAL
C0202791|CHEST X-RAY 1 VIEW FRONTAL
C0202791|X-ray of chest, 1 view, front
C0202791|Retired procedure [P5-20070]
C0202791|Retired procedure (procedure) [P5-20070]
C0202822|Radiologic examination; sternoclavicular joint or joints, minimum of three views
C0202822|Radiologic examination; sternoclavicular joint or joints, minimum of 3 views
C0202822|RADEX STERNOCLAVICULAR JT/JTS MINIMUM 3 VIEWS
C0202822|X-RAY STRENOCLAVIC JT 3/>VWS
C0202822|Retired procedure [P5-20674]
C0202822|Retired procedure (procedure) [P5-20674]
C0202822|X-ray of sternoclavicular joint, minimum of 3 views
C0202799|Radiologic examination, chest, special views (eg, lateral decubitus, Bucky studies)
C0202799|RADEX CHEST SPECIAL VIEWS
C0202799|CHEST X-RAY SPECIAL VIEWS
C0202799|Retired procedure [P5-20160]
C0202799|Retired procedure (procedure) [P5-20160]
C0202795|Radiologic examination, chest, two views, frontal and lateral; with oblique projections
C0202795|Radiologic examination, chest, 2 views, frontal and lateral; with oblique projections
C0202795|CHEST X-RAY FRNT LAT OBLIQUE
C0202795|RADEX CH 2 VIEWS FRONTAL & LATERAL OBLIQUE PRJCJ
C0202795|Retired procedure [P5-20120]
C0202795|Retired procedure (procedure) [P5-20120]
C0202794|Radiologic examination, chest, two views, frontal and lateral; with apical lordotic procedure
C0202794|Radiologic examination, chest, 2 views, frontal and lateral; with apical lordotic procedure
C0202794|RADEX CH 2 VIEWS FRNT & LAT APICAL LORDOTIC PX
C0202794|CHEST X-RAY FRNT LAT LORDOTC
C0202794|Retired procedure [P5-20110]
C0202794|Retired procedure (procedure) [P5-20110]
C0202792|Radiologic examination, chest, two views, frontal and lateral
C0202792|Radiologic examination, chest, 2 views, frontal and lateral
C0202792|RADIOLOGIC EXAM CHEST 2 VIEWS FRONTAL&LATERAL
C0202792|CHEST X-RAY 2VW FRONTAL&LATL
C0202792|Retired procedure [P5-20080]
C0202792|Retired procedure (procedure) [P5-20080]
C3838010|cxr bowel present in chest (procedure)
C3838010|cxr bowel present in chest
C3838009|chest x-ray for chest diameter measurement (procedure)
C3838009|chest x-ray for chest diameter measurement
C3838009|cxr diameter
C3838008|cxr liver present in chest
C3838008|cxr liver present in chest (procedure)
C3863804|CXR on expiration (procedure)
C3863804|CXR on expiration
C3863771|CXR with nipple markers
C3863771|CXR with nipple markers (procedure)
C3863812|cxr four or more views
C3863812|CXR, four or more views (procedure)
C3863812|CXR, four or more views
C3863775|cxr two views (procedure)
C3863775|cxr two views
C3863810|CXR, four views
C3863810|cxr four views
C3863810|CXR, four views (procedure)
C3863773|CXR, two views, with nipple markers
C3863773|CXR, two views, with nipple markers (procedure)
C3863773|cxr two views with nipple markers
C3863779|cxr single view
C3863779|CXR, single view
C3863779|CXR, single view (procedure)
C3863777|cxr two or more views
C3863777|CXR, two or more views
C3863777|CXR, two or more views (procedure)
C3863803|CXR on inspiration
C3863803|CXR on inspiration (procedure)
C3863809|cxr left lateral upright view
C3863809|CXR, left lateral upright view
C3863809|CXR, left lateral upright view (procedure)
C3863815|CXR, AP left lateral decubitus view (procedure)
C3863815|CXR, AP left lateral decubitus view
C3863815|cxr ap left lateral decubitus view
C3863770|CXR with oral contrast
C3863770|CXR with oral contrast (procedure)
C3863820|CXR with AP right lateral decubitus views
C3863820|CXR with AP right lateral decubitus views (procedure)
C3863820|cxr anteroposterior and right lateral decubitus views
C3863813|CXR during surgery (procedure)
C3863813|CXR during surgery
C3863774|cxr two views with apical view
C3863774|CXR, two views with apical view
C3863774|CXR, two views with apical view (procedure)
C3863817|CXR, AP and AP right lateral decubitus views (procedure)
C3863817|CXR, AP and AP right lateral decubitus views
C3863817|cxr ap and ap right lateral decubitus views
C3863818|CXR with AP, lateral, and right and left oblique views
C3863818|cxr anteroposterior, lateral, right and left oblique views
C3863818|CXR with AP, lateral, and right and left oblique views (procedure)
C3863778|CXR, three views
C3863778|cxr three views
C3863778|CXR, three views (procedure)
C3863802|CXR on inspiration and expiration
C3863802|CXR on inspiration and expiration (procedure)
C3863816|CXR, AP and PA upright views (procedure)
C3863816|CXR, AP and PA upright views
C3863816|cxr ap and pa upright views
C3863814|CXR with AP right and left lateral decubitus views (procedure)
C3863814|cxr, ap right and left lateral decubitus views
C3863814|CXR with AP right and left lateral decubitus views
C1629851|X-ray of chest and abdomen
C1629851|x-ray chest and abdomen
C1629851|chest and abdomen x-ray (procedure)
C1629851|chest and abdomen x-ray
C1629851|X-ray of chest and abdomen (procedure)
C4029408|cxr diagnostic
C4029408|diagnostic chest x-ray (procedure)
C4029408|diagnostic chest x-ray
C0202813|Radiography of ribs
C0202813|X-ray;ribs
C0202813|Ribs X-ray (procedure)
C0202813|Ribs X-ray
C0202813|X-ray of ribs
C0202813|X-ray of ribs (procedure)
C0202813|X-ray of rib
C0202813|X-ray of rib (procedure)
C0202813|Radiography of ribs (procedure)
C0202813|Radiography of ribs, NOS
C0202813|X-ray of the ribs
C4075943|X-ray guided localization of iodine 125 radioactive seed to breast lesion
C4075943|Localisation of iodine 125 radioactive seed to breast lesion using X-ray guidance
C4075943|Localization of iodine 125 radioactive seed to breast lesion using X-ray guidance
C4075943|X-ray guided localisation of iodine 125 radioactive seed to breast lesion
C4075943|Localization of iodine 125 radioactive seed to breast lesion using X-ray guidance (procedure)
C0203292|Radiologic examination; calcaneus, minimum of 2 views
C0203292|Retired procedure (procedure) [P5-90208]
C0203292|Retired procedure [P5-90208]
C0203292|X-ray of calcaneus, minimum of 2 views
C0203292|X-RAY EXAM OF HEEL
C0203292|RADEX CALCANEUS MINIMUM 2 VIEWS
C0203270|Radiologic examination; lower extremity, infant, minimum of 2 views
C0203270|X-RAY EXAM OF LEG INFANT
C0203270|RADEX LOWER EXTREMITY INFANT MINIMUM 2 VIEWS
C0203270|Retired procedure (procedure) [P5-90122]
C0203270|Retired procedure [P5-90122]
C0203270|X-ray of lower extremity of infant, minimum of 2 views
C0203294|Radiologic examination; toe(s), minimum of 2 views
C0203294|X-ray of toes, minimum of 2 views
C0203294|Retired procedure [P5-90222]
C0203294|Retired procedure (procedure) [P5-90222]
C0203294|X-ray of toe, minimum of 2 views
C0203294|X-RAY EXAM OF TOE(S)
C0203294|RADEX TOE MINIMUM 2 VIEWS
C0203278|Radiologic examination; tibia and fibula, 2 views
C0203278|RADIOLOGIC EXAMINATION TIBIA & FIBULA 2 VIEWS
C0203278|X-ray of tibia and fibula, 2 views
C0203278|X-RAY EXAM OF LOWER LEG
C0202769|Radiologic examination; pharynx or larynx, including fluoroscopy and/or magnification technique
C0202769|Retired procedure (procedure) [P5-10640]
C0202769|Retired procedure [P5-10640]
C0202769|THROAT X-RAY & FLUOROSCOPY
C0202769|RADEX PHARYNX/LARX W/FLUOR&/MAGNIFICATION TQ
C0202747|Radiologic examination; orbits, complete, minimum of four views
C0202747|Radiologic examination; orbits, complete, minimum of 4 views
C0202747|RADEX ORBITS COMPLETE MINIMUM 4 VIEWS
C0202747|Retired procedure (procedure) [P5-10410]
C0202747|Retired procedure [P5-10410]
C0202747|X-RAY EXAM OF EYE SOCKETS
C0373198|Radiologic examination; pharynx and/or cervical esophagus
C0373198|RADEX PHARYNX&/CERVICAL ESOPHAGUS
C0373198|CONTRST X-RAY EXAM OF THROAT
C0203217|Radiologic examination; upper extremity, infant, minimum of 2 views
C0203217|X-RAY EXAM OF ARM INFANT
C0203217|RADEX UPPER EXTREMITY INFANT MINIMUM 2 VIEWS
C0203217|X-ray of arm in infant minimum of 2 views
C0203217|Retired procedure [P5-80036]
C0203217|Retired procedure (procedure) [P5-80036]
C0203217|X-ray of upper extremity of infant, minimum of 2 views
C0373176|Radiologic examination; scapula, complete
C0373176|RADEX SCAPULA COMPLETE
C0373176|X-RAY EXAM OF SHOULDER BLADE
C0373179|Radiologic examination; acromioclavicular joints, bilateral, with or without weighted distraction
C0373179|RADEX A-C JOINTS BI W/WO WEIGHTED DISTRCJ
C0373179|X-RAY EXAM OF SHOULDERS
C0203226|Radiologic examination; clavicle, complete
C0203226|RADEX CLAVICLE COMPLETE
C0203226|Radiologic examination of clavicle, complete
C0203226|Radiography of clavicle, complete
C0203226|Radiologic examination of clavicle, complete (procedure)
C0203226|X-RAY EXAM OF COLLAR BONE
C0203216|Radiologic examination; humerus, minimum of 2 views
C0203216|RADEX HUMERUS MINIMUM 2 VIEWS
C0203216|Retired procedure (procedure) [P5-80034]
C0203216|Retired procedure [P5-80034]
C0203216|X-ray of humerus, minimum of 2 views
C0203216|X-RAY EXAM OF HUMERUS
C3515830|Radiologic examination; forearm, 2 views
C3515830|RADEX FOREARM 2 VIEWS
C3515830|X-ray of forearm, 2 views
C3515830|X-RAY EXAM OF FOREARM
C2729424|Pet tumor init tx strat
C2729424|Positron emission tomography (pet) or pet/computed tomography (ct) to inform the initial treatment strategy of tumors that are biopsy proven or strongly suspected of being cancerous based on other diagnostic testing
C0412534|ultrasound abdominal liver
C0412534|abdominal ultrasound liver
C0412534|Ultrasound liver
C0412534|hepatic ultrasound
C0412534|liver ultrasound
C0412534|ultrasound of abdomen: appearance of liver (procedure)
C0412534|ultrasound of abdomen: appearance of liver
C0412534|US scan of liver
C0412534|US scan of liver (procedure)
C0412534|LUSS - Ultrasound scan of liver
C0412534|Ultrasonography of liver
C0412534|Liver US scan
C0412534|Ultrasonography of liver (procedure)
C0412534|ultrasound of the liver
C0412534|Ultrasound;liver
C0411889|Liver soft tissue X-ray
C0411889|Liver soft tissue X-ray (procedure)
C0412760|Thermography - hepatic region (procedure)
C0412760|Thermography - hepatic region
C0412694|MRI of liver (procedure)
C0412694|Magnetic resonance imaging of liver (procedure)
C0412694|Magnetic Resonance Imaging (MRI) of Liver
C0412694|MRI of liver
C0412694|Magnetic resonance imaging of liver
C0203765|Liver and spleen imaging
C0203765|Imaging of liver and spleen
C0203765|Liver and spleen imaging (procedure)
C0203758|liver scanning
C0203758|Radioisotope function study of liver
C0203758|Liver scan/isotope funct
C0203758|liver imaging
C0203758|Radioisotope function study of liver (procedure)
C0203758|Radionuclide hepatic function study
C0203758|Liver scan
C0203758|Radionuclide liver studies
C0203758|Liver isotope studies
C0203758|Liver scan NOS
C0203758|Scan liver NOS
C0203758|Radioisotope study of liver (procedure)
C0203758|Radioisotope study of liver
C0203758|Liver scan and radioisotope function study
C2316126|Single photon emission computed tomography (SPECT) of hemangioma of liver
C2316126|Single photon emission computed tomography of hemangioma of liver
C2316126|Single photon emission computed tomography of haemangioma of liver
C2316126|Single photon emission computed tomography of hemangioma of liver (procedure)
C2316126|Single photon emission computed tomography (SPECT) of haemangioma of liver
C0203761|Liver imaging; with vascular flow
C0203761|LIVER IMAGING W/VASCULAR FLOW
C0203761|Imaging of liver blood flow
C0203761|Liver imaging with vascular flow
C0203761|Liver imaging with vascular flow (procedure)
C0203761|LIVER IMAGING WITH FLOW
C0202977|venography of liver (procedure)
C0202977|venography of liver
C0202977|Hepatic venography
C0202977|Hepatic venogram
C0202977|Hepatic venography (procedure)
C0202977|Hepatic phlebography
C0203759|Liver imaging; static only
C0203759|Isotope static scan liver
C0203759|LIVER IMAGING STATIC ONLY
C0203759|Isotope static scan liver (procedure)
C0203759|Retired procedure (procedure) [P5-D5051]
C0203759|Retired procedure [P5-D5051]
C0203759|Liver imaging
C4039140|Liver angiography
C4039140|Angiography of liver (procedure)
C4039140|Angiography of liver
C4039879|Imaging guided percutaneous fine needle aspiration biopsy of liver
C4039879|Percutaneous fine needle aspiration biopsy of liver using imaging guidance (procedure)
C4039879|Percutaneous fine needle aspiration biopsy of liver using imaging guidance
C2315171|Single photon emission computed tomography of liver and spleen
C2315171|Single photon emission computed tomography of liver and spleen (procedure)
C2315171|Single photon emission computed tomography (SPECT) of liver and spleen
C2317182|Magnetic resonance imaging (MRI) of liver and spleen
C2317182|Magnetic resonance imaging of liver and spleen (procedure)
C2317182|Magnetic resonance imaging of liver and spleen
C2317182|MRI of liver and spleen
C0473930|Tc99m-labeled colloid liver and spleen study - dynamic (procedure)
C0473930|Tc99m-labelled colloid liver and spleen study - dynamic (procedure)
C0473930|Tc99m-labeled colloid liver and spleen study - dynamic
C0473930|Tc99m-labelled colloid liver and spleen study - dynamic
C0412394|Radionuclide study of liver, spleen and biliary tract
C0412394|Radionuclide study of liver, spleen and biliary tract (procedure)
C0203767|Liver and spleen imaging; with vascular flow
C0203767|LIVER & SPLEEN IMAGING W/VASCULAR FLOW
C0203767|Liver and spleen imaging with vascular flow
C0203767|Liver and spleen imaging with vascular flow (procedure)
C0203767|LIVER & SPLEEN IMAGE/FLOW
C0473931|Tc99m-labeled colloid liver and spleen study - static (procedure)
C0473931|Tc99m-labelled colloid liver and spleen study - static
C0473931|Tc99m-labelled colloid liver and spleen study - static (procedure)
C0473931|Tc99m-labeled colloid liver and spleen study - static
C0203766|Liver and spleen imaging; static only
C0203766|LIVER & SPLEEN IMAGING STATIC ONLY
C0203766|Retired procedure [P5-D5064]
C0203766|Retired procedure (procedure) [P5-D5064]
C0203766|Liver and spleen imaging
C1644183|Radionuclide liver and spleen imaging procedure (procedure)
C1644183|Radionuclide liver and spleen imaging procedure
C1644183|Radionuclide liver and spleen study
C0476419|[D]Abnormal liver scan (context-dependent category)
C0476419|[D]Abnormal liver scan (situation)
C0476419|[D]Abnormal liver scan
C0476419|Scan liver NOS abnormal
C0476419|Liver scan abnormal
C0476419|Liver scan NOS abnormal
C0476419|Abnormal liver scan
C3648818|imaging studies nonspecific abnormal findings liver
C3648818|imaging studies: nonspecific abnormal findings of liver
C3648818|nonspecific abnormal imaging findings of liver
C3648818|imaging studies: nonspecific abnormal findings of liver (procedure)
C4076645|Ultrasonography of liver abnormal (finding)
C4076645|Ultrasonography of liver abnormal
C2227710|abdominal x-ray, AP view: biliary calcification
C2227710|abdominal x-ray, AP view: biliary calcification (procedure)
C0495790|Abnormal findings on diagnostic imaging of liver and biliary tract
C0495790|Abnormal findings on dx imaging of liver and biliary tract
C0495790|Abnormal findings diagnostic imaging of liver and biliary tract
C0495790|Abnormal findings diagnostic imaging of liver+biliary tract
C0495790|Abnormal findings diagnostic imaging of liver+biliary tract (finding)
C0495790|Abnormal findings diagnostic imaging of liver and biliary tract (finding)
C1385723|diagnostic imaging; abnormal, bile ducts (common) (hepatic)
C1385723|abnormal; diagnostic imaging, bile ducts (common) (hepatic)
C1385728|diagnostic imaging; abnormal, liver
C1385728|abnormal; diagnostic imaging, liver
C0347946|[D]Gallbladder nonvisualization (context-dependent category)
C0347946|Nonvisualization of gallbladder
C0347946|[D]Gallbladder nonvisualisation
C0347946|[D]Gallbladder nonvisualization (situation)
C0347946|[D]Gallbladder nonvisualization
C0347946|Nonvisualisation of gallbladder
C0347946|Nonvisualization of gallbladder (finding)
C0347946|nonvisualization; gallbladder
C2047961|imaging studies: nonspecific abnormal finding of biliary tract (procedure)
C2047961|imaging studies: nonspecific abnormal finding of biliary tract
C2585276|Radionuclide study of perfusion of liver
C2585276|Radionuclide study of perfusion of liver (procedure)
C2108323|radioisotope scan of liver (procedure)
C2108323|radioisotope scan of liver
C2054285|technetium scan of liver (procedure)
C2054285|technetium scan of liver
C0412396|Isotope dynamic liver scan (procedure)
C0412396|Isotope dynamic liver scan
C0203760|Liver function study with serial images
C0203760|Liver function study with serial images (procedure)
C0589338|Dynamic non-imaging isotope: liver (& [study]) (procedure)
C0589338|Dynamic non-imaging isotope: liver (& [study])
C0589338|Dynamic non-imaging isotope study: liver (procedure)
C0589338|Dynamic non-imaging isotope study: liver
C0589338|Dynam.non-im.isotope: liver
C0581583|Tc99m-labelled colloid liver study - dynamic
C0581583|Tc99m-labeled colloid liver study - dynamic
C0581583|Tc99m-labeled colloid liver study - dynamic (procedure)
C0581583|Tc99m-labelled colloid liver study - dynamic (procedure)
C0581584|Tc99m-labeled colloid liver study - static
C0581584|Tc99m-labelled colloid liver study - static
C0581584|Tc99m-labelled colloid liver study - static (procedure)
C0581584|Tc99m-labeled colloid liver study - static (procedure)
C0203764|Radiolabeled Rose Bengal study
C0203764|Radioiodinated rose bengal study of liver
C0203764|Radiolabelled Rose Bengal study
C0203764|Radioiodinated rose bengal study of liver (procedure)
C0679575|neuroimaging
C0600032|Diagnostic imaging NOS
C0600032|Diagnostic imaging, not elsewhere classified
C2350266|Terahertz Imaging
C2350266|Imaging, Terahertz
C2350397|Respiratory Gated Imaging Techniques
C2350397|Techniques, Respiratory-Gated Imaging
C2350397|Respiratory-Gated Imaging Techniques
C2350397|Technique, Respiratory-Gated Imaging
C2350397|Imaging Technique, Respiratory-Gated
C2350397|Imaging Techniques, Respiratory-Gated
C2350397|Respiratory-Gated Imaging Technique
C2350397|Gated Imaging Techniques, Respiratory
C0020910|Computer-Assisted Image Interpretation
C0020910|Computer-Assisted Image Interpretations
C0020910|Image Interpretation, Computer-Assisted
C0020910|Image Interpretations, Computer-Assisted
C0020910|Interpretation, Computer-Assisted Image
C0020910|Interpretations, Computer-Assisted Image
C0020910|IMAGE INTERP
C0020910|Image Interpretation, Computer Assisted
C0026018|Microscopies
C0026018|Microscopy
C0026018|Microscopic Examination
C0026018|Microscopy (procedure)
C0026018|Microscopic examination (procedure)
C0026018|MIEXAM
C0026018|Optical microscopy
C0031749|Photographies
C0031749|Photography
C0034606|Imaging, Gamma Camera
C0034606|Imaging, Radionuclide
C0034606|Radionuclide Imaging
C0034606|Isotope scan
C0034606|scintigraphy
C0034606|SCINTIGR
C0034606|Radionuclide Scanning
C0034606|Scan
C0034606|Scanning
C0034606|radionuclide scan
C0034606|radionuclide scan (procedure)
C0034606|Radioisotope scan
C0034606|radionuclide imaging/scanning
C0034606|Radioisotope scans
C0034606|Radionuclide scans
C0034606|Nuclear Scans
C0034606|Radionuclide study
C0034606|Isotope study
C0034606|Radioisotope study
C0034606|Nuclear medicine
C0034606|NM - Nuclear medicine
C0034606|Radioisotope study (procedure)
C0034606|Radionuclide scanning (procedure)
C0034606|Radioisotope scanning
C0034606|nuclear medicine scan
C0034606|radioimaging
C0034606|Radioisotope scan NOS
C0034606|Scintigraphy NOS
C0034606|RI scan
C0034606|Scanning, Radioisotope
C0034606|Gamma Camera Imaging
C0034606|Nuclear medicine imaging procedure (procedure)
C0034606|Nuclear medicine imaging procedure
C0034606|Radionuclide scanning, NOS
C0038603|Subtraction Technics
C0038603|Subtraction Technique
C0038603|Subtraction Techniques
C0038603|Technic, Subtraction
C0038603|Technics, Subtraction
C0038603|Technique, Subtraction
C0038603|Techniques, Subtraction
C0038603|Subtraction Technic
C0039810|Thermography
C0039810|Thermogram
C0039810|THERMOGR
C0039810|Thermography imaging
C0039810|Thermography imaging - action
C0039810|thermography (procedure)
C0039810|Mapping, Temperature
C0039810|Temperature Mappings
C0039810|Mappings, Temperature
C0039810|Thermography NOS
C0039810|Thermography NOS (procedure)
C0039810|Temperature Mapping
C0039810|Thermography technique
C0039810|Thermography imaging - action (qualifier value)
C0039810|Thermography, NOS
C0039810|Thermogram, NOS
C0376519|NIR Spectroscopies
C0376519|Near-Infrared Spectrometries
C0376519|Near-Infrared Spectrometry
C0376519|Near-Infrared Spectroscopies
C0376519|Near-Infrared Spectroscopy
C0376519|Spectrometries, Near-Infrared
C0376519|Spectrometry, Near Infrared
C0376519|Spectroscopies, NIR
C0376519|Spectroscopies, Near-Infrared
C0376519|Spectroscopy, NIR
C0376519|Spectroscopy, Near Infrared
C0376519|Spectroscopy, Near-Infrared
C0376519|NIR spectroscopy
C0376519|near infrared spectrometry
C0376519|near infrared spectroscopy
C0376519|near-infrared spectroscopy (procedure)
C0376519|Spectrometry, Near-Infrared
C0887832|3 D Imaging
C0887832|3-D Imagings
C0887832|Imaging, 3-D
C0887832|Imaging, Three Dimensional
C0887832|Imaging, Three-Dimensional
C0887832|Imagings, 3-D
C0887832|Imagings, Three-Dimensional
C0887832|Three-Dimensional Imaging
C0887832|Three-Dimensional Imagings
C0887832|3D imaging
C0887832|3-D Imaging
C0887832|Medical Imaging, Three Dimensional
C0887832|Three Dimensional Imaging
C1450459|Stroboscopy
C0011923|Diagnostic Imaging
C0011923|DIAG IMAGING
C0011923|IMAGING DIAG
C0011923|Imaging by method
C0011923|Imaging
C0011923|Imaging procedure
C0011923|Diagnostic imaging (procedure)
C0011923|Imaging by method (procedure)
C0011923|Clinical imaging
C0011923|Medical Imaging
C0011923|Imaging, Diagnostic
C0011923|Imaging (procedure)
C0011923|Diagnostic imaging, NOS
C0024485|Magnetic Resonance Imaging
C0024485|Imaging, Magnetic Resonance
C0024485|MRI
C0024485|TOMOGR MR
C0024485|MR TOMOGR
C0024485|NMRI
C0024485|NMR Imaging
C0024485|TOMOGR NMR
C0024485|ZEUGMATOGR
C0024485|Imaging, NMR
C0024485|NMR TOMOGR
C0024485|Magnetic resonance imaging - action
C0024485|NMR
C0024485|Nuclear magnetic resonance imaging
C0024485|MRI Scan
C0024485|Magnetic resonance imaging procedure
C0024485|Nuclear magnetic resonance
C0024485|Nuclear magnetic resonance NOS
C0024485|Nuclear magnetic resonance NOS (procedure)
C0024485|NMR Scan
C0024485|Magnetic resonance study (procedure)
C0024485|Magnetic resonance: [imaging] or [study]
C0024485|Magnetic resonance study
C0024485|Magnetic resonance: [imaging] or [study] (procedure)
C0024485|MRI scan (procedure)
C0024485|Tomography, NMR
C0024485|MR Tomography
C0024485|Tomography, MR
C0024485|Zeugmatography
C0024485|NMR Tomography
C0024485|MR - Magnetic resonance
C0024485|MRI - Magnetic resonance imaging
C0024485|NMR - Nuclear magnetic resonance
C0024485|Magnetic resonance technique
C0024485|Magnetic resonance imaging (procedure)
C0024485|Magnetic resonance imaging - action (qualifier value)
C0024485|Magnetic resonance imaging, NOS
C0024485|MRI, NOS
C0024485|Magnetic Resonance Imaging Scan
C0024485|Medical Imaging, Magnetic Resonance / Nuclear Magnetic Resonance
C0040706|Diaphanoscopies
C0040706|Transillumination
C0040706|Transilluminations
C0040706|Diaphanoscopy
C0040706|Light scanning
C0040706|Transillumination scanning
C0040706|Optical transillumination (procedure)
C0040706|Optical transillumination
C0040706|Optical transillumination, NOS
C0203669|whole body scanning
C0203669|Total body scan
C0203669|Whole Body Scan
C0203669|whole body imaging
C0203669|Total body scan (procedure)
C0203669|Scan NOS whole body
C0203669|Radioisotope scan of total body
C0203669|Radioisotope scan of total body (procedure)
C0203669|Total body scan (procedure) [Ambiguous]
C0203669|Imaging, Whole Body
C0203669|Imagings, Whole Body
C0203669|Scan, Whole Body
C0203669|Scans, Whole Body
C0203669|Whole Body Imagings
C2350395|Cardiac Gated Imaging Techniques
C2350395|Technique, Cardiac-Gated Imaging
C2350395|Techniques, Cardiac-Gated Imaging
C2350395|Imaging Techniques, Cardiac-Gated
C2350395|Cardiac-Gated Imaging Techniques
C2350395|Cardiac-Gated Imaging Technique
C2350395|Imaging Technique, Cardiac-Gated
C0040399|Emission-Computed Tomography, Single-Photon
C0040399|SPECT
C0040399|Tomography, Emission-Computed, Single-Photon
C0040399|Tomography, Single-Photon Emission-Computed
C0040399|single photon emission computed tomography
C0040399|CT SINGLE PHOTON EMISS
C0040399|RADIONUCLIDE TOMOGR SINGLE PHOTON EMISS
C0040399|SINGLE PHOTON EMISS CT
C0040399|EMISS CT SINGLE PHOTON
C0040399|Single photon emission computed tomography - action
C0040399|Single Photon Emission Computer Assisted Tomography
C0040399|Single Photon Emission Computerized Tomography
C0040399|Single Photon Emission CT Scan
C0040399|CT Scan, Single Photon Emission
C0040399|CAT Scan, Single Photon Emission
C0040399|Single photon emission computerised tomogram
C0040399|SPET
C0040399|Single Photon Emission Tomography
C0040399|Radionuclide Tomography, Single Photon Emission Computed
C0040399|Single-photon emission computed tomography
C0040399|Single photon emission computerized tomogram
C0040399|Single photon emission computerised tomography
C0040399|SPECT SCAN
C0040399|Single-Photon Emission CT Scan
C0040399|Single-Photon Emission Computer-Assisted Tomography
C0040399|Radionuclide Tomography, Single-Photon Emission-Computed
C0040399|Single-Photon Emission Computerized Tomography
C0040399|CT Scan, Single-Photon Emission
C0040399|Single-Photon Emission-Computed Tomography
C0040399|CAT Scan, Single-Photon Emission
C0040399|Tomography, Single-Photon, Emission-Computed
C0040399|SPET - Single photon emission computed tomography
C0040399|Single photon emission computed tomography - action (qualifier value)
C0040399|Single photon emission computerized tomography (procedure)
C0040399|tomography, emission computed, single photon
C0040399|SPECT imaging
C0040399|Single photon emission computerized tomography, NOS
C0040399|Medical Imaging, Single Photon Emission Computed Tomography
C0040399|Single photon emission computed tomography (SPECT)
C2717949|Vm Mapping, Optical
C2717949|Mapping, Optical Vm
C2717949|Mappings, Optical Vm
C2717949|Vm Mappings, Optical
C2717949|Voltage-Sensitive Dye Imaging
C2717949|Optical Vm Mappings
C2717949|Imaging, Voltage-Sensitive Dye
C2717949|Voltage Sensitive Dye Imaging
C2717949|Optical Vm Mapping
C2717949|Optical Mapping, Transmembrane Potential
C2717949|Transmembrane Potential Optical Mapping
C2717949|Optical Transmembrane Potential Mapping
C1537028|Imaging, Molecular
C1537028|Molecular Imaging
C1533147|Specific imaging methods NOS (procedure)
C1533147|Specific imaging methods (procedure)
C1533147|Specific imaging methods NOS
C1533147|Specific imaging methods
C0730031|Bone density scan
C0730031|Bone density scan (procedure)
C0006117|Brain Mapping
C0006117|Mapping, Brain
C0006117|Brain mapping (procedure)
C0581609|Radionuclide water and electrolyte study
C0581609|Radionuclide water and electrolyte study (procedure)
C2936236|Imaging Techniques, Cardiac
C2936236|Technique, Cardiac Imaging
C2936236|Cardiac Imaging Techniques
C2936236|Cardiac Imaging Technique
C2936236|Imaging Technique, Cardiac
C2936236|Techniques, Cardiac Imaging
C0581589|Radionuclide urinary tract study
C0581589|Urinary isotope studies
C0581589|Urinary isotope studies (procedure)
C0581589|Radionuclide urinary tract study (procedure)
C0203668|bone scanning
C0203668|Radioisotope scan of bone
C0203668|Bone scan
C0203668|Radioisotope bone scan
C0203668|Scan;bone(s)
C0203668|skeletal imaging
C0203668|bone imaging
C0203668|Radionuclide bone study
C0203668|Radionuclide bone study (procedure)
C0203668|Bone isotope studies
C0203668|isotopic bone scan (procedure)
C0203668|isotopic bone scan
C0203668|Bone scan NOS
C0203668|Scan NOS bone
C0203668|Nuclear medicine imaging bone
C0203668|Isotope bone scan
C0203668|Radioisotope scan of bone (procedure)
C0203668|Radioisotope scan of bone, NOS
C0203668|Bone scan, NOS
C0203668|Bone imaging, NOS
C0203668|skeletal scanning
C0203779|nuclear thyroid imaging (procedure)
C0203779|nuclear thyroid imaging only
C0203779|nuclear thyroid imaging only (procedure)
C0203779|nuclear thyroid imaging
C0203779|thyroid imaging
C0203779|thyroid imaging only
C0203779|Thyroid scan/isotop func
C0203779|radionuclide scan of thyroid
C0203779|radionuclide scan of thyroid (procedure)
C0203779|Thyroid isotope studies
C0203779|Radionuclide thyroid study
C0203779|Radionuclide thyroid study (procedure)
C0203779|Scan thyroid gland
C0203779|Scan NOS thyroid gland
C0203779|Radionuclide thyroid imaging study
C0203779|Thyroid scan and radioisotope function studies
C0203779|Radionuclide thyroid imaging (procedure)
C0203779|Radionuclide thyroid imaging
C0203779|Thyroid scan
C0203779|Thyroid scan and radioisotope function studies, NOS
C0203779|Thyroid scan, NOS
C0430470|Radionuclide study of heart
C0430470|Heart isotope studies
C0430470|Cardiac isotope studies
C0430470|Radionuclide study of heart (procedure)
C0412375|Lymphoscintigraphy
C0412375|lymphoscintigraphy (procedure)
C0412375|Lymphatic system scan
C0412375|Lymphoscintigraphies
C0412375|Radioisotope scan of lymphatic system
C0412375|Radionuclide study of lymphatic system (procedure)
C0412375|Radionuclide lymphogram
C0412375|Lymph isotope studies
C0412375|Radionuclide study of lymphatic system
C0412375|Radioisotope scan of lymphatic system (procedure)
C0412375|Radionuclide lymphogram (procedure)
C0412375|Radionuclide lymphangiogram
C0412375|Scan of lymphatic system
C0412375|Radioisotope scan of lymphatic system (procedure) [Ambiguous]
C0412324|Cystographic isotope studies
C0412324|Cystogr.isotope studies
C0412324|Cystographic isotope studies (procedure)
C1571763|Iron isotope studies
C0412331|CSF isotope study (procedure)
C0412331|Cerebrospinal fluid isotope study (procedure)
C0412331|Cerebrospinal fluid isotope study
C0412331|CSF isotope study
C0412400|radioisotope scan of spleen
C0412400|isotopic scans spleen
C0412400|radioisotope scan of spleen (procedure)
C0412400|Spleen isotope studies
C0412400|Radionuclide spleen studies
C0412400|Spleen scan or function study
C1881134|Image Study
C1881134|Imaging Study
C1881134|imaging studies (procedure)
C1881134|imaging studies
C2985362|ProstaScint Scan
C0162481|Doppler Ultrasound
C0162481|Doppler Ultrasound (procedure)
C0162481|Ultrasound Doppler
C0162481|US.doppler
C0162481|Doppler scan
C0162481|Ultrasound Doppler NOS
C0162481|Diagnostic Doppler ultrasonography
C0162481|Ultrasonic Doppler
C0162481|Diagnostic Doppler ultrasonography (procedure)
C0162481|Diagnostic Doppler ultrasonography, NOS
C0162481|Doppler ultrasound, NOS
C3494219|Optical Imaging
C3494219|Imaging, Optical
C0203790|Thyroid carcinoma metastases imaging; whole body
C0203790|whole body nuclear imaging for metastatic thyroid carcinoma
C0203790|whole body nuclear imaging for metastatic thyroid carcinoma (procedure)
C0203790|THYROID MET IMAGING BODY
C0203790|THYROID CARCINOMA METASTASES IMG WHOLE BODY
C0203790|Thyroid imaging for metastatic carcinoma, whole body
C0203790|Thyroid imaging for metastatic carcinoma, whole body (procedure)
C1299233|Radionuclide bone marrow study
C1299233|Scan bone marrow
C1299233|Radioisotope scan of bone marrow
C1299233|Radioisotope scan of bone marrow (procedure)
C1299233|Bone marrow scan or function study
C0203788|Chest imaging for metastatic carcinoma of thyroid
C0203788|Chest imaging for metastatic carcinoma of thyroid (procedure)
C0581646|X-ray face eyes
C0581646|x-ray of eye (procedure)
C0581646|x-ray of eye
C0581646|X-ray;eye
C0581646|Ophthalmic plain film
C0581646|Ophthalmic plain film (procedure)
C0203382|Carotid imaging
C0203382|Imaging of carotid arteries (procedure)
C0203382|Imaging of carotid arteries
C0203382|Imaging of carotid arteries, NOS
C0200189|eye fundus photography
C0200189|Fundus photography
C0200189|fundus photography (procedure)
C0200189|Ocular fundus photography
C0200189|Ocular fundus photography (procedure)
C0031753|Photomicrographies
C0031753|Photomicrography
C0031753|PHOTOMICROGR
C0031753|Photography, microscopic (procedure)
C0031753|Photography, microscopic
C0031753|Photography, microscopic, NOS
C0031753|Photomicrography, NOS
C0203787|Neck imaging for metastatic carcinoma of thyroid
C0203787|Neck imaging for metastatic carcinoma of thyroid (procedure)
C1443932|Radiologic procedure on chest
C1443932|Radiologic procedure on chest (procedure)
C0203793|Adrenal imaging
C0203793|Adrenal imaging (procedure)
C0203793|Adrenal imaging, NOS
C3665374|Diagn. nuclear medicine NOS
C3665374|diagnostic service sources radiology labs radionuclide imaging
C3665374|diagnostic service sources radiology labs radionuclide imaging (procedure)
C3665374|radionuclide imaging
C3665374|Diagnostic nuclear medicine procedures
C3665374|Diagnostic nuclear medicine NOS
C3665374|Diagnostic nuclear medicine NOS (procedure)
C3665374|Diagnostic nuclear med.
C3665374|Isotope diagnostic rad.
C3665374|Nuclear med.-diagnostic
C3665374|Isotope diagnostic radiology
C3665374|Diagnostic nuclear medicine
C3665374|Nuclear medicine diagnostic procedure (procedure)
C3665374|Diagn. nuclear medicine NOS (procedure)
C3665374|Diagnostic radionuclide study
C3665374|Nuclear medicine diagnostic procedure
C3665374|Diagnostic nuclear medicine procedure
C3665374|Isotope study
C3665374|Diagnostic radionuclide study, NOS
C0204141|Diagnostic dental photographs
C0204141|Diagnostic dental photography (procedure)
C0204141|Diagnostic dental photography
C0007800|Cerebral Ventriculographies
C0007800|Cerebral Ventriculography
C0007800|Ventriculographies, Cerebral
C0007800|ventriculography
C0007800|VENTRICULOGR CEREBRAL
C0007800|CEREBRAL VENTRICULOGR
C0007800|brain ventriculography
C0007800|Ventriculography, Cerebral
C0007800|Ventriculography of brain
C0007800|Cerebral ventriculography (procedure)
C0007800|Ventriculography of brain (procedure)
C0007800|Ventriculogram
C1533606|Endoscopy of pancreas, NOS
C1533606|Endoscopy of pancreas (procedure)
C1533606|Endoscopy of pancreas
C1533606|Endoscopy of pancreas (procedure) [Ambiguous]
C0016313|Fluorescein Angiography
C0016313|FA - Fluorescein angiogram
C0016313|Fluorescein angiogram
C0016313|FLUORESCEIN ANGIOGR
C0016313|ANGIOGR FLUORESCEIN
C0016313|fluorescein angiography of eye (procedure)
C0016313|fluorescein angiography of eye
C0016313|Angiography, Fluorescein
C0431056|Clinical photography, NOS
C0431056|Medical photography of patient, NOS
C0431056|Photography of patient (procedure)
C0431056|Medical photography (procedure)
C0431056|Photography of patient
C0431056|Medical photography
C0431056|Clinical photography
C0431056|Photography of patient (procedure) [Ambiguous]
C0412379|Radionuclide salivary gland imaging procedure
C0412379|Salivary gland imaging
C0412379|Radionuclide salivary gland study
C0412379|Salivary gland imaging (procedure)
C0412379|Radionuclide salivary gland imaging procedure (procedure)
C0202639|Muscle thermography
C0202639|muscle thermography (procedure)
C0203042|Placentography
C0203042|Placentography NOS (procedure)
C0203042|Placentography NOS
C0203042|Placentography (procedure)
C0203042|Placentogram
C0203042|Placental imaging
C0009618|Computer Assisted Image Analysis
C0009618|Computer-Assisted Image Analyses
C0009618|Image Analyses, Computer-Assisted
C0009618|Image Analysis, Computer Assisted
C0009618|COMPUTER ASSISTED IMAGE ANAL
C0009618|IMAGE ANAL COMPUTER ASSISTED
C0009618|ANAL COMPUTER ASSISTED IMAGE
C0009618|Analysis, Computer-Assisted Image
C0009618|Computer-Assisted Image Analysis
C0009618|Computer assisted image analysis (procedure)
C0009618|Image Analysis, Computer-Assisted
C0438661|Clinical X-ray application NOS
C0438661|Clinical X-ray application NOS (procedure)
C0438661|Clinical X-ray application NOS (situation)
C0408190|Examination of joint under image intensifier
C0408190|Examination of joint under image intensifier (procedure)
C1293911|Ocular photography AND/OR evaluation (procedure)
C1293911|Ocular photography AND/OR evaluation
C0184973|Endoscopy and photography
C0184973|Endoscopy and photography (procedure)
C0559963|Retinal photography (procedure)
C0559963|Retinal photography
C0559963|Photography;retinal
C0203300|magnetic resonance imaging of joint of lower extremity
C0203300|magnetic resonance imaging of joint of lower extremity (procedure)
C0203300|MRI of joint of lower extremity
C0203391|Imaging of arteries of extremities (procedure)
C0203391|Imaging of arteries of extremities
C0203391|Imaging of arteries of extremities, NOS
C0560563|Fluoroscopic guidance
C0560563|procedure with fluoroscopic guidance
C0560563|procedure with fluoroscopic guidance (treatment)
C0560563|Fluoroscopic guidance (procedure)
C0454120|radiation therapy treatment planning using magnetic resonance imaging (treatment)
C0454120|radiation therapy treatment planning using magnetic resonance imaging
C0454120|Radiotherapy planning MRI scan
C0454120|Radiotherapy planning using magnetic resonance imaging
C0454120|Radiotherapy planning using magnetic resonance imaging (procedure)
C0411316|Therapeutic barium enema
C0411316|Enema for intussusception
C0411316|Therapeutic barium enema (procedure)
C0411330|Percutaneous imaging guided therapeutic drainage
C0411330|Percutaneous imaging guided therapeutic drainage (procedure)
C0202726|MRI TMJ
C0202726|magnetic resonance imaging of temporomandibular joint
C0202726|magnetic resonance imaging of temporomandibular joint (procedure)
C0202726|MAGNETIC IMAGE JAW JOINT
C0202726|Magnetic resonance (eg, proton) imaging, temporomandibular joint(s)
C0202726|MRI TEMPOROMANDIBULAR JOINT
C0202726|MRI of temporomandibular joint
C0202726|MRI of temporomandibular joints
C0202726|MRI scan of jaw joints
C0203854|Testicular imaging
C0203854|Testicular imaging (procedure)
C0412751|Miscellaneous imaging procedures
C0412751|Miscellaneous imaging procedures (procedure)
C0203256|MRI of joint of upper extremity
C0203256|Magnetic resonance imaging of joint of upper extremity
C0203256|Magnetic resonance imaging of joint of upper extremity (procedure)
C0456852|Image-Guided Biopsies
C0456852|Biopsy, Imaging Guided
C0456852|Image Guided Biopsy
C0456852|Biopsy, Image-Guided
C0456852|Imaging Guided Biopsies
C0456852|Guided Biopsy, Imaging
C0456852|Guided Biopsies, Imaging
C0456852|Image-Guided Biopsy
C0456852|Biopsies, Image-Guided
C0456852|Biopsies, Imaging Guided
C0456852|Imaging Guided Biopsy
C0456852|Imaging guided biopsy (procedure)
C1513743|Multimodal Imaging
C1513743|Imagings, Multimodal
C1513743|Multimodal Imagings
C1513743|Imaging, Multimodal
C1513743|Multimodality
C2047967|3-dimensional rendering
C2047967|imaging study with 3-dimensional rendering
C2047967|3-D rendering
C2047967|imaging study with 3-dimensional rendering (procedure)
C2015796|other imaging studies (procedure)
C2015796|other imaging studies
C3697941|Postmortem imaging procedure (procedure)
C3697941|Postmortem imaging procedure
C3687804|Post Processing of Image or Image Sets
C3534891|Image Capture Only
C3642491|Image Capture With Interpretation
C3534890|Interpretation and Report Only
C3898703|Intraoperative Imaging
C3897151|X-Ray PCI
C3897151|Phase-Contrast X-Ray Imaging
C3897151|Phase-Sensitive X-Ray Imaging
C3897151|X-Ray Phase-Contrast Imaging
C3898624|Laser Doppler Imaging
C3898624|Scanning Laser Doppler
C1328868|Diffuse Optical Tomography
C3897187|Video-Based 3-Dimensional Surface Imaging
C3897187|Video-Based 3D Surface Imaging
C0430876|Fluorescence imaging
C0430876|Imaging, Fluorescence
C0430876|Fluorescence imaging (procedure)
C0430876|Ophthalmic fluorescence imaging
C3898640|Kv/Mv Imaging
C3897255|Ultrasound Tomography
C3889415|Biodynamic Imaging
C3889415|BDI
C3899943|Bioelectric Field Imaging
C3897003|Dynamic Contrast-Enhanced Ultrasound Imaging
C3898477|Magnetic Resonance Thermal Imaging
C3899379|Diffuse Optical Imaging
C3854375|Laser speckle contrast imaging
C3854375|LSCI
C3854375|Laser Speckle Imaging
C3898096|Optical Doppler Tomography
C3897256|Ultrasound Elasticity Imaging
C3897929|Photoacoustic Imaging
C3898216|Multispectral Imaging
C3897769|Real-Time Position-Tracking Imaging
C4064207|reflectance confocal microscopy
C4064207|reflectance confocal microscopy (procedure)
C0412412|Renal scan/isotope funct
C0412412|Renal scan
C0412412|Renal isotope studies
C0412412|Kidney isotope studies
C0412412|Radionuclide dynamic renal study
C0412412|Kidney radioisotope scan
C0412412|Renal isotope studies (procedure)
C0412412|Radionuclide dynamic renal study (procedure)
C0412412|Renal scan and radioisotope function study
C0412412|Radionuclide renal studies
C0412412|Kidney imaging with function study (procedure)
C0412412|Renal radioisotope scan
C0412412|Kidney imaging with function study
C0412412|Renal scan NOS
C0412412|Scan NOS renal
C0412412|radionuclide renal function study
C0412412|Isotopic renogram
C0412412|Kidney scan
C0412412|Isotopic renogram, NOS
C0442972|Imaging guidance procedure
C0442972|Imaging guidance
C0442972|Imaging guidance (procedure)
C0442972|Imaging guidance procedure (procedure)
C1299525|Imaging by body site (procedure)
C1299525|Imaging by body site
C0203512|Special dosimetry
C0203512|radiation therapy special dosimetry (treatment)
C0203512|radiation therapy special dosimetry
C0203512|Special dosimetry (procedure)
C0203512|Special dosimetry, NOS
C1299527|Video imaging procedure
C1299527|Video imaging procedure (procedure)
C1299527|Video imaging
C0411282|Endovascular radiologic intervention
C0411282|Endovascular intervention
C0411282|Endovascular therapeutic radiology
C0411282|Endovascular radiological intervention
C0411282|Endovascular radiologic intervention (procedure)
C0411282|Endovascular intervention (procedure)
C0400689|Endoscopic retrograde cholangiography and biopsy of lesion of bile duct
C0400689|Endoscopic retrograde cholangiography and biopsy of lesion of bile duct (procedure)
C0412467|Metabolic studies
C0412467|Radionuclide metabolic studies
C0412467|Radionuclide metabolic studies (procedure)
C1266825|Nuclear medicine diagnostic procedure on endocrine AND/OR haematopoietic system
C1266825|Nuclear medicine diagnostic procedure on endocrine AND/OR hematopoietic system (procedure)
C1266825|Nuclear medicine diagnostic procedure on endocrine AND/OR hematopoietic system
C0412323|Isotope uptake/excretion studies
C0412323|Isotope uptake/excretion studies (procedure)
C0400803|Endoscopic retrograde cholangiopancreatography and biopsy of lesion of ampulla of Vater
C0400803|Endoscopic retrograde cholangiopancreatography and biopsy of lesion of ampulla of Vater (procedure)
C0203639|Radionuclide special dynamic function study (procedure)
C0203639|Radionuclide special dynamic function study
C0203639|Radionuclide special dynamic function study, NOS
C0581576|Regional nuclear medicine
C0581576|Regional nuclear medicine (procedure)
C0473940|Blood isotope studies
C0473940|Radionuclide studies in haematology
C0473940|Radionuclide studies in hematology
C0473940|Radionuclide studies in hematology (procedure)
C0400540|Endoscopic retrograde pancreatography and biopsy of lesion of pancreas
C0400540|Endoscopic retrograde pancreatography and biopsy of lesion of pancreas (procedure)
C0203831|Radionuclide study, protein kinetics
C0203831|Radionuclide study, protein kinetics (procedure)
C0203647|Radionuclide volume dilution study (procedure)
C0203647|Radionuclide volume dilution study
C0203647|Radionuclide volume dilution study, NOS
C0203646|Radionuclide dynamic function study with multiple probes (procedure)
C0203646|Radionuclide dynamic function study with multiple probes
C0203646|Radionuclide dynamic function study with multiple probes, NOS
C1831737|infrared thermography
C1522706|1H-nuclear magnetic resonance spectroscopic imaging
C1522706|magnetic resonance spectroscopic imaging
C1522706|proton magnetic resonance spectroscopic imaging
C1522706|Magnetic Resonance Spectroscopy
C1522706|MRS
C1522706|MRSI
C1522706|MRS Imaging
C1522706|1H- Nuclear Magnetic Resonance Spectroscopic Imaging
C1510486|DEXA
C1510486|DXA
C1510486|Dual X-Ray Absorptiometry
C1510486|Dual-Energy X-Ray Absorptiometry
C1510486|DEXA scan
C1510486|Dual Energy X Ray Absorptiometry
C1510486|X Ray Absorptiometry, Dual Energy
C1510486|Dual X Ray Absorptiometry
C1510486|X-Ray Absorptiometry, Dual
C1510486|Absorptiometry, Dual X Ray
C1510486|Absorptiometries, DPX
C1510486|Absorptiometry, DPX
C1510486|Absorptiometry, Dual Energy X Ray
C1510486|Dual Energy X-ray Absorptiometry
C1510486|DXA SCAN
C1510486|dual energy x-ray absorptiometric scan
C1510486|bone mineral density scan
C1510486|BMD scan
C1510486|Dual X-Ray Absorptometry
C1510486|Absorptiometry, Dual-Energy X-Ray
C1510486|Absorptiometry, Dual X-Ray
C1510486|X-Ray Absorptiometry, Dual-Energy
C1510486|DPX Absorptiometry
C0920367|optical coherence tomography
C0920367|TOMOGR OPTICAL COHERENCE
C0920367|OPTICAL COHERENCE TOMOGR
C0920367|OCT TOMOGR
C0920367|optical coherence tomography (procedure)
C0920367|Doppler OCT
C0920367|Tomography, Optical Coherence
C0920367|OCT
C0920367|OCT Tomography
C0920367|Tomography, OCT
C0920367|Coherence Tomography, Optical
C0920367|OCT - Optical coherence tomography
C0037812|Spectrum Analysis
C0037812|spectroscopy
C0037812|SPECTRUM ANAL
C0037812|ANAL SPECTRUM
C0037812|Analysis, Spectrum
C1514690|Radiation Ionizing, Diagnostic Imaging
C1455714|Thallium stress test
C1455714|Exercise Thallium
C1455714|Stress Thallium Test
C1455714|Thallium Myocardial Perfusion Imaging Stress Test
C1455714|Thallium stress test with or without transesophageal pacing
C1881135|Imaging Biomarker Analysis
C1514691|Radiation Non-Ionizing, Diagnostic Imaging
C0400786|ERCP sphincterotomy sphincter of Oddi and calculus removal (procedure)
C0400786|ERCP sphincterotomy sphincter of Oddi and calculus removal
C0400786|Endoscopic retrograde cholangiopancreatography sphincterotomy sphincter of Oddi and calculus removal (procedure)
C0400786|Endoscopic retrograde cholangiopancreatography sphincterotomy sphincter of Oddi and calculus removal
C0400786|Endoscopic retrograde cholangiopancreatography (ERCP) sphincterotomy sphincter of Oddi and calculus removal
C0400786|Endoscopic retrograde cholangiopancreatography (ERCP) sphincterotomy sphincter of Oddi and calculus removal (procedure)
C2348290|Digital Image Analysis
C2346479|Implanted Fiducial-Based Imaging System
C2349125|Vibration Response Imaging
C2348715|Frequency-Domain Photon Migration
C2348715|FDPM
C2094547|radionuclide scan of liver and spleen with vascular flow (procedure)
C2094547|radionuclide scan of liver and spleen with vascular flow
C0361418|Technetium[99mTc] tin colloid injection BP (product)
C0361418|Technetium[99mTc] tin colloid injection BP
C0361418|Technetium[99mTc] tin colloid injection BP (substance)
C0361413|Technetium[99mTc] albumin millimicrospheres injection (product)
C0361413|Technetium[99mTc] albumin millimicrospheres injection
C0361413|Technetium[99mTc] albumin millimicrospheres injection (substance)
C0361331|Technetium[99mTc] rhenium sulfide colloid injection (product)
C0361331|Technetium[99mTc] rhenium sulphide colloid injection
C0361331|Technetium[99mTc] rhenium sulfide colloid injection
C0361331|Technetium[99mTc] rhenium sulfide colloid injection (substance)
C0361420|Technetium[99mTc] albumin colloid injection
C0361420|Technetium[99mTc] albumin colloid injection (product)
C0361420|Technetium[99mTc] albumin colloid injection (substance)
C1444888|Technetium[99mTc] sulfur colloid diagnostic kit
C1444888|Technetium[99mTc] sulfur colloid injection (product)
C1444888|Technetium[99mTc] sulfur colloid injection
C1444888|Technetium[99mTc] sulphur colloid diagnostic kit
C1444888|Technetium[99mTc] sulphur colloid injection
C2314954|Magnetic resonance imaging (MRI) of liver with contrast
C2314954|Magnetic resonance imaging of liver with contrast (procedure)
C2314954|abdominal MRI liver with contrast
C2314954|magnetic resonance imaging of liver with contrast
C2314954|MRI of liver with contrast
C2318037|abdominal MRI liver without contrast
C2318037|magnetic resonance imaging of liver without contrast (procedure)
C2318037|magnetic resonance imaging of liver without contrast
C2318039|abdominal MRI liver without, then with contrast
C2318039|magnetic resonance imaging of liver without, then with contrast (procedure)
C2318039|magnetic resonance imaging of liver without, then with contrast
C2584955|Ablation of liver using magnetic resonance imaging guidance (procedure)
C2584955|MRI guided ablation of liver
C2584955|Ablation of liver using magnetic resonance imaging guidance
C2711639|Magnetic resonance imaging of heart and liver for assessment of cardiac and hepatic iron load (procedure)
C2711639|Magnetic resonance imaging of heart and liver for assessment of cardiac and hepatic iron load
C2711639|MRI of heart and liver for assessment of cardiac and hepatic iron load
C2094545|radionuclide scan of liver and spleen (procedure)
C2094545|radionuclide scan of liver and spleen
C2094546|static radionuclide scan of liver and spleen (procedure)
C2094546|static radionuclide scan of liver and spleen
C2315791|Magnetic resonance imaging (MRI) of liver and biliary tract with contrast
C2315791|Hepatobiliary magnetic resonance imaging (MRI) with contrast
C2315791|Magnetic resonance imaging of liver and biliary tract with contrast (procedure)
C2315791|Magnetic resonance imaging of liver and biliary tract with contrast
C2315791|MRI of liver and biliary tract with contrast
C2584862|Focused ultrasound ablation of liver using magnetic resonance imaging guidance (procedure)
C2584862|Focused ultrasound ablation of liver using magnetic resonance imaging guidance
C2584862|MRI guided focused ultrasound ablation of liver
