C0020538|Hypertensive disease
C1963138|Hypertension Adverse Event	
C0085580|Essential hypertension
C0085580|primary hypertension
C0085580|Essential (primary) hypertension
C0085580|HYPERTENSION, ESSENTIAL
C0085580|idiopathic hypertension
C0085580|essential hypertension (diagnosis)
C0085580|Hypertension NOS
C0085580|Hypertension;essential
C0085580|Essential hypertension (disorder)
C0085580|Essential hypertension NOS (disorder)
C0085580|Essential hypertension NOS
C0085580|EHT
C0085580|Essential hypertension, unspecified
C0085580|Unspecified essential hypertension
C0085580|Systemic primary arterial hypertension
C0085580|Essential hypertension, NOS
C0085580|Primary hypertension, NOS
C0020541|Hypertension, Portal
C0020541|Hypertensions, Portal
C0020541|Portal Hypertensions
C0020541|Portal hypertension
C0020541|portal hypertension (diagnosis)
C0020541|Hypertension, Portal [Disease/Finding]
C0020541|Hypertension;portal
C0020541|Portal hypertension (disorder)
C0020541|Hypertension portal
C0020541|PHT - Portal hypertension
C0020541|hypertension; portal
C0020541|portal; hypertension
C0020542|Hypertension, Pulmonary
C0020542|pulmonary hypertension
C0020542|Pulmonary artery hypertension
C0020542|HYPERTENSION PULM
C0020542|PULM HYPERTENSION
C0020542|pulmonary hypertension (diagnosis)
C0020542|Hypertension, Pulmonary [Disease/Finding]
C0020542|Pulmonary hypertension NOS
C0020542|Pulmonary hypertensions
C0020542|Hypertension pulmonary
C0020542|Cardio/pulm: Pulmonary hypertension
C0020542|PHT - Pulmonary hypertension
C0020542|Pulmonary hypertension (disorder)
C0020542|hypertension; pulmonary
C0020542|pulmonary; hypertension
C0020542|Pulmonary hypertension, NOS
C0020544|Hypertension, Renal
C0020544|Hypertensions, Renal
C0020544|Renal Hypertensions
C0020544|Renal Hypertension
C0020544|Hypertension, Renal [Disease/Finding]
C0020544|Hypertension;cardiorenal
C0020544|secondary hypertension to renal disorders
C0020544|hypertension secondary to renal disorders
C0020544|hypertension secondary to renal disorders (diagnosis)
C0020544|Renal hypertension NOS
C0020544|Hypertension renal
C0020544|Renal hypertension (disorder)
C0020544|cardiorenal; hypertension
C0020544|hypertension; renal
C0020544|renal; hypertension
C0264641|Endocrine hypertension
C0264641|adrenal hypertension
C0264641|Endocrine hypertension (disorder)
C0264641|endocrine; disorder hypertension
C0264641|hypertension; endocrine disorders
C0596515|environment associated hypertension
C0598428|familial hypertension
C0598428|congenital hypertension
C0598428|genetic hypertension
C0597048|neurogenic hypertension
C0596088|angiotensin/renin/aldosterone hypertension
C0032914|Pre Eclampsia
C0032914|Pre-Eclampsia
C0032914|preeclampsia
C0032914|Pre-eclampsia, unspecified
C0032914|PREECLAMPSIA/ECLAMPSIA 1
C0032914|PEE1
C0032914|PREGN TOXEMIAS
C0032914|pre-eclampsia (diagnosis)
C0032914|Unspecified pre-eclampsia, unspecified trimester
C0032914|Unspecified pre-eclampsia
C0032914|EPH Gestosis
C0032914|Hypertension-Edema-Proteinuria Gestosis
C0032914|Pre-Eclampsia [Disease/Finding]
C0032914|Pregnancy Toxemias
C0032914|EPH Toxemias
C0032914|Edema-Proteinuria-Hypertension Gestosis
C0032914|Toxemias, Pregnancy
C0032914|EPH Complex
C0032914|Proteinuria-Edema-Hypertension Gestosis
C0032914|Gestosis, EPH
C0032914|Toxaemia (in);pregnancy
C0032914|pregnancy toxemia/hypertension
C0032914|pregnancy toxemia
C0032914|Toxemia Of Pregnancy
C0032914|Toxemia
C0032914|Toxaemia NOS
C0032914|EPH - Oedema, proteinuria and hypertension of pregnancy
C0032914|Pre-eclampsia NOS (disorder)
C0032914|Toxemia NOS (disorder)
C0032914|Toxaemia of pregnancy
C0032914|Pre-eclamptic toxaemia
C0032914|Toxemia NOS
C0032914|Proteinuric hypertension of pregnancy (disorder)
C0032914|Pre-eclampsia (disorder)
C0032914|Pre-eclampsia NOS
C0032914|EPH - Edema, proteinuria and hypertension of pregnancy
C0032914|PET - Pre-eclamptic toxaemia
C0032914|PET - Pre-eclamptic toxemia
C0032914|PE - Pre-eclampsia
C0032914|Proteinuric hypertension of pregnancy
C0032914|Pre-eclamptic toxemia
C0032914|PEE
C0032914|PREG1
C0032914|Hypertensive disorder of pregnancy
C0032914|Pre-eclampsia toxaemia
C0032914|Pre-eclampsia toxemia
C0032914|Of Pregnancy, Toxemia
C0032914|1s, Preeclampsia Eclampsia
C0032914|Of Pregnancies, Toxemia
C0032914|Preeclampsia Eclampsia 1
C0032914|Eclampsia 1, Preeclampsia
C0032914|Pregnancies, Toxemia Of
C0032914|Pregnancy, Toxemia Of
C0032914|Toxemia Of Pregnancies
C0032914|Eclampsia 1s, Preeclampsia
C0032914|1, Preeclampsia Eclampsia
C0032914|Preeclampsia Eclampsia 1s
C0032914|Toxemia of pregnancy (disorder)
C0032914|maternal; toxemia
C0032914|pre-eclamptic; toxemia
C0032914|pregnancy; pre-eclampsia
C0032914|pregnancy; toxemia
C0032914|toxemia; maternal
C0032914|toxemia; pre-eclamptic
C0032914|toxemia; pregnancy
C0032914|Pre-eclampsia, NOS
C0032914|Pre-eclamptic toxemia, NOS
C0032914|Toxemia of pregnancy, NOS
C0032914|Toxaemia of pregnancy, NOS
C0032914|Edema Proteinuria Hypertension Gestosis
C0032914|EPH Toxemia
C0032914|Gestosis, Edema-Proteinuria-Hypertension
C0032914|Gestosis, Hypertension-Edema-Proteinuria
C0032914|Gestosis, Proteinuria-Edema-Hypertension
C0032914|Hypertension Edema Proteinuria Gestosis
C0032914|Proteinuria Edema Hypertension Gestosis
C0032914|Toxemia, EPH
C0032914|Toxemia, Pregnancy
C0032914|Toxemias, EPH
C0032914|Pre-eclamptic NOS
C0032914|Toxemia (in);pregnancy
C0032914|toxemia in pregnancy
C0032914|toxaemia in pregnancy
C0810002|Hypertension with complications and secondary hypertension
C0152105|Hypertensive heart disease
C0152105|hypertensive heart disease (diagnosis)
C0152105|Hypertensive heart disease NOS
C0152105|Hypertension;heart disease
C0152105|Hypertensive heart disease NOS (disorder)
C0152105|Hypertensive heart disease (disorder)
C0152105|Hypertensive heart disease, unspecified
C0152105|Unspecified hypertensive heart disease
C0152105|Hypertensive cardiopathy
C0152105|Hypertensive cardiovascular disease
C0152105|HHD - Hypertensive heart disease
C0152105|heart; hypertension
C0152105|Hypertensive heart disease, NOS
C0848548|Hypertensive renal disease
C0848548|HYPERTENSIVE NEPHROPATHY
C0848548|hypertensive nephropathy (diagnosis)
C0848548|hypertensive kidney disease (diagnosis)
C0848548|hypertensive kidney disease
C0848548|Hypertensive renal disease NOS
C0848548|Hypertension;renal disease
C0848548|Hypertension;nephropathy
C0848548|HNP1
C0848548|Hypertensive renal disease NOS (disorder)
C0848548|Hypertensive renal disease, unspecified
C0848548|Nephropathy hypertensive
C0848548|Hypertensive renal disease (disorder)
C0848548|renal disease; hypertension
C0848548|Hypertensive nephropathy, NOS
C0848548|Hypertensive renal disease, NOS
C0848548|hypertension secondary to renal disease
C0155601|Hypertensive heart and renal disease
C0155601|Hypertensive heart and renal disease NOS
C0155601|Hypertensive heart and renal disease, unspecified
C0155601|cardiorenal disease
C0155601|Hypertensive heart AND renal disease (disorder)
C0155601|Hypertensive heart and renal disease NOS (disorder)
C0155601|hypertensive heart disease; with hypertensive kidney disease
C0155601|kidney; hypertension, with hypertensive heart disease
C0155601|Cardiorenal disease, NOS
C0155601|Hypertensive heart and renal disease, NOS
C0155601|Hypertensive heart AND renal disease [dup] (disorder)
C0155616|Secondary hypertension
C0155616|Secondary hypertension, unspecified
C0155616|unspecified secondary hypertension (diagnosis)
C0155616|secondary hypertension (diagnosis)
C0155616|unspecified secondary hypertension
C0155616|Secondary hypertension (disorder)
C0155616|Secondary hypertension NOS
C0155616|Secondary hypertension NOS (disorder)
C0155616|Hypertension secondary
C0155616|hypertension; secondary
C0155616|secondary; hypertension
C0155616|Secondary hypertension, NOS
C0155616|Hypertension;secondary
C0020540|Hypertension, Malignant
C0020540|Malignant Hypertension
C0020540|Accelerated hypertension
C0020540|Hypertension, Malignant [Disease/Finding]
C0020540|Hypertension;malignant
C0020540|Malignant hypertension (disorder)
C0020540|hypertension (systemic) malignant
C0020540|malignant hypertension (diagnosis)
C0020540|Hypertension malignant
C0020540|Malignant hypertension NOS
C0852036|HYPERTENSION, PREGNANCY-INDUCED
C0852036|HYPERTENSION PREGN IND
C0852036|pregnancy-induced hypertension
C0852036|pregnancy-induced hypertension (diagnosis)
C0852036|Pregnancy associated hypertension
C0852036|Induced Hypertension, Pregnancy
C0852036|Induced Hypertensions, Pregnancy
C0852036|Hypertensions, Pregnancy Induced
C0852036|gestational hypertension NOS
C0852036|Hypertension, Pregnancy-Induced [Disease/Finding]
C0852036|Gestational Hypertension
C0852036|Pregnancy Induced Hypertension
C0852036|Hypertension of pregnancy
C0852036|Hypertension of pregnancy NOS
C0852036|Hypertension induced by pregnancy
C0852036|Hypertension induced by pregnancy (disorder)
C0852036|Hypertension of preg.
C0852036|Hypertension of pregnancy NOS (disorder)
C0852036|Hypertension gestational
C0852036|Gestational hypertension (disorder)
C0852036|PIH Pregnancy induced hypertension
C0852036|GH - Gestational hypertension
C0852036|PIH - Pregnancy-induced hypertension
C0852036|Pregnancy-induced hypertension (disorder)
C0852036|pregnancy; hypertension
C0852036|Pregnancy-induced hypertension, NOS
C0852036|Hypertension, Gestational
C0852036|Hypertension, Pregnancy Induced
C0020538|High blood pressure
C0020538|Hypertension
C0020538|Hypertensive diseases
C0020538|Systemic hypertension
C0020538|Hypertensive disorder, systemic arterial
C0020538|HTN
C0020538|hyperpiesia
C0020538|hyperpiesis
C0020538|Hypertensive disease
C0020538|systemic HTN
C0020538|systemic hypertension (diagnosis)
C0020538|HBP
C0020538|HT
C0020538|Surg comp - hypertension
C0020538|Blood Pressure, High
C0020538|Hypertension [Disease/Finding]
C0020538|Hypertensive diseases (I10-I15)
C0020538|Complications affecting other specified body systems, not elsewhere classified, hypertension
C0020538|Hypertensive disease NOS (disorder)
C0020538|Hypertensive disease NOS
C0020538|Hypertension NOS
C0020538|Hypertensive disease (disorder)
C0020538|(Hypertensive disease) or (hypertension)
C0020538|(Hypertensive disease) or (hypertension) (disorder)
C0020538|[X]Hypertensive diseases (disorder)
C0020538|[X]Hypertensive diseases
C0020538|Increased Blood Pressure
C0020538|Blood Pressure, Increased
C0020538|Pressure, High Blood
C0020538|Elevated blood pressure
C0020538|Hypertension arterial
C0020538|Blood pressure high
C0020538|Cardio/pulm: Hypertensive disorder
C0020538|Hypertensive vascular degeneration
C0020538|Hypertensive vascular disease
C0020538|BP - High blood pressure
C0020538|High blood pressure disorder
C0020538|Systemic arterial hypertension
C0020538|HBP - High blood pressure
C0020538|BP+ - Hypertension
C0020538|HT - Hypertension
C0020538|Hypertensive disorder, systemic arterial (disorder)
C0020538|Hypertensive disorder
C0020538|HTN - Hypertension
C0020538|blood pressure; high
C0020538|high; arterial tension
C0020538|high; blood pressure
C0020538|Hypertension, NOS
C0020538|Hypertensive disease, NOS
C0020538|Raised blood pressure (disorder)
C0020538|Blood Pressures, High
C0020538|High Blood Pressures
C0020538|Vascular Hypertensive Disorder
C0745138|Hypertensive urgency (disorder)
C0745138|Hypertensive urgency
C0745138|hypertensive urgency (diagnosis)
C3695318|Hypertensive chronic kidney disease
C3695318|hypertensive chronic kidney disease (diagnosis)
C3695318|Hypertensive chronic kidney disease NOS
C3695318|Chronic kidney disease due to hypertension
C3695318|Chronic kidney disease due to hypertension (disorder)
C3695318|Hypertensive chronic kidney disease (disorder)
C1719469|Hypertensive heart and chronic kidney disease
C1719469|hypertensive heart and chronic kidney disease (diagnosis)
C1719469|Hypertensive heart and chronic kidney disease (disorder)
C2169401|reactive hypertension
C2169401|reactive hypertension (diagnosis)
C2931417|Faye-Petersen Ward Carey syndrome
C1171349|Kallikrein attenuated hypertension
C1171349|Kallikrein hypertension
C2931778|Tachycardia hypertension microphthalmos hyperglycinuria
C2931778|Adams Nance syndrome
C0152132|Hypertensive Retinopathy
C0152132|hypertensive retinopathy (diagnosis)
C0152132|Retinopathy hypertensive
C0152132|Retinopathy, Hypertensive
C0152132|Hypertensive Retinopathies
C0152132|Retinopathies, Hypertensive
C0152132|Retinopathy;hypertensive
C0152132|Hypertensive Retinopathy [Disease/Finding]
C0152132|Hypertensive retinopathy (disorder)
C0152132|Hypertensive retinopathy [Ambiguous]
C0745121|iatrogenic hypertension (diagnosis)
C0745121|iatrogenic hypertension
C0262534|white coat hypertension
C0262534|Clinic Hypertension, Isolated
C0262534|Syndrome, White Coat
C0262534|Hypertension, White Coat
C0262534|Hypertension, Isolated Clinic
C0262534|White Coat Hypertension [Disease/Finding]
C0262534|White Coat Syndrome
C0262534|Isolated Clinic Hypertension
C0262534|White coat hypertension (disorder)
C0262534|Labile hypertension due to being in a clinical environment (disorder)
C0262534|Labile hypertension due to being in a clinical environment
C0262534|Hypertension;white coat
C3178811|Hypertension, Masked
C3178811|Hypertensions, Masked
C3178811|Masked Hypertension
C3178811|Masked Hypertensions
C3178811|Masked Hypertension [Disease/Finding]
C2186383|reported a history of intermittent hypertension
C2186383|reported history of intermittent hypertension (history)
C2186383|reported history of intermittent hypertension
C2186383|intermittent hypertension
C0745136|Hypertensive emergency (disorder)
C0745136|Hypertensive emergency
C0919726|Postoperative hypertension
C0919726|Postoperative hypertension (disorder)
C0155583|Benign essential hypertension (disorder)
C0155583|benign essential hypertension (diagnosis)
C0155583|benign essential hypertension
C0155583|Benign hypertension
C0155583|Essential hypertension, benign
C0333301|Hypertensive ischemic ulcer -RETIRED-
C0333301|Hypertensive ischaemic ulcer -RETIRED-
C0333301|Hypertensive ischemic ulcer
C0333301|Hypertensive ischaemic ulcer
C0333301|Hypertensive ischemic ulcer (disorder)
C0333301|Ulcer of skin caused by ischemia due to hypertension
C0333301|Ulcer of skin caused by ischaemia due to hypertension
C0333301|Ulcer of skin caused by ischaemia due to hypertensive disease
C0333301|Ulcer of skin caused by ischemia due to hypertensive disease (disorder)
C0333301|Ulcer of skin caused by ischemia due to hypertensive disease
C0333301|ulcer of skin caused by ischemia due to hypertensive disease. dl (disorder)
C0392682|Elevated blood-pressure reading, without diagnosis of hypertension
C0392682|Increased blood pressure (not hypertension)
C0392682|Elevated blood pressure reading without diagnosis of hypertension
C0392682|Elevated blood-pressure reading without diagnosis of hypertension (finding)
C0392682|Elevated blood pressure reading without diagnosis of hypertension (situation)
C0392682|Elev bl pres w/o hypertn
C0392682|Elevated blood-pressure reading, w/o diagnosis of htn
C0392682|elevated blood pressure reading without diagnosis of hypertension (physical finding)
C0392682|Elevated blood-pressure reading w/out diagn of hypertension (disorder)
C0392682|Elevated blood-pressure reading w/out diagn of hypertension
C0392682|Elevated blood-pressure reading without diagnosis of hypertension
C0392682|blood pressure; high, incidental reading, without diagnosis of hypertension
C0392682|increased; blood pressure, reading, no diagnosis of hypertension
C0392682|Elevated blood pressure (not hypertension)
C0392682|Elevated blood-pressure reading without diagnosis of hypertension (disorder)
C0476453|[D]Raised blood pressure reading (context-dependent category)
C0476453|[D]Raised blood pressure reading (situation)
C0476453|Raised blood pressure reading (disorder)
C0476453|[D]Raised blood pressure reading
C0476453|Raised blood pressure reading
C0340272|Other specified hypertensive disease
C0340272|Other specified hypertensive disease (disorder)
C0497247|Elevated blood pressure
C0497247|Raised blood pressure
C0497247|Increased blood pressure
C0497247|Increase in blood pressure
C0497247|Blood pressure increased
C0497247|Blood pressure elevation
C0497247|Raised blood pressure (finding)
C0497247|Finding of increased blood pressure
C0497247|Elevated BP
C0497247|Rise in blood pressure
C0497247|Pressure blood increased
C0497247|Blood pressure raised
C0497247|Pressure arterial increased
C0497247|Arterial pressure high
C0497247|Rise in BP
C0497247|Arterial pressure NOS increased
C0497247|BP raised
C0497247|Raised BP
C0497247|Finding of increased blood pressure (finding)
C0497247|blood pressure; increased
C0497247|increased; blood pressure
C2887335|Postprocedural hypertension
C2887335|hypertension iatrogenic postprocedural
C2887335|postprocedural hypertension (diagnosis)
C3661921|Perioperative hypertension
C3661921|Perioperative hypertension (disorder)
C3665418|Labile hypertension
C3665418|labile hypertension (physical finding)
C3665418|labile hypertension was observed
C3665418|Hypertension;labile
C3665418|labile hypertension (diagnosis)
C3665418|Labile hypertension (disorder)
C3665418|White coat hypertension
C1301626|Hypertension with albuminuria
C1301626|Hypertension with albuminuria (diagnosis)
C1301626|Hypertension with albuminuria (disorder)
C0264637|Benign hypertension (disorder)
C0264637|Hypertension;benign
C0264637|benign hypertension
C0264637|benign hypertension (diagnosis)
C0264637|benign; hypertension
C0264637|hypertension; benign
C0235222|Diastolic hypertension
C0235222|diastolic hypertension (diagnosis)
C0235222|hypertenion diastolic
C0235222|Hypertension diastolic
C0235222|Diastolic hypertension (disorder)
C0235222|Diastolic hypertension, NOS
C0520539|Hypertensive episode
C0520539|hypertensive episode (diagnosis)
C0520539|Hypertensive episodes
C0520539|Hypertensive episode (disorder)
C1997276|Exertional hypertension
C1997276|Exertional hypertension (disorder)
C1997276|exertional hypertension (diagnosis)
C0221155|Systolic hypertension
C0221155|Systolic hypertension (disorder)
C0221155|systolic hypertension (diagnosis)
C0221155|hypertension systolic
C0520540|rebound hypertension (diagnosis)
C0520540|Rebound hypertension
C0520540|Hypertension rebound
C0520540|Rebound hypertension (disorder)
C0152170|Transient hypertension
C0152170|transient hypertension (diagnosis)
C0152170|Transient hypertension (disorder)
C3669043|Intermittent hypertension (disorder)
C3669043|Intermittent hypertension
C1862170|HYPERTENSION WITH BRACHYDACTYLY
C1862170|Bilginturan syndrome
C1862170|Brachydactyly type E with short stature and hypertension
C1862170|Brachydactyly with hypertension
C1862170|Brachydactyly, Type E, With Short Stature And Hypertension
C1862170|HTNB
C1837739|HYPERTENSION, DIASTOLIC, RESISTANCE TO
C1839021|HYPOMAGNESEMIA, HYPERTENSION, AND HYPERCHOLESTEROLEMIA, MITOCHONDRIAL
C1839021|HYPERTENSION, HYPERCHOLESTEROLEMIA, AND HYPOMAGNESEMIA, MITOCHONDRIAL
C1833688|OSTEOCHONDRODYSPLASIA, RHIZOMELIC, WITH CALLOSAL AGENESIS, THROMBOCYTOPENIA, HYDROCEPHALUS, AND HYPERTENSION
C3501739|Tachycardia, Hypertension, Microphthalmia, And Hyperglycinuria
C1854631|HYPERTENSION, EARLY-ONSET, AUTOSOMAL DOMINANT, WITH SEVERE EXACERBATION IN PREGNANCY
C1834155|HYPERTENSION, RESISTANT TO CONVENTIONAL THERAPY
C1834155|HYPERTENSION RESISTANT TO CONVENTIONAL THERAPY
C1865267|ARTERIAL OCCLUSIVE DISEASE, PROGRESSIVE, WITH HYPERTENSION, HEART DEFECTS, BONE FRAGILITY, AND BRACHYSYNDACTYLY
C1865267|Grange Occlusive Arterial Syndrome
C3831106|Chronic Maternal Hypertension with Superimposed Preeclampsia
C3827254|Chronic Maternal Hypertension
C3837203|hypertension (systemic) susceptibility
C3837203|hypertension (systemic) susceptibility (diagnosis)
C3874846|Hypertension in chronic kidney disease due to type 2 diabetes mellitus (disorder)
C3874846|Hypertension in chronic kidney disease due to type II diabetes mellitus
C3874846|Hypertension in chronic kidney disease due to type 2 diabetes mellitus
C3874779|Hypertension in chronic kidney disease due to type 1 diabetes mellitus (disorder)
C3874779|Hypertension in chronic kidney disease due to type I diabetes mellitus
C3874779|Hypertension in chronic kidney disease due to type 1 diabetes mellitus
C0020546|Hypertensive crisis
C0020546|Hypertensive crisis (disorder)
C0020546|Crisis hypertensive
C2902961|Page kidney
C2902961|page kidney (diagnosis)
C2902961|Hypertension due to compression of renal parenchyma
C2902961|Hypertension due to compression of renal parenchyma (disorder)
C1857175|Hypertension, episodic
C1857175|Episodic hypertension
C4025693|Hypertension associated with pheochromocytoma
C0020545|Hypertension, Renovascular
C0020545|Renovascular Hypertension
C0020545|renovascular hypertension (diagnosis)
C0020545|secondary hypertension renovascular
C0020545|Hypertension, Renovascular [Disease/Finding]
C0020545|Secondary renovascular hypertension NOS
C0020545|Secondary renovascular hypertension NOS (disorder)
C0020545|Hypertension due to renal artery hyperplasia
C0020545|Hypertension due to renovascular disease
C0020545|Renovascular hypertension (disorder)
C0020545|hypertension; renovascular disorders
C0020545|hypertension; renovascular
C0020545|renal disease; hypertension, arterial
C0020545|renovascular; hypertension
C1840375|Elevated diastolic blood pressure
C1840376|Elevated mean arterial pressure
C1840374|Elevated systolic blood pressure
C4076686|Supine hypertension
C4076686|Supine hypertension (disorder)
C0151620|Hypertensive encephalopathy
C0151620|HYPERTENSIVE ENCEPH
C0151620|ENCEPH HYPERTENSIVE
C0151620|hypertensive encephalopathy (diagnosis)
C0151620|Hypertens encephalopathy
C0151620|Encephalopathy, Hypertensive
C0151620|Hypertensive Encephalopathy [Disease/Finding]
C0151620|Hypertensive encephalopathy (disorder)
C0151620|Encephalopathy hypertensive
C0151620|encephalopathy; hypertensive
C0494575|Hypertensive heart and renal disease, unspecified, with congestive heart failure
C0494575|Hypertensive heart and renal disease with (congestive) heart failure
C0494575|Hypertensive heart and renal disease with (congestive) heart failure (disorder)
C0494575|failure; cardiorenal, hypertensive, with heart failure
C0264650|Unspecified hypertensive heart disease with congestive heart failure
C0264650|Hypertensive heart disease with (congestive) heart failure
C0264650|Hypertensive heart disease NOS with congestive cardiac failure (disorder)
C0264650|Hypertensive heart disease NOS with congestive cardiac failure
C0264650|Hypertensive heart disease with congestive heart failure
C0264650|hypertensive heart dis with congestive heart failure
C0264650|hypertensive heart dis with congestive heart failure (diagnosis)
C0264650|Hypertensive heart disease with congestive heart failure (disorder)
C0494574|Hypertensive renal disease without renal failure
C0494574|Hy kid NOS w cr kid I-IV
C0494574|Hypertensive renal disease, unspecified, without mention of renal failure
C0494574|Hypertensive chronic kidney disease, unspecified, with chronic kidney disease stage I through stage IV, or unspecified
C0348586|Other unspecified secondary hypertension
C0348586|Other secondary hypertension
C0348586|Second hypertension NEC
C0348586|[X]Other secondary hypertension
C0348586|[X]Other secondary hypertension (disorder)
C0155591|Hypertensive heart disease without (congestive) heart failure
C0155591|Hypertensive heart disease NOS without congestive cardiac failure
C0155591|Hypertensive heart disease NOS without congestive cardiac failure (disorder)
C0155591|Hypertensive heart disease without congestive heart failure
C0155591|Hypertensive heart disease without congestive heart failure (diagnosis)
C0155591|Unspecified hypertensive heart disease without congestive heart failure
C0155591|Hypertensive heart disease without congestive heart failure (disorder)
C0155620|Secondary benign hypertension
C0155620|benign secondary hypertension (diagnosis)
C0155620|benign secondary hypertension
C0155620|secondary hypertension benign
C0155620|Secondary benign hypertension NOS
C0155620|Secondary benign hypertension NOS (disorder)
C0155620|Benign secondary hypertension (disorder)
C0155620|Secondary hypertension, benign
C0155620|Secondary benign hypertension (disorder)
C0544618|Orthostatic hypertension
C0262395|Borderline hypertension
C0262395|borderline; hypertension
C0262395|hypertension; borderline
C1171328|catecholamine hypertension
C0597290|prostaglandin hypertension
C0155622|Other benign secondary hypertension
C0155622|Benign second hypert NEC
C0221154|paroxysmal hypertension (physical finding)
C0221154|paroxysmal hypertension
C0221154|paroxysmal hypertension was observed
C0221154|Hypertension paroxysmal
C0221154|Paroxysmal hypertension (disorder)
C0341909|Hypertension complicating pregnancy, childbirth, and the puerperium
C0341909|Unspecified hypertension complicating pregnancy, childbirth and the puerperium NOS
C0341909|Unspecified hypertension complicating pregnancy, childbirth and the puerperium unspecified (disorder)
C0341909|Unspecified hypertension complicating pregnancy, childbirth and the puerperium unspecified
C0341909|Unspecified hypertension complicating pregnancy, childbirth and the puerperium (disorder)
C0341909|Unspecified hypertension complicating pregnancy, childbirth and the puerperium NOS (disorder)
C0341909|Unspecified hypertension complicating pregnancy, childbirth and the puerperium
C0341909|Hypertension complicating pregnancy; childbirth and the puerperium
C0341909|Hypertension complicating pregnancy, childbirth and the puerperium
C0341909|Hypertension complicating pregnancy, childbirth and the puerperium (disorder)
C1443005|Non-proteinuric hypertension of pregnancy (disorder)
C1443005|Hypertension in the obstetric context
C1443005|Hypertension in the obstetric context (disorder)
C1443005|Non-proteinuric hypertension of pregnancy
C1443005|Hypertension without albuminuria AND without oedema in the obstetric context
C1443005|Hypertension without albuminuria AND without edema in the obstetric context
C1443005|Hypertension in the obstetric context, NOS
C1443005|Hypertension without albuminuria or edema in the obstetric context, NOS
C1443005|Hypertension in the obstetric context (disorder) [Ambiguous]
C1443005|Non-proteinuric hypertension of pregnancy [Ambiguous]
C1171326|bradykinin hypertension
C1171351|kinin hypertension
C0349368|Hypertension secondary to endocrine disorders
C0349368|hypertension secondary to endocrine disorders (diagnosis)
C0349368|secondary hypertension to endocrine disorders
C0349368|hypertension; secondary, due to endocrine disorders
C0349368|secondary; hypertension, due to endocrine disorders
C0349368|Hypertension secondary to endocrine disorder (disorder)
C0349368|Hypertension secondary to endocrine disorder
C0349368|Hypertension secondary to endocrine disorders (disorder)
C0348587|Hypertension secondary to other renal disorders
C0348587|[X]Hypertension secondary to other renal disorders (disorder)
C0348587|[X]Hypertension secondary to other renal disorders
C0348587|hypertension; secondary, due to renal disorders
C0348587|secondary; hypertension, due to renal disorders
C0348860|Hypertensive renal disease, unspecified, with renal failure
C0348860|Hypertensive renal disease with renal failure
C0348860|Hyp kid NOS w cr kid V
C0348860|Hypertensive chronic kidney disease, unspecified, with chronic kidney disease stage V or end stage renal disease
C0348860|hypertensive kidney disease with renal failure (diagnosis)
C0348860|hypertensive kidney disease with renal failure
C0348860|Hypertensive renal disease with renal failure (disorder)
C0348860|hypertension; renal disease, hypertensive, with renal failure
C0348860|insufficiency; renal, chronic, hypertensive
C0348860|insufficiency; renal, with hypertension
C0348860|kidney; hypertension, with renal failure
C0348879|Hypertensive heart and renal disease, unspecified, with renal failure
C0348879|Hypertensive heart and renal disease with renal failure
C0348879|hypertensive heart and renal disease with renal failure (diagnosis)
C0348879|hypertensive heart and chronic kidney disease with renal failure
C0348879|Hy ht/kd NOS st V w/o hf
C0348879|Hypertensive heart and chronic kidney disease, unspecified, without heart failure and with chronic kidney disease stage V or end stage renal disease
C0348879|Hypertensive heart and renal disease with renal failure (disorder)
C0348879|failure; cardiorenal, hypertensive, with renal failure
C0348879|insufficiency; renal, with hypertensive heart disease
C0348879|kidney; insufficiency, with hypertensive heart disease
C0494576|Hypertensive heart and renal disease, unspecified, with congestive heart failure and renal failure
C0494576|Hypertensive heart and renal disease with both (congestive) heart failure and renal failure
C0494576|Hyp ht/kd NOS st V w hf
C0494576|Hypertensive heart and chronic kidney disease, unspecified, with heart failure and chronic kidney disease stage V or end stage renal disease
C0494576|Hypertensive heart and renal disease, unspecified, with heart failure and renal failure
C0494576|Hypertensive heart and renal disease with both (congestive) heart failure and renal failure (disorder)
C0494576|insufficiency; renal, with hypertensive heart disease and heart failure
C0494576|kidney; insufficiency, with hypertensive heart disease and heart failure
C0452204|Neonatal hypertension
C0452204|Hypertension neonatal
C0452204|neonatal hypertension (diagnosis)
C0452204|Hypertension, neonatal
C0452204|Neonatal hypertension (disorder)
C0452204|hypertension; neonatal
C0452204|hypertension; newborn
C0452204|neonatal; hypertension
C0452204|newborn; hypertension
C0269660|Eclampsia added to pre-existing hypertension
C0269660|Eclampsia added to pre-existing hypertension (disorder)
C0156689|Hypertens NOS-antepartum
C0156689|Unspecified hypertension complicating pregnancy, childbirth, or the puerperium, antepartum condition or complication
C0156689|Unspecified antepartum hypertension
C0497248|Hypertension;uncomplicated
C0497248|Uncomplicated hypertension
C1335457|Postpartum Hypertension
C0028840|Hypertensions, Ocular
C0028840|Ocular Hypertension
C0028840|Ocular Hypertensions
C0028840|preglaucoma ocular hypertension (diagnosis)
C0028840|preglaucoma ocular hypertension
C0028840|Hypertension, Ocular
C0028840|Ocular Hypertension [Disease/Finding]
C0028840|Hypertension ocular
C0028840|Pressure Behind Eyeballs
C0028840|OH - Ocular hypertension
C0028840|OHT - Ocular hypertension
C0028840|Ocular hypertension (disorder)
C0028840|hypertension; ocular
C0028840|ocular; hypertension
C2227904|American College of Physicians (ACP) staging stage 1 hypertension: 140-159/90-99 (physical finding)
C2227904|American College of Physicians (ACP) staging stage 1 hypertension: 140-159/90-99
C2227904|ACP staging stage 1 hypertension: 140-159 / 90-99
C2227905|American College of Physicians (ACP) staging stage 2 hypertension: greater than equal to 160/100
C2227905|American College of Physicians (ACP) staging stage 2 hypertension: greater than equal to 160/100 (physical finding)
C2227905|ACP staging stage 2 hypertension: greater than or = 160/100
C2216285|elevation of both systolic and diastolic blood pressures (physical finding)
C2216285|elevation of both systolic and diastolic BP
C2216285|combined systolic and diastolic elevation
C2216285|elevation of both systolic and diastolic blood pressures
C2216285|combined systolic and diastolic elevation was observed
C0341934|Transient hypertension of pregnancy
C0341934|TRANSIENT HYPERTENSION PREGN
C0341934|pregnancy complicated by transient hypertension (diagnosis)
C0341934|pregnancy complicated by transient hypertension
C0341934|Transient hypertension of pregnancy (disorder)
C0341934|Transient hypertension of pregnancy NOS (disorder)
C0341934|Transient hypertension of pregnancy unspecified (disorder)
C0341934|Transient hypertension of pregnancy unspecified
C0341934|Transient hypertension of pregnancy NOS
C0341934|Transient Hypertension, Pregnancy
C0341934|pregnancy; hypertension, transient
C0341934|Transient hypertension of pregnancy (disorder) [Ambiguous]
C0341934|Hypertension, Pregnancy Transient
C0341934|Pregnancy Transient Hypertension
C1556272|CTCAE Grade 1 Hypertension
C1556272|Grade 1 Hypertension
C1556275|CTCAE Grade 4 Hypertension
C1556275|Grade 4 Hypertension
C1556276|CTCAE Grade 5 Hypertension
C1556276|Grade 5 Hypertension
C1556274|CTCAE Grade 3 Hypertension
C1556274|Grade 3 Hypertension
C1556273|CTCAE Grade 2 Hypertension
C1556273|Grade 2 Hypertension
