C0019151|Hepatic Encephalopathy
C3266165|Hepatic encephalopathy in fulminant hepatic failure
C2729507|hepatic encephalopathy with coma
C3888788|Minimal hepatic encephalopathy
C4024937|Chronic hepatic encephalopathy
C3889995|CDISC SDTM West Haven Hepatic Encephalopathy Grade Terminology
C3890564|West Haven Hepatic Encephalopathy Grade
C4086961|West Haven Criteria - West Haven Hepatic Encephalopathy Grade
C3151062|INFECTIONS, RECURRENT, WITH ENCEPHALOPATHY, HEPATIC DYSFUNCTION, AND CARDIOVASCULAR MALFORMATIONS
C3889290|West Haven Hepatic Encephalopathy Grade 3
C3889292|West Haven Hepatic Encephalopathy Grade 1
C3889293|West Haven Hepatic Encephalopathy Grade 4
C3889824|West Haven Hepatic Encephalopathy Grade 2
C3890401|West Haven Hepatic Encephalopathy Grade 0
C4016797|INFECTIONS, RECURRENT, ASSOCIATED WITH ENCEPHALOPATHY, HEPATIC DYSFUNCTION, AND CARDIOVASCULAR MALFORMATIONS
C4086072|CDISC Clinical Classification West Haven Criteria Test Code Terminology
C4086073|CDISC Clinical Classification West Haven Criteria Test Name Terminology
C3854121|Documentation of medical reason(s) for not receiving annual screening for hcv infection (e.g., decompensated cirrhosis indicating advanced disease [i.e., ascites, esophageal variceal bleeding, hepatic encephalopathy], hepatocellular carcinoma, waitlist for organ transplant, limited life expectancy, other medical reasons)
C3871346|Documentation of medical reason(s) for not receiving one-time screening for hcv infection (e.g., decompensated cirrhosis indicating advanced disease [ie, ascites, esophageal variceal bleeding, hepatic encephalopathy], hepatocellular carcinoma, waitlist for organ transplant, limited life expectancy, other medical reasons)
C0019151|Encephalopathies, Hepatic
C0019151|Encephalopathies, Portosystemic
C0019151|Hepatic Encephalopathies
C0019151|Hepatic Encephalopathy
C0019151|Portosystemic Encephalopathies
C0019151|ENCEPH HEPATOCEREBRAL
C0019151|ENCEPH PORTAL SYSTEMIC
C0019151|HEPATIC ENCEPH
C0019151|PORTOSYSTEMIC ENCEPH
C0019151|ENCEPH PORTOSYSTEMIC
C0019151|PORTAL SYSTEMIC ENCEPH
C0019151|HEPATOCEREBRAL ENCEPH
C0019151|ENCEPH HEPATIC
C0019151|hepatic encephalopathy (diagnosis)
C0019151|Hepatocerebral encephalopathy -RETIRED-
C0019151|Encephalopathies, Hepatocerebral
C0019151|Hepatocerebral Encephalopathies
C0019151|Encephalopathies, Portal-Systemic
C0019151|Portal Systemic Encephalopathy
C0019151|Portal-Systemic Encephalopathies
C0019151|hepatic encephalopathy NOS
C0019151|Portosystemic Encephalopathy
C0019151|Encephalopathy, Hepatocerebral
C0019151|Hepatocerebral Encephalopathy
C0019151|Hepatic Encephalopathy [Disease/Finding]
C0019151|Portal-Systemic Encephalopathy
C0019151|Encephalopathy, Hepatic
C0019151|Encephalopathy, Portal-Systemic
C0019151|Encephalopathy, Portosystemic
C0019151|hepatic coma/encephalopathy
C0019151|Encephalopathy, Portal Systemic
C0019151|Gaustad's syndrome
C0019151|Portal systemic encephalopathy (disorder)
C0019151|Transient hepatargy syndrome
C0019151|Encephalopathy - hepatic
C0019151|Hepatocerebral encephalopathy (disorder)
C0019151|Encephalopathy hepatic
C0019151|HE - Hepatic encephalopathy
C0019151|Hepatic encephalopathy (disorder)
C0019151|encephalopathy; hepatic
C0019151|encephalopathy; portosystemic
C0019151|hepatic; encephalopathy
C0019151|portosystemic; encephalopathy
C2729507|hepatic encephalopathy with coma (diagnosis)
C2729507|hepatic encephalopathy with coma
C0019147|Comas, Hepatic
C0019147|Hepatic Comas
C0019147|Coma, Hepatic
C0019147|Hepatic coma
C0019147|Coma hepatic
C0019147|Hepatic coma NOS
C0019147|Coma;hepatic
C0019147|Hepatic coma (disorder)
C0019147|Hepatocerebral intoxication
C0019147|coma; hepatic
C0019147|hepatic; coma
C3266165|Hepatic encephalopathy in fulminant hepatic failure
C3266165|Hepatic encephalopathy in fulminant hepatic failure (disorder)
C0751198|Hepatic Stupors
C0751198|Stupor, Hepatic
C0751198|Stupors, Hepatic
C0751198|Hepatic Stupor
C1836797|COXPD1
C1836797|COMBINED OXIDATIVE PHOSPHORYLATION DEFICIENCY 1
C1836797|Hepatoencephalopathy, Early Fatal Progressive
C4024937|Chronic hepatic encephalopathy
C3888788|Minimal hepatic encephalopathy
C3889824|West Haven Hepatic Encephalopathy Grade 2
C3889824|GRADE 2
C3890401|GRADE 0
C3890401|West Haven Hepatic Encephalopathy Grade 0
C3889292|GRADE 1
C3889292|West Haven Hepatic Encephalopathy Grade 1
C3889290|GRADE 3
C3889290|West Haven Hepatic Encephalopathy Grade 3
C3889293|West Haven Hepatic Encephalopathy Grade 4
C3889293|GRADE 4
C3854121|Documentation of medical reason(s) for not receiving annual screening for hcv infection (e.g., decompensated cirrhosis indicating advanced disease [i.e., ascites, esophageal variceal bleeding, hepatic encephalopathy], hepatocellular carcinoma, waitlist for organ transplant, limited life expectancy, other medical reasons)
C3854121|Doc med reas no ann srn hcv
C3871346|Documentation of medical reason(s) for not receiving one-time screening for hcv infection (e.g., decompensated cirrhosis indicating advanced disease [ie, ascites, esophageal variceal bleeding, hepatic encephalopathy], hepatocellular carcinoma, waitlist for organ transplant, limited life expectancy, other medical reasons)
C3871346|Doc med reas no scrn hcv
