C0015879|Ferritin
C0373607|Ferritin measurement
C0003590|Ferritins, apo-
C0003590|Apoferritins
C0003590|Apoferritins [Chemical/Ingredient]
C0003590|Apoferritin
C0015879|Ferritin
C0015879|Ferritins
C0015879|ferritin (medication)
C0015879|hematinics ferritin
C0015879|Ferritins [Chemical/Ingredient]
C0015879|Ferritin (substance)
C2607715|ferritin A, E coli
C2607715|FtnA protein, E coli
C2607715|EcFtnA protein, E coli
C1987810|Ferritin &#x7C; bld-ser-plas
C1987811|Ferritin &#x7C; Red Blood Cells
C2357527|Ferritin &#x7C; Body Fluid
C3657120|FER1 protein, Arabidopsis
C3657120|At5g01600 protein, Arabidopsis
C3180177|mitochondrial ferritin, human
C3180177|FtMt protein, human
C4077042|AtFer3 protein, Arabidopsis
C4077042|Fer3 protein, Arabidopsis
C4077041|Fer4 protein, Arabidopsis
C4077041|AtFer4 protein, Arabidopsis
C0071525|cationized ferritin
C0071525|polycationic ferritin
C0056922|cytochrome b-1
C0056922|bacterioferritin
C0056922|cytochrome b1
C0060262|ferritin-protein conjugates
C0101243|isoferritin, acidic
C0101243|acidic isoferritin
C0071012|phytoferritin
C0620494|DA-Fe conjugate
C0620494|daunomycin-ferretin conjugate
C0620494|ferretin-daunomycin conjugate
C0621939|fucosyl ferritin
C0051915|anionized ferritin
C0060260|ferritin hydrazide
C0625267|ferritin-peanut agglutinin conjugate
C0625267|peanut-lectin-ferritin conjugate
C0627610|protamine-ferritin conjugate
C0627610|ferritin-protamine
C0119873|ferritin, glycosylated
C0119873|glycosylated ferritin
C0119873|glycosylated ferritins
C0081681|avidin-ferritin biotin
C0630489|ferritin-Con A conjugate
C0630489|concanavalin A-ferritin conjugate
C0630489|ferritin-concanavalin A conjugate
C0631398|ferritin-wheat germ agglutinin
C0631398|wheat germ agglutinin-ferritin
C0636154|phytosiderin
C0649838|CHA-ferritin
C0649838|ferritin-cyclohexyladenosine
C0166450|heme ferritin
C0166450|hemoferritin
C0166450|haemoferritin
C0963515|cold shock protein, Listeria
C0963515|ferritin-like protein, Listeria
C0963515|18-kDa CSP protein, Listeria
C0968127|ferritin pfr, Helicobacter pylori
C0968127|pfr protein, Helicobacter pylori
C1448299|HuHF protein, human
C1448299|FTH1 protein, human
C1448299|PLIF protein, human
C1448299|ferritin, heavy polypeptide 1, human
C1448299|placenta immunoregulatory factor, human
C1448299|placental immunomodulatory ferritin protein, human
C1504956|PLIF protein, mouse
C1504956|placental immunomodulatory ferritin protein, mouse
C0105254|Basic Isoferritin
C0105254|Isoferritin, Basic
C0063967|Isoferritin
C0373607|Ferritin
C0373607|Ferritin measurement
C0373607|Test;ferritin
C0373607|ASSAY OF FERRITIN
C0373607|Ferritin (blood protein) level
C0373607|Measurement of ferritin
C0373607|Ferritin level
C0373607|Ferritin measurement (procedure)
C0373607|ferritin test
C1276043|Plasma ferritin level
C1276043|Plasma ferritin measurement (procedure)
C1276043|Plasma ferritin measurement
C0696113|Serum ferritin
C0696113|serum ferritin level (lab test)
C0696113|serum ferritin level
C0696113|Serum ferritin level (procedure)
C0696113|Ferritin - serum
C0696113|Serum ferritin measurement (procedure)
C0696113|Serum ferritin measurement
C0696113|Serum ferritin each test
C0696113|serum ferritin ea.tst
C0565897|Serum ferritin/TIBC measurement (procedure)
C0565897|Serum ferritin/Total iron binding capacity measurement
C0565897|Serum ferritin/Total iron binding capacity measurement (procedure)
C0565897|Serum ferritin/TIBC
C0565897|Serum ferritin/TIBC measurement
