C0338831|Manic
C0564408|Manic mood
C0241934|Hypomania
C0154436|atypical manic disorder
C0154436|atypical manic disorder (diagnosis)
C0154436|Atypical manic disorder (disorder)
C0338831|Mania
C0338831|Manias
C0338831|Manic States
C0338831|State, Manic
C0338831|States, Manic
C0338831|Manic
C0338831|Manic State
C0338831|Mania NOS
C0338831|Mania (disorder)
C0349208|Manic episode, unspecified
C0349208|Manic episode
C0349208|manic episode (diagnosis)
C0349208|[X]Mania NOS
C0349208|[X]Manic episode, unspecified
C0349208|[X]Manic episode
C0349208|[X] Mania: [episode, unspecified] or [NOS]
C0349208|[X]Manic episode, unspecified (disorder)
C0349208|[X] Mania: [episode, unspecified] or [NOS] (disorder)
C0349208|episode; manic
C0349208|manic; episode
C0005586|Bipolar Disorders
C0005586|MANIC DEPRESSIVE ILLNESS
C0005586|Bipolar Affective Psychosis
C0005586|Bipolar Disorder
C0005586|Manic Depressive Psychosis
C0005586|Manic-Depressive Psychoses
C0005586|Psychoses, Bipolar Affective
C0005586|Psychoses, Manic Depressive
C0005586|Psychosis, Bipolar Affective
C0005586|Psychosis, Manic Depressive
C0005586|Bipolar affective disorder
C0005586|Disorder, Bipolar
C0005586|Manic-depressive psychosis
C0005586|Bipolar affective disorder, unspecified
C0005586|BIPOLAR DIS
C0005586|Manic-Depression
C0005586|manic depressive disorder
C0005586|BPAD
C0005586|unspecified bipolar disorder
C0005586|unspecified bipolar disorder (diagnosis)
C0005586|bipolar disorder not otherwise specified
C0005586|Manic depressive
C0005586|Bipolar disorder NOS
C0005586|manic-depressive reaction
C0005586|manic-depressive illness
C0005586|Bipolar disorder, unspecified
C0005586|Affective Psychosis, Bipolar
C0005586|Bipolar Disorder [Disease/Finding]
C0005586|Psychoses, Manic-Depressive
C0005586|Psychosis, Manic-Depressive
C0005586|Disorder;bipolar
C0005586|Depression;manic
C0005586|Psychosis;manic depressive
C0005586|Bi-polar Disorder
C0005586|Bipolar disorder (disorder)
C0005586|Unspecified bipolar affective disorder
C0005586|Depressive-manic psych.
C0005586|Unspecified bipolar affective disorder (disorder)
C0005586|Unspecified bipolar affective disorder, unspecified
C0005586|[X]Bipolar affective disorder, unspecified
C0005586|[X]Bipolar affective disorder, unspecified (disorder)
C0005586|Unspecified bipolar affective disorder, unspecified (disorder)
C0005586|Unspecified bipolar affective disorder, NOS
C0005586|Manic-depress.psychoses
C0005586|Unspecified bipolar affective disorder, NOS (disorder)
C0005586|Manic depression
C0005586|Manic depressive reaction
C0005586|Reaction manic-depressive
C0005586|Psychosis manic-depressive
C0005586|MDI - Manic-depressive illness
C0005586|bipolar; disorder, affective
C0005586|bipolar; disorder
C0005586|disorder; bipolar, affective
C0005586|disorder; bipolar
C0005586|manic-depressive; disorder
C0005586|manic-depressive; psychosis
C0005586|manic-depressive; syndrome
C0005586|psychosis; manic-depressive
C0005586|syndrome; manic-depressive
C0005586|Bipolar disorder, NOS
C0005586|Bipolar Mood Disorder
C0005586|Manic-depressive reaction NOS
C0005586|Manic-depressive syndrome NOS
C0236756|Manic disorder, single episode, unspecified degree
C0236756|bipolar I disorder with single manic episode (diagnosis)
C0236756|bipolar I disorder with single manic episode
C0236756|Bipol I single manic NOS
C0236756|Bipolar I disorder, single manic episode, unspecified
C0236756|Bipolar 1 disorder, single manic episode
C0236756|Manic disorder, single episode NOS (disorder)
C0236756|Manic disorder, single episode
C0236756|Manic disorder, single episode NOS
C0236756|Single manic episode, unspecified
C0236756|Single manic episode, unspecified (disorder)
C0236756|Manic disorder, single episode (diagnosis)
C0236756|manic episode single
C0236756|Bipolar I disorder, single manic episode
C0236756|Manic disorder, single episode (disorder)
C0236756|Bipolar I disorder, single manic episode (disorder)
C0338846|Manic stupor
C0338846|Manic stupor (diagnosis)
C0338846|manic episode stupor
C0338846|Manic stupor (disorder)
C0338846|manic; stupor
C0338846|stupor; manic
C0338832|manic disorder with recurrent episode
C0338832|manic disorder, recurrent episode
C0338832|manic disorder with recurrent episode (diagnosis)
C0338832|Recurrent manic episodes NOS
C0338832|Recurrent manic episode NOS (disorder)
C0338832|Recurrent manic episodes, unspecified (disorder)
C0338832|[X]Recurrent manic episodes
C0338832|Recurrent manic episode NOS
C0338832|Recurrent manic episodes, unspecified
C0338832|Recurrent manic episodes
C0338832|Recurrent manic episodes (disorder)
C0270601|AMOK
C0270601|manic episode amok
C0270601|Amok (diagnosis)
C0270601|Cafard
C0270601|Cathard
C0270601|Iich'aa
C0270601|Mal de pelea
C0270601|Amok (disorder)
C0270601|Amuck
C0241934|Hypomania
C0241934|Hypomania (disorder)
C0241934|Hypomania (diagnosis)
C0241934|manic episode hypomania
C0241934|Hypomanic Mood
C0241934|Hypomanic mood (finding)
C0865308|Mania NOS single episode or unspecified
C0865309|Monopolar mania NOS single episode or unspecified
C2874863|Manic episode without psychotic symptoms
C2874863|Manic episode without psychotic symptoms, unspecified
C2874863|manic episode without psychotic symptoms (diagnosis)
C0564408|Manic mood
C0564408|Manic
C0564408|Manic mood (finding)
C0865305|Hypomania NOS single episode or unspecified
C0865306|Mild hypomania NOS single episode or unspecified
C0865307|Hypomanic psychosis single episode or unspecified
C1389907|bipolar; disorder, single manic episode, mild
C1389907|disorder; bipolar, single manic episode, mild
C1396834|episode; hypomanic
C1396834|hypomanic; episode
C1400223|excitement; hypomanic
C1400223|hypomanic; excitement
C0683410|Hypomanic psychoses
C0683410|Hypomanic psychosis
C0683410|hypomanic; psychosis
C0683410|psychosis; hypomanic
C1400224|hypomanic; reaction
C1400224|reaction; hypomanic
