C0004002|Aspartate Transaminase
C0201899|Aspartate aminotransferase measurement
C0684153|GLUTAMATE OXALOACETATE TRANS 002
C0684153|Aspartate Aminotransferase, Mitochondrial [Chemical/Ingredient]
C0684153|Glutamate Oxaloacetate Transaminase-2
C0684153|Aspartate Aminotransferase, Mitochondrial
C0684153|Aminotransferase, Mitochondrial Aspartate
C0684153|Glutamate Oxaloacetate Transaminase 2
C0684153|Mitochondrial Aspartate Aminotransferase
C0684153|Oxaloacetate Transaminase-2, Glutamate
C0684153|Transaminase-2, Glutamate Oxaloacetate
C0684153|Plasma Membrane-Associated Fatty Acid-Binding Protein
C0684153|EC 2.6.1.1
C0684153|Aspartate Aminotransferase 2
C0684153|mAspAT
C0684153|FABP-1
C0684153|FABPpm
C0684153|Fatty Acid-Binding Protein
C0684153|Transaminase A
C0684153|GOT2
C0684153|Mitochondrial Glutamic-Oxaloacetic Transaminase 2
C0949643|GLUTAMATE OXALOACETATE TRANS 001
C0949643|Aspartate Aminotransferase, Cytoplasmic
C0949643|Aspartate Aminotransferase, Cytoplasmic [Chemical/Ingredient]
C0949643|Glutamate Oxaloacetate-Transaminase-1
C0949643|Aminotransferase, Cytoplasmic Aspartate
C0949643|Cytoplasmic Aspartate Aminotransferase
C0949643|Oxaloacetate-Transaminase-1, Glutamate
C0949643|Aspartate Aminotransferase 1
C0949643|EC 2.6.1.1
C0949643|Glutamate Oxaloacetate Transaminase 1
C0949643|Transaminase A
C0949643|GOT1
C0949643|Glutamate Oxaloacetate Transaminase-1
C0949643|Soluble Glutamic-Oxaloacetic Transaminase 1
C0004002|Aminotransferase, Aspartate
C0004002|Aminotransferase, L-Aspartate-2-Oxoglutarate
C0004002|Apoaminotransferase, Aspartate
C0004002|Aspartate Aminotransferase
C0004002|Aspartate Transaminase
C0004002|Glutamic-Oxaloacetic Transaminase
C0004002|Transaminase, Aspartate
C0004002|Transaminase, Glutamate-Aspartate
C0004002|Transaminase, Glutamic-Oxaloacetic
C0004002|Glutamate Aspartate Transaminase
C0004002|Glutamic Oxaloacetic Transaminase
C0004002|L Aspartate 2 Oxoglutarate Aminotransferase
C0004002|L-Aspartate:2-oxoglutarate aminotransaminase
C0004002|GLUTAMIC OXALOACETIC TRANS 000
C0004002|transaminase A
C0004002|glutamic aspartic transaminase
C0004002|Aspartate Aminotransferases
C0004002|Glutamate-Aspartate Transaminase
C0004002|L-Aspartate-2-Oxoglutarate Aminotransferase
C0004002|Aspartate Apoaminotransferase
C0004002|Aspartate Aminotransferases [Chemical/Ingredient]
C0004002|Aminotransferases, Aspartate
C0004002|ASAT - Aspartate aminotransferase
C0004002|AST - Aspartate transaminase
C0004002|GOT
C0004002|Glutamate oxaloacetate transaminase
C0004002|Glutamic-aspartic transaminase
C0004002|L-aspartate:2-oxoglutarate aminotransferase
C0004002|Aspartate aminotransferase (substance)
C1981807|Aspartate aminotransferase &#x7C; peritoneal fluid
C1981801|Aspartate aminotransferase &#x7C; bld-ser-plas
C1981802|Aspartate aminotransferase &#x7C; body fluid
C1981810|Aspartate aminotransferase &#x7C; red blood cells
C1981806|Aspartate aminotransferase &#x7C; gastric fluid
C1981813|Aspartate aminotransferase &#x7C; urine
C1981814|Aspartate aminotransferase.macromolecular &#x7C; Bld-Ser-Plas
C1981808|Aspartate aminotransferase &#x7C; pleural fluid
C1981812|Aspartate aminotransferase &#x7C; synovial fluid
C1981800|Aspartate aminotransferase &#x7C; amniotic fluid
C1981803|Aspartate aminotransferase &#x7C; cerebral spinal fluid
C1981804|Aspartate aminotransferase &#x7C; dialysis fluid
C1952687|Aspartate aminotransferase.macromolecular
C1952687|Macromolecular aspartate aminotransferase (substance)
C1952687|Macromolecular aspartate aminotransferase
C0201899|serum SGOT
C0201899|serum AST
C0201899|Aspartate aminotransferase
C0201899|GOT
C0201899|AST
C0201899|Aspartate Aminotransferase Measurement
C0201899|Transferase; aspartate amino (AST) (SGOT)
C0201899|TRANSFERASE ASPARTATE AMINO AST SGOT
C0201899|Liver enzyme (SGOT), level
C0201899|Measurement of aspartate amino transferase
C0201899|Measurement of aspartate amino transferase (AST) (SGOT)
C0201899|AST - aspartate transam SGOT (& level) (procedure)
C0201899|AST - aspartate transam SGOT (& level)
C0201899|Transferase (ast) (sgot)
C0201899|SGOT
C0201899|ASPT
C0201899|Aspartate transferase
C0201899|Asp transferase
C0201899|Serum glutamic-oxaloacetic transferase
C0201899|Glutamic-oxaloacetic transferase
C0201899|Serum Aspartate Transaminase Test
C0201899|AST measurement
C0201899|Glutamic oxaloacetic transaminase measurement
C0201899|GOT measurement
C0201899|SGOT measurement
C0201899|Aspartate aminotransferase measurement (procedure)
C1261155|AST serum measurement (procedure)
C1261155|Serum Aspartate Transaminase Measurement
C1261155|Serum Aspartate Aminotransferase Measurement
C1261155|Serum SGOT Measurement
C1261155|AST serum level
C1261155|AST serum level (procedure)
C1261155|Aspartate aminotransferase (AST) serum measurement (procedure)
C1261155|Aspartate aminotransferase serum measurement (procedure)
C1261155|Aspartate aminotransferase (AST) serum measurement
C1261155|Aspartate aminotransferase serum measurement
C1261155|AST serum measurement
C0523517|Aspartate amino transferase/alanine amino transferase ratio measurement
C0523517|Aspartate amino transferase/alanine amino transferase ratio measurement (procedure)
C1278050|Plasma aspartate transaminase level (procedure)
C1278050|Plasma aspartate transaminase level
C1278050|Plasma aspartate transaminase measurement (procedure)
C1278050|Plasma aspartate transaminase measurement
