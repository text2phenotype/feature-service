C0079304|Esophagogastroduodenoscopy
C0009378|colonoscopy
C0079304|Esophagogastroduodenoscopies
C0079304|Esophagogastroduodenoscopy
C0079304|Oesophagogastroduodenoscopy
C0079304|Fibreoptic oesophagogastroduodenoscopy (procedure)
C0079304|Fiberoptic esophagogastroduodenoscopy (procedure)
C0079304|Endoscopy upper gastrointestinal tract
C0079304|EGD
C0079304|Upper GI endoscopy
C0079304|Endoscopic examination of oesophagus, stomach and duodenum
C0079304|Endoscopic examination of esophagus, stomach and duodenum (procedure)
C0079304|Combined upper GI endoscopy
C0079304|OGD - Esophagogastroduodenoscopy
C0079304|OGD - Oesophagogastroduodenoscopy
C0079304|Oesophagogastroduodenoscopy (procedure)
C0079304|Endoscopic examination of upper GI tract
C0079304|Fibreoptic oesophagogastroduodenoscopy
C0079304|Fiberoptic esophagogastroduodenoscopy
C0079304|Endoscopic examination of esophagus, stomach and duodenum
C0079304|Upper Gastrointestinal endoscopy
C0079304|Esophagogastroduodenoscopy Procedures
C0079304|diagnostic esophagogastroduodenoscopy (procedure)
C0079304|diagnostic esophagogastroduodenoscopy
C0079304|esophagogastroduodenoscopy (treatment)
C0079304|Upper gastrointestinal tract endoscopy
C0079304|Esophagogastroduodenoscopy (procedure)
C0472993|Fiberoptic endoscopic snare resection of lesion of esophagus
C0472993|Fibreoptic endoscopic snare resection of lesion of oesophagus
C0472993|Fiberoptic esophagoscopy and snare resection
C0472993|Fibreoptic oesophagoscopy and snare resection
C0472993|Fiberoptic esophagoscopy and snare resection (procedure)
C0472984|Fiberoptic endoscopic laser destruction of lesion of esophagus
C0472984|Fibreoptic endoscopic laser destruction of lesion of oesophagus
C0472984|Fiberoptic esophagoscopy and laser
C0472984|Fibreoptic oesophagoscopy and laser
C0472984|Fiberoptic esophagoscopy and laser (procedure)
C0472981|Fiberoptic endoscopic cauterization of lesion of esophagus
C0472981|Fibreoptic endoscopic cauterisation of lesion of oesophagus
C0472981|Fibreoptic oesophagoscopy and cauterisation
C0472981|Fiberoptic esophagoscopy and cauterization
C0472981|Fiberoptic esophagoscopy and cauterization (procedure)
C0472989|Fiberoptic endoscopic injection sclerotherapy to esophageal varices
C0472989|Fibreoptic endoscopic injection sclerotherapy to oesophageal varices
C0472989|Fiberoptic esophagoscopy and injection sclerotherapy of varices
C0472989|Fibreoptic oesophagoscopy and injection sclerotherapy of varices
C0472989|Fiberoptic esophagoscopy and injection sclerotherapy of varices (procedure)
C0472952|Fiberoptic endoscopic banding of esophageal varices
C0472952|Fibreoptic endoscopic banding of oesophageal varices
C0472952|Fiberoptic esophagoscopy and banding of esophageal varices
C0472952|Fibreoptic oesophagoscopy and banding of oesophageal varices
C0472952|Fiberoptic esophagoscopy and banding of esophageal varices (procedure)
C0472966|Fiberoptic endoscopic removal of foreign body from esophagus
C0472966|Fibreoptic endoscopic removal of foreign body from oesophagus
C0472966|Fiberoptic esophagoscopy and removal of foreign body
C0472966|Fibreoptic oesophagoscopy and removal of foreign body
C0472966|Fiberoptic esophagoscopy and removal of foreign body (procedure)
C0472973|Fiberoptic endoscopic balloon dilation of esophagus
C0472973|Fibreoptic endoscopic balloon dilation of oesophagus
C0472973|Fiberoptic esophagoscopy and balloon dilatation
C0472973|Fibreoptic oesophagoscopy and balloon dilatation
C0472973|Fiberoptic esophagoscopy and balloon dilatation (procedure)
C0472962|Diagnostic fiberoptic endoscopic examination of esophagus and biopsy of lesion of esophagus
C0472962|Diagnostic fibreoptic endoscopic examination of oesophagus and biopsy of lesion of oesophagus
C0472962|Fiberoptic esophagoscopy and biopsy
C0472962|Fibreoptic oesophagoscopy and biopsy
C0472962|Fiberoptic esophagoscopy and biopsy (procedure)
C0472992|Endoscopic snare resection of lesion of esophagus using rigid esophagoscope
C0472992|Endoscopic snare resection of lesion of oesophagus using rigid oesophagoscope
C0472992|Rigid esophagoscopy and snare resection
C0472992|Rigid oesophagoscopy and snare resection
C0472992|Rigid esophagoscopy and snare resection (procedure)
C0472983|Endoscopic laser destruction of lesion of esophagus using rigid esophagoscope
C0472983|Endoscopic laser destruction of lesion of oesophagus using rigid oesophagoscope
C0472983|Rigid esophagoscopy and laser
C0472983|Rigid oesophagoscopy and laser
C0472983|Rigid esophagoscopy and laser (procedure)
C0472980|Endoscopic cauterisation of lesion of oesophagus using rigid oesophagoscope
C0472980|Endoscopic cauterization of lesion of esophagus using rigid esophagoscope
C0472980|Rigid oesophagoscopy and cauterisation
C0472980|Rigid esophagoscopy and cauterization
C0472980|Rigid esophagoscopy and cauterization (procedure)
C0472988|Endoscopic injection sclerotherapy to varices of esophagus using rigid esophagoscope
C0472988|Endoscopic injection sclerotherapy to varices of oesophagus using rigid oesophagoscope
C0472988|Rigid esophagoscopy and injection sclerotherapy of varices
C0472988|Rigid oesophagoscopy and injection sclerotherapy of varices
C0472988|Rigid esophagoscopy and injection sclerotherapy of varices (procedure)
C0472951|Rigid esophagoscopic banding of esophageal varices
C0472951|Rigid oesophagoscopic banding of oesophageal varices
C0472951|Rigid esophagoscopy and banding of esophageal varices
C0472951|Rigid oesophagoscopy and banding of oesophageal varices
C0472951|Rigid esophagoscopy and banding of esophageal varices (procedure)
C0472965|Rigid esophagoscopy with removal of foreign body
C0472965|esophagoscopy foreign body removal
C0472965|rigid esophagoscopy with foreign body removal (treatment)
C0472965|rigid esophagoscopy with foreign body removal
C0472965|Endoscopic removal of foreign body from esophagus using rigid esophagoscope
C0472965|Endoscopic removal of foreign body from oesophagus using rigid oesophagoscope
C0472965|Rigid esophagoscopy and removal of foreign body
C0472965|Rigid oesophagoscopy and removal of foreign body
C0472965|Rigid esophagoscopy and removal of foreign body (procedure)
C0472972|Endoscopic balloon dilation of esophagus using rigid esophagoscope
C0472972|Endoscopic balloon dilation of oesophagus using rigid oesophagoscope
C0472972|Rigid esophagoscopy and balloon dilatation
C0472972|Rigid oesophagoscopy and balloon dilatation
C0472972|Rigid esophagoscopy and balloon dilatation (procedure)
C0472961|Rigid esophagoscopy with biopsy
C0472961|Diagnostic endoscopic examination of esophagus and biopsy of lesion of esophagus using rigid esophagoscope
C0472961|Diagnostic endoscopic examination of oesophagus and biopsy of lesion of oesophagus using rigid oesophagoscope
C0472961|Rigid esophagoscopy and biopsy
C0472961|Rigid oesophagoscopy and biopsy
C0472961|Rigid esophagoscopy and biopsy (procedure)
C0472857|Fiberoptic endoscopic examination of upper gastrointestinal tract and biopsy of lesion of upper gastrointestinal tract
C0472857|Fibreoptic endoscopic examination of upper gastrointestinal tract and biopsy of lesion of upper gastrointestinal tract
C0472857|Fiberoptic endoscopic examination of upper gastrointestinal tract and biopsy of lesion of upper gastrointestinal tract (procedure)
C0399776|Diagnostic endoscopic examination of duodenum NOS (procedure)
C0399776|Diagnostic endoscopic examination of duodenum NOS
C0399776|Diagnostic duodenoscopy
C0399776|Diagnostic endoscopic examination of duodenum
C0399776|Diagnostic endoscopic examination of duodenum (procedure)
C0192310|Esophagoscopy for removal of polypoid lesion
C0192310|Oesophagoscopy for removal of polypoid lesion
C0192310|Esophagoscopy for removal of polypoid lesion (procedure)
C0475192|Fiberoptic endoscopic insertion of tubal prosthesis into esophagus
C0475192|Fibreoptic endoscopic insertion of tubal prosthesis into oesophagus
C0475192|Fiberoptic esophagoscopy and insertion of tube prosthesis
C0475192|Fibreoptic oesophagoscopy and insertion of tube prosthesis
C0475192|Fiberoptic esophagoscopy and insertion of tube prosthesis (procedure)
C0472996|Endoscopic insertion of tubal prosthesis into esophagus using rigid esophagoscope
C0472996|Endoscopic insertion of tubal prosthesis into oesophagus using rigid oesophagoscope
C0472996|Rigid esophagoscopy and insertion of tube prosthesis
C0472996|Rigid oesophagoscopy and insertion of tube prosthesis
C0472996|Rigid esophagoscopy and insertion of tube prosthesis (procedure)
C0472855|Diagnostic fiberoptic endoscopic examination of upper gastrointestinal tract NOS
C0472855|Diagnostic fibreoptic endoscopic examination of upper gastrointestinal tract NOS
C0472855|Diagnostic fiberoptic endoscopic examination of upper gastrointestinal tract NOS (procedure)
C0472855|Diagnostic fibreoptic endoscopic examination of upper gastrointestinal tract
C0472855|Diagnostic fiberoptic endoscopic examination of upper gastrointestinal tract
C0472855|Diagnostic fiberoptic endoscopic examination of upper gastrointestinal tract (procedure)
C0192317|Esophagoscopy for direct dilation
C0192317|Oesophagoscopy for direct dilation
C0192317|Esophagoscopy for direct dilation (procedure)
C0192467|upper gastrointestinal endoscopy with directed placement of percutaneous gastrostomy-tube (treatment)
C0192467|upper gastrointestinal endoscopy with directed placement of percutaneous gastrostomy-tube
C0192467|upper GI endoscopy with directed placement of percutaneous gastrostomy-tube
C0192467|upper gastrointestinal endoscopy with directed placement of percutaneous gastrostomy tube
C0192467|Upper gastrointestinal endoscopy for directed placement of percutaneous gastrostomy tube
C0192467|Upper gastrointestinal endoscopy for directed placement of percutaneous gastrostomy tube (procedure)
C2733057|Esophagogastroduodenoscopy with endoscopic ultrasound of upper gastrointestinal tract (procedure)
C2733057|Esophagogastroduodenoscopy with endoscopic ultrasound of upper gastrointestinal tract
C2733057|Oesophagogastroduodenoscopy with endoscopic ultrasound of upper gastrointestinal tract
C2733463|Esophagogastroduodenoscopy with directed submucosal injection (procedure)
C2733463|Oesophagogastroduodenoscopy with directed submucosal injection
C2733463|Esophagogastroduodenoscopy with directed submucosal injection
C0192318|Esophagoscopy for insertion of wire to guide dilation
C0192318|ESOPH ENDOSCOPY DILATION
C0192318|Esophagoscopy, flexible, transoral; with insertion of guide wire followed by passage of dilator(s) over guide wire
C0192318|ESOPHAGOSCOPY FLEXIBLE GUIDE WIRE DILATION
C0192318|Oesophagoscopy for insertion of wire to guide dilation
C0192318|Esophagoscopy for insertion of wire to guide dilation (procedure)
C0192312|FB - Esophoscopy and removal of foreign body
C0192312|FB - Esophagoscopy and removal of foreign body
C0192312|Esophagoscopy for removal of foreign body
C0192312|Remov intralum esoph FB
C0192312|Endoscopic removal of intraluminal foreign body from esophagus without incision
C0192312|Endoscopic removal of intraluminal foreign body from oesophagus without incision
C0192312|Oesophagoscopy for removal of foreign body
C0192312|Esophagoscopy and removal of foreign body
C0192312|FB - Oesophoscopy and removal of foreign body
C0192312|Oesophagoscopy and removal of foreign body
C0192312|Esophagoscopy for removal of foreign body (procedure)
C0192312|Removal of intraluminal foreign body from esophagus without incision
C0192316|Esophagoscopy for injection of esophageal varices
C0192316|Injection of sclerosing agent into esophageal varices by endoscopy
C0192316|Endoscopic injection of esophageal varices
C0192316|Injection of esophageal varices by endoscopy
C0192316|Injection of varicose veins of esophagus by endoscopy
C0192316|Endoscopic injection of oesophageal varices
C0192316|Injection of oesophageal varices by endoscopy
C0192316|Injection of sclerosing agent into oesophageal varices by endoscopy
C0192316|Injection of varicose veins of oesophagus by endoscopy
C0192316|Oesophagoscopy for injection of oesophageal varices
C0192316|Esophagoscopy for injection of esophageal varices (procedure)
C0192316|Injection of esophageal varices by endoscopic approach
C2732453|Esophagogastroduodenoscopy with insertion of guide wire and dilation of esophagus (procedure)
C2732453|Oesophagogastroduodenoscopy with insertion of guide wire and dilation of oesophagus
C2732453|Esophagogastroduodenoscopy with insertion of guide wire and dilation of esophagus
C2122145|fiberoptic duodenoscopy (procedure)
C2122145|fiberoptic duodenoscopy
C2122145|fiberoptic examinations duodenoscopy
C0472844|fiberoptic esophagoscopy (procedure)
C0472844|fiberoptic examinations esophagoscopy
C0472844|fiberoptic esophagoscopy
C0472844|Fibreoptic oesophagoscopy
C0472844|Flexible esophagoscopy
C0472844|Flexible oesophagoscopy
C0017195|Gastroscopies
C0017195|Gastroscopy
C0017195|fiberoptic examinations gastroscopy
C0017195|gastroscopy (procedure)
C0017195|Endoscopy of stomach
C0017195|Endoscopy of stomach (procedure)
C0017195|upper endoscopy
C0017195|Endoscopy of stomach, NOS
C0017195|Gastroscopy, NOS
C2207161|esophagogastroduodenoscopy w/ directed submucousal injection
C2207161|esophagogastroduodenoscopy with directed submucousal injection (procedure)
C2207161|esophagogastroduodenoscopy with directed submucousal injection
C2207161|esophagogastroduodenoscopy with directed submucousal injection(s)
C0192674|esophagogastroduodenoscopy with biopsy (procedure)
C0192674|esophagogastroduodenoscopy with biopsy
C0192674|Upper gastrointestinal endoscopy with biopsy
C0192674|Retired procedure (procedure) [P1-56735]
C0192674|Retired procedure [P1-56735]
C0192674|Biopsy of the esophagus, stomach, and/or upper small bowel using an endoscope
C0192674|Upper gastrointestinal endoscopy; biopsy
C0399616|Gastresophagoscopy via gastrotomy
C0399616|Gastroesophagoscopy via gastrotomy
C0399616|Gastrooesophagoscopy via gastrotomy
C0399616|Esophagogastroscopy via gastrotomy
C0399616|Oesophagogastroscopy via gastrotomy
C0399616|Oesophagogastroscopy via gastrotomy (procedure)
C0399616|Esophagogastroscopy via gastrotomy (procedure)
C0192470|Esophagogastroscopy through stoma
C0192470|Oesophagogastroscopy through stoma
C0192470|Esophagogastroscopy through stoma (procedure)
C0472851|rigid esophagoscopy (treatment)
C0472851|rigid esophagoscopy
C0472851|Rigid oesophagoscopy
C0472851|Rigid esophagoscopy (procedure)
C0192656|Oesophagogastroduodenoscopy through stoma
C0192656|Esophagogastroduodenoscopy through stoma
C0192656|Esophagogastroduodenoscopy through stoma (procedure)
C0192656|Esophagogastroduodenoscopy through stoma (procedure) [Ambiguous]
C2960085|Endoscopy of upper gastrointestinal tract and excision of polyp of esophagus
C2960085|Endoscopy of upper gastrointestinal tract and excision of polyp of oesophagus
C2960085|Oesophagogastroduodenoscopy and polypectomy of oesophagus
C2960085|Esophagogastroduodenoscopy and polypectomy of esophagus
C2960085|Endoscopy of upper gastrointestinal tract and excision of polyp of esophagus (procedure)
C2960784|Endoscopy and biopsy of upper gastrointestinal tract (procedure)
C2960784|Esophagogastroduodenoscopy and biopsy
C2960784|Endoscopy and biopsy of upper gastrointestinal tract
C2960784|Oesophagogastroduodenoscopy and biopsy
C2959366|Endoscopy of upper gastrointestinal tract and dilation of esophageal stricture (procedure)
C2959366|Endoscopy of upper gastrointestinal tract and dilation of oesophageal stricture
C2959366|Endoscopy of upper gastrointestinal tract and dilation of esophageal stricture
C2959366|Esophagogastroduodenoscopy and dilation of esophageal stricture
C2959366|Oesophagogastroduodenoscopy and dilation of oesophageal stricture
C2959746|Esophagogastroduodenoscopy and mucosectomy of duodenum
C2959746|Endoscopy of upper gastrointestinal tract and excision of mucosa of duodenum (procedure)
C2959746|Oesophagogastroduodenoscopy and mucosectomy of duodenum
C2959746|Endoscopy of upper gastrointestinal tract and excision of mucosa of duodenum
C2960325|Endoscopy of upper gastrointestinal tract and excision of mucosa of stomach (procedure)
C2960325|Endoscopy of upper gastrointestinal tract and excision of mucosa of stomach
C2960325|Esophagogastroduodenoscopy and mucosectomy of stomach
C2960325|Oesophagogastroduodenoscopy and mucosectomy of stomach
C2959681|Endoscopy of upper gastrointestinal tract and excision of polyp of duodenum
C2959681|Oesophagogastroduodenoscopy and polypectomy of duodenum
C2959681|Endoscopy of upper gastrointestinal tract and excision of polyp of duodenum (procedure)
C2959681|Esophagogastroduodenoscopy and polypectomy of duodenum
C2959668|Endoscopy of upper gastrointestinal tract and removal of foreign body from esophagus
C2959668|Endoscopy of upper gastrointestinal tract and removal of foreign body from esophagus (procedure)
C2959668|Endoscopy of upper gastrointestinal tract and removal of foreign body from oesophagus
C2959668|Oesophagogastroduodenoscopy and removal of foreign body from oesophagus
C2959668|Esophagogastroduodenoscopy and removal of foreign body from esophagus
C2960120|Oesophagogastroduodenoscopy and insertion of oesophageal stent
C2960120|Endoscopy of upper gastrointestinal tract and insertion of esophageal stent
C2960120|Endoscopy of upper gastrointestinal tract and insertion of oesophageal stent
C2960120|Esophagogastroduodenoscopy and insertion of esophageal stent
C2960120|Endoscopy of upper gastrointestinal tract and insertion of esophageal stent (procedure)
C2960528|Oesophagogastroduodenoscopy and dilation of gastric cardia
C2960528|Endoscopy of upper gastrointestinal tract and dilation of gastric cardia
C2960528|Esophagogastroduodenoscopy and dilation of gastric cardia
C2960528|Endoscopy of upper gastrointestinal tract and dilation of gastric cardia (procedure)
C2960061|Endoscopy of upper gastrointestinal tract and tattooing (procedure)
C2960061|Endoscopy of upper gastrointestinal tract and tattooing
C2960061|Esophagogastroduodenoscopy and tattooing
C2960061|Oesophagogastroduodenoscopy and tattooing
C2959967|Endoscopy of upper gastrointestinal tract and dilation of gastric stoma
C2959967|Endoscopy of upper gastrointestinal tract and dilation of gastric stoma (procedure)
C2960407|Esophagogastroduodenoscopy and injection of gastric varices
C2960407|Endoscopy of upper gastrointestinal tract and injection of varix of stomach (procedure)
C2960407|Oesophagogastroduodenoscopy and injection of gastric varices
C2960407|Endoscopy of upper gastrointestinal tract and injection of gastric varices
C2960407|Endoscopy of upper gastrointestinal tract and injection of varix of stomach
C2959433|Endoscopy of upper gastrointestinal tract and excision of mucosa of esophagus (procedure)
C2959433|Endoscopy of upper gastrointestinal tract and excision of mucosa of oesophagus
C2959433|Esophagogastroduodenoscopy and mucosectomy of esophagus
C2959433|Endoscopy of upper gastrointestinal tract and excision of mucosa of esophagus
C2959433|Oesophagogastroduodenoscopy and mucosectomy of oesophagus
C2960354|Endoscopy of upper gastrointestinal tract and excision of polyp of stomach (procedure)
C2960354|Esophagogastroduodenoscopy and polypectomy of stomach
C2960354|Endoscopy of upper gastrointestinal tract and excision of polyp of stomach
C2960354|Oesophagogastroduodenoscopy and polypectomy of stomach
C2959632|Endoscopy of upper gastrointestinal tract and banding of varix of esophagus (procedure)
C2959632|Esophagogastroduodenoscopy and banding of esophageal varices
C2959632|Endoscopy of upper gastrointestinal tract and banding of varix of oesophagus
C2959632|Endoscopy of upper gastrointestinal tract and banding of esophageal varices
C2959632|Endoscopy of upper gastrointestinal tract and banding of oesophageal varices
C2959632|Endoscopy of upper gastrointestinal tract and banding of varix of esophagus
C2959632|Oesophagogastroduodenoscopy and banding of oesophageal varices
C2959721|Endoscopy of upper gastrointestinal tract and injection of varix of esophagus (procedure)
C2959721|Esophagogastroduodenoscopy and injection of esophageal varices
C2959721|Endoscopy of upper gastrointestinal tract and injection of esophageal varices
C2959721|Endoscopy of upper gastrointestinal tract and injection of varix of oesophagus
C2959721|Endoscopy of upper gastrointestinal tract and injection of oesophageal varices
C2959721|Endoscopy of upper gastrointestinal tract and injection of varix of esophagus
C2959721|Oesophagogastroduodenoscopy and injection of oesophageal varices
C2959927|Oesophagogastroduodenoscopy and banding of gastric varices
C2959927|Endoscopy of upper gastrointestinal tract and banding of varix of stomach
C2959927|Endoscopy of upper gastrointestinal tract and banding of gastric varices
C2959927|Endoscopy of upper gastrointestinal tract and banding of varix of stomach (procedure)
C2959927|Esophagogastroduodenoscopy and banding of gastric varices
C2960375|Oesophagogastroduodenoscopy and ligation of duodenal varices
C2960375|Endoscopy of upper gastrointestinal tract and ligation of duodenal varices
C2960375|Endoscopy of upper gastrointestinal tract and ligation of varix of duodenum (procedure)
C2960375|Endoscopy of upper gastrointestinal tract and ligation of varix of duodenum
C2960375|Esophagogastroduodenoscopy and ligation of duodenal varices
C0014873|Esophagoscopies
C0014873|Esophagoscopy
C0014873|Oesophagoscopy
C0014873|esophagoscopy (treatment)
C0014873|Endoscopy Procedures on the Esophagus
C0014873|Endoscopic examination of esophagus
C0014873|Endoscopic examination of oesophagus
C0014873|Endoscopy of esophagus (procedure)
C0014873|Endoscopy of esophagus
C0014873|Endoscopy of oesophagus
C0014873|Endoscopy of esophagus, NOS
C0014873|Esophagoscopy, NOS
C0014873|Oesophagoscopy, NOS
C0192471|esophagogastroscopy operative
C0192471|esophagogastroscopy operative (treatment)
C0192471|Operative esophagogastroscopy
C0192471|Operative oesophagogastroscopy
C0192471|Operative esophagogastroscopy (procedure)
C0013301|Duodenoscopies
C0013301|Duodenoscopy
C0013301|Duodenoscopy (procedure)
C0013301|Endoscopy of duodenum
C0013301|Duodenoscopy, NOS
C0013301|Endoscopy of duodenum, NOS
C0192655|esophagogastroduodenoscopy operative
C0192655|esophagogastroduodenoscopy operative (treatment)
C0192655|Operative esophagogastroduodenoscopy
C0192655|Operative oesophagogastroduodenoscopy
C0192655|Operative esophagogastroduodenoscopy (procedure)
C2095043|upper gastrointestinal endoscopy, simple primary exam
C2095043|upper gastrointestinal endoscopy, simple primary exam (procedure)
C2095043|upper GI endoscopy, simple primary exam
C2095643|upper gastrointestinal endoscopy (diagnostic)
C2095643|upper GI endoscopy diagnostic
C2095643|upper gastrointestinal diagnostic endoscopy
C2095643|upper gastrointestinal diagnostic endoscopy (procedure)
C2095643|Diagnostic upper gastrointestinal endoscopy
C3507762|esophagogastroduodenoscopy with optic endomicroscopy
C3507762|esophagogastroduodenoscopy with optic endomicroscopy (procedure)
C0192466|Oesophagogastroscopy
C0192466|Esophagogastroscopy
C0192466|Endoscopic examination of esophagus and stomach
C0192466|Endoscopic examination of oesophagus and stomach
C0192466|Esophagogastroscopy (procedure)
C0192466|esophagogastroscopy (treatment)
C3694781|esophagogastroduodenoscopy transoral flex w/ optic endomicroscopy (procedure)
C3694781|esophagogastroduodenoscopy transoral flex w/ optic endomicroscopy
C3694780|esophagogastroduodenoscopy transoral flexible (procedure)
C3694780|esophagogastroduodenoscopy transoral flexible
C3694780|Esophagogastroduodenoscopy, flexible, transoral
C4038699|Esophagogastroduodenoscopy and dilatation of duodenum
C4038699|Endoscopy of upper gastrointestinal tract and dilatation of duodenum (procedure)
C4038699|Endoscopy of upper gastrointestinal tract and dilatation of duodenum
C4038699|Oesophagogastroduodenoscopy and dilatation of duodenum
C4065150|esophagogastroduodenoscopy with esophagogastric fundoplasty
C4065150|esophagogastroduodenoscopy with esophagogastric fundoplasty (treatment)
C0810405|Esophagogastroduodenoscopy (EGD) with biopsy
C0176784|Egd with closed biopsy
C0176784|Esophagogastroduodenoscopy [EGD] with closed biopsy
C0176784|Esophagogastroduodenoscopy with closed biopsy
C0176784|Biopsy of one or more sites involving esophagus, stomach and/or duodenum
C0399617|Diagnostic gastroscopy via stoma
C0399617|Diagnostic gastroscopy via stoma (procedure)
C0009556|complete colonoscopy
C0009556|complete colonoscopy (treatment)
C0009556|Total colonoscopy
C0009556|Total colonoscopy (procedure)
C0192910|COLONOSCOPY STOMA W/RMVL FOREIGN BODY
C0192910|Colonoscopy through stoma with removal of foreign body
C0192910|Retired procedure (procedure) [P1-57731]
C0192910|Retired procedure [P1-57731]
C0192910|Colonoscopy through stoma; with removal of foreign body(s)
C0192910|COLONOSCOPY FOR FOREIGN BODY
C0016234|Flexible Fiberoptic Sigmoidoscopy
C0016234|fiberoptic examinations sigmoidoscopy
C0016234|fiberoptic sigmoidoscopy (procedure)
C0016234|fiberoptic sigmoidoscopy
C0016234|fiberoptic sigmoidoscopy (treatment)
C0016234|Flexible sigmoidoscopy
C0016234|Sigmoidoscopy, flexible
C0016234|Fibreoptic sigmoidoscopy
C0016234|FS - Flexible sigmoidoscopy
C0016234|FOS - Fiberoptic sigmoidoscopy
C0016234|FOS - Fibreoptic sigmoidoscopy
C0016234|Flexible fiberoptic sigmoidoscopy (procedure)
C0016234|Flexible fibreoptic sigmoidoscopy
C0372134|Flexible colonoscopy proximal to splenic flexure with removal of foreign body
C0372134|Colonoscopy, flexible; with removal of foreign body(s)
C0372134|COLONOSCOPY FLX W/REMOVAL OF FOREIGN BODY(S)
C0372134|COLONOSCOPY W/FB REMOVAL
C0192899|colonoscopy with rigid sigmoidoscope through colotomy (procedure)
C0192899|Colonoscopy with rigid sigmoidoscope through colotomy
C0192901|colonoscopy (fiberoptic) with biopsy
C0192901|fiberoptic colonoscopy with biopsy (procedure)
C0192901|fiberoptic colonoscopy with biopsy
C0192901|Fibreoptic colonoscopy with biopsy
C0192902|Retired procedure [P1-57722]
C0192902|Retired procedure (procedure) [P1-57722]
C0192903|Retired procedure (procedure) [P1-57723]
C0192903|Retired procedure [P1-57723]
C0192904|Retired procedure (procedure) [P1-57724]
C0192904|Retired procedure [P1-57724]
C0192905|Retired procedure [P1-57725]
C0192905|Retired procedure (procedure) [P1-57725]
C0192906|Retired procedure [P1-57726]
C0192906|Retired procedure (procedure) [P1-57726]
C0192909|fiberoptic colonoscopy via colostomy (procedure)
C0192909|fiberoptic colonoscopy via colostomy
C0192909|fiberoptic examinations colonoscopy via colostomy
C0192909|Fiberoptic colonoscopy through colostomy
C0192909|Endoscopy of colon through artificial stoma
C0192909|Colonoscopy through artificial stoma
C0192909|Fiberoptic colonoscopy through colostomy (procedure)
C0192909|Fibreoptic colonoscopy through colostomy
C0192913|Retired procedure [P1-57734]
C0192913|Retired procedure (procedure) [P1-57734]
C0192914|Retired procedure (procedure) [P1-57735]
C0192914|Retired procedure [P1-57735]
C0192915|Retired procedure (procedure) [P1-57736]
C0192915|Retired procedure [P1-57736]
C0192916|Retired procedure [P1-57737]
C0192916|Retired procedure (procedure) [P1-57737]
C0037075|Proctosigmoidoscopies
C0037075|Proctosigmoidoscopy
C0037075|Sigmoidoscopies
C0037075|Sigmoidoscopy
C0037075|Sigmoidoscopy (procedure)
C0037075|SIGGY - Sigmoidoscopy
C0037075|SIGy - Sigmoidoscopy
C0037075|Sigmoidoscopy, NOS
C0009378|Colonoscopies
C0009378|Colonoscopy
C0009378|Colonoscopy (procedure)
C0009378|colonoscopy (treatment)
C0009378|Endoscopy Procedures on the Rectum
C0009378|Endoscopic examination of colon
C0009378|Endoscopy of colon
C0009378|Colonoscopy, NOS
C0009378|Endoscopy of colon, NOS
C0009378|Colonoscopy [Ambiguous]
C0751041|SURG PROCEDURES COLONOSCOPIC
C0751041|SURG COLONOSCOPIC
C0751041|COLONOSCOPIC SURG PROCEDURES
C0751041|COLONOSCOPIC SURG
C0751041|Colonoscopic Surgical Procedure
C0751041|Procedure, Colonoscopic Surgical
C0751041|Procedures, Colonoscopic Surgical
C0751041|Surgical Procedure, Colonoscopic
C0751041|Colonoscopic Surgeries
C0751041|Surgeries, Colonoscopic
C0751041|Colonoscopic Surgery
C0751041|Surgical Procedures, Colonoscopic
C0751041|Surgery, Colonoscopic
C0751041|Colonoscopic Surgical Procedures
C2732814|Colonoscopy through colostomy with endoscopic biopsy of colon
C2732814|Colonoscopy through colostomy with endoscopic biopsy of colon (procedure)
C2732814|colonoscopy via colostomy with endoscopic biopsy (procedure)
C2732814|colonoscopy via colostomy with endoscopic biopsy
C1882982|Screening Colonoscopy
C1882982|Screening colonoscopy (procedure)
C1882982|Screening colonoscopy NOS
C2960146|Colonoscopy and excision of mucosa of colon
C2960146|Colonoscopy and excision of mucosa of colon (procedure)
C2960146|Colonoscopy and colonic mucosectomy
C2960146|colonoscopy with excision of mucosa of colon (treatment)
C2960146|colonoscopy with excision of mucosa of colon
C2960408|Colonoscopy and biopsy of colon (procedure)
C2960408|Colonoscopy and biopsy of colon
C2960062|Colonoscopy and tattooing (procedure)
C2960062|Colonoscopy and tattooing
C2960062|colonoscopy (fiberoptic) with tattooing (procedure)
C2960062|colonoscopy (fiberoptic) with tattooing
C3274817|Index Colonoscopy
C3274817|Baseline Colonoscopy
C0399623|intraoperative colonoscopy
C0399623|intraoperative colonoscopy (procedure)
C0399623|Transab lg bowel endosc
C0399623|Operative endoscopy of colon
C0399623|Operative colonoscopy
C0399623|Transabdominal endoscopy of large intestine
C0399623|Intraoperative endoscopy of large intestine
C1298662|Endoscopic insertion of temporary colonic stent (procedure)
C1298662|Endoscopic insertion of temporary colonic stent
C0585464|Laparoscopic right hemicolectomy
C0585464|Lap right hemicolectomy
C0585464|Laparoscopic-assisted right colectomy
C0585464|Laparoscopic-assisted right colectomy (procedure)
C1298663|Endoscopic insertion of permanent colonic stent (procedure)
C1298663|Endoscopic insertion of permanent colonic stent
C0192929|Proctosigmoidoscopy with biopsy
C0192929|Proctosigmoidoscopy with biopsy (procedure)
C0035622|rigid proctosigmoidoscopy (treatment)
C0035622|rigid proctosigmoidoscopy
C0035622|Rigid proctosigmoidoscpy
C0035622|Proctosigmoidoscopy.rigid
C0035622|Proctosigmoidoscopy, rigid
C0035622|Rigid proctosigmoidoscopy (procedure)
C0192927|Proctosigmoidoscopy by transabdominal approach
C0192927|Proctosigmoidoscopy by transabdominal approach (procedure)
C0578726|Endoscopic biopsy of lesion of colon
C0578726|Endoscopic biopsy of lesion of colon (procedure)
C0192933|Proctosigmoidoscopy for dilation
C0192933|Proctosigmoidoscopy for dilation (procedure)
C0521258|Laparoscopic-assisted left colectomy
C0521258|Laparoscopic-assisted left colectomy (procedure)
C0192900|Fiberoptic colonoscopy
C0192900|Fiberoptic colonoscopy, NOS
C0192900|Fibreoptic colonoscopy, NOS
C0192900|fiberoptic colonoscopy (procedure)
C0192900|Fibreoptic colonoscopy
C0192900|Colonoscopy (procedure)
C0192900|Fiberoptic colonoscopy (procedure) [Ambiguous]
C0192900|Flexible fiberoptic colonoscopy
C2095474|complete colonoscopy of hepatic flexure (treatment)
C2095474|complete colonoscopy of hepatic flexure
C2095866|complete colonoscopy of sigmoid colon with dilation (treatment)
C2095866|complete colonoscopy of sigmoid colon with dilation
C2095475|complete colonoscopy of transverse colon (treatment)
C2095475|complete colonoscopy of transverse colon
C2095473|complete colonoscopy of ascending colon
C2095473|complete colonoscopy of ascending colon (treatment)
C2095478|complete colonoscopy of sigmoid colon
C2095478|complete colonoscopy of sigmoid colon (treatment)
C2095476|complete colonoscopy of splenic flexure (treatment)
C2095476|complete colonoscopy of splenic flexure
C2095477|complete colonoscopy of descending colon
C2095477|complete colonoscopy of descending colon (treatment)
C0588165|Check colonoscopy (procedure)
C0588165|Check colonoscopy
C0588165|colonoscopy check
C0588165|check colonoscopy (treatment)
C0554063|Therapeutic Colonoscopy
C0554063|colonoscopy therapeutic
C0554063|Therapeutic colonoscopy (treatment)
C0554063|Therapeutic colonoscopy (procedure)
C0399622|open colonoscopy (treatment)
C0399622|Open colonoscopy
C0399622|Open colonoscopy (procedure)
C3869456|Colonoscopy, flexible
C4040527|Colonoscopy and dilatation of stricture of colon
C4040527|Colonoscopy and dilatation of stricture of colon (procedure)
C4039452|Colonoscopy using X-ray guidance
C4039452|Colonoscopy using X-ray guidance (procedure)
C4038675|Colonoscopy using fluoroscopic guidance
C4038675|Fluoroscopy guided colonoscopy
C4038675|Colonoscopy using fluoroscopic guidance (procedure)
C0400018|Diagnostic Colonoscopy
C0400018|Diagnostic endoscopic examination on colon
C0400018|Diagnostic endoscopic examination of colon NOS
C0400018|Diagnostic endoscopic examination of colon NOS (procedure)
C0400018|diagnostic endoscopy of colon
C0400018|colon endoscopy (diagnostic)
C0400018|diagnostic endoscopy of colon (procedure)
C0400018|Diagnostic endoscopic examination on colon (procedure)
C0399625|colonoscopy (fiberoptic) limited
C0399625|limited colonoscopy (fiberoptic) (procedure)
C0399625|limited colonoscopy (fiberoptic)
C0399625|Limited colonoscopy
C0399625|Limited colonoscopy (procedure)
C0863836|Endoscopy of descending colon
C1960976|Diagnostic endoscopic examination of colonic pouch and biopsy of colonic pouch using fiberoptic sigmoidoscope (procedure)
C1960976|Diagnostic endoscopic examination of colonic pouch and biopsy of colonic pouch using fiberoptic sigmoidoscope
C1960976|Diagnostic endoscopic examination of colonic pouch and biopsy of colonic pouch using fibreoptic sigmoidoscope
C1960975|Diagnostic endoscopic examination of colonic pouch and biopsy of colonic pouch using colonoscope (procedure)
C1960975|Diagnostic endoscopic examination of colonic pouch and biopsy of colonic pouch using colonoscope
C1960975|colonoscopy (fiberoptic) of colonic pouch with biopsy
C1960975|colonoscopy (fiberoptic) of colonic pouch with biopsy (procedure)
C1960974|Diagnostic endoscopic examination of colonic pouch and biopsy of colonic pouch using rigid sigmoidoscope (procedure)
C1960974|Diagnostic endoscopic examination of colonic pouch and biopsy of colonic pouch using rigid sigmoidoscope
