C0489786|Height
C0005890|Body Height
C0424645|Standing height
C0231248|Body height normal for age
C0487985|Body height:Length:Point in time:^Patient:Quantitative
C0424639|Height / growth measure
C1861519|Short stature, moderate
C1861519|Moderately short stature
C1861519|Moderate short stature
C1849937|Short-limbed dwarfism
C1849937|Short stature, disproportionate short limb
C1849937|Short stature, disproportionate short-limb
C1849937|Short limb dwarfism, disproportionate
C1849937|Short-limb dwarfism
C1849937|Short limb dwarfism
C1849937|Dwarfism, short-limbed
C1849937|Dwarfism, micromelic
C1849937|Dwarfism, short-limb
C1849937|Dwarfism, disproportionate short-limb
C1849937|Brachymelic dwarfism
C1849937|Micromelic dwarfism
C1849937|Disproportionate short-limb short stature
C1849937|Disproportionate short limb dwarfism
C1853173|Normal birth length
C1853173|Birth length normal
C2678391|Birth length below 5th percentile
C2673388|Average adult height 114 cm
C2676293|Birth length below 0.3 percentile
C2673284|Short stature (type II, infantile and juvenile)
C2673718|Decreased stature
C0557899|Increased height
C0557899|Height increased
C0557899|Height increased (finding)
C2675900|Normal or reduced
C2674444|Short stature (childhood)
C2674444|Short stature in childhood
C2674444|Short stature (in childhood)
C2678144|Short stature (5th percentile)
C2732728|Body height decreased
C2732728|Decreased body height
C2732728|Decreased height
C2732728|Short for age
C2732728|Short stature for age
C2732728|Short stature for age (finding)
C2732728|Decreased;height
C2677758|Short stature, final adult height 150-160cm
C1861927|Short limb dwarfism, prenatal onset
C1861927|Dwarfism, short-limb, prenatal onset
C2674171|Dwarfism, lethal micromelic
C2674171|Lethal short-limbed dwarfism
C2674171|Lethal micromelic dwarfism
C2674171|Lethal short-limbed short stature
C2030323|height ___ percentile for age
C2030323|height percentile for age
C2030323|height percentile for age (physical finding)
C2030328|height proportional to weight
C2030328|height proportional to weight (physical finding)
C2030328|the height was proportional to the weight
C2367600|father's height
C2367600|father's height (physical finding)
C2367341|mother's height
C2367341|mother's height (physical finding)
C2367313|mid-parental height
C2367313|mid-parental height (physical finding)
C2243104|span (physical finding)
C2243104|span
C2243104|span - body measurement finding
C2017863|span versus height
C2017863|span versus height (physical finding)
C2030327|height of upper segment of body greater than lower segment (physical finding)
C2030327|height of upper segment of body greater than lower segment
C2030327|the upper body segment height was greater than the lower body segment
C2030326|height of lower segment of body greater than upper segment (physical finding)
C2030326|height of lower segment of body greater than upper segment
C2030326|the lower body segment height was greater than the upper body segment
C2228524|excessive height
C2228524|excessive height (physical finding)
C0349588|Short stature
C0349588|[D]Short stature (context-dependent category)
C0349588|Height less than 3rd percentile
C0349588|short stature (physical finding)
C0349588|short stature was noted
C0349588|Short stature NOS
C0349588|Short;stature
C0349588|Small stature
C0349588|[D]Short stature (situation)
C0349588|[D]Short stature
C0349588|Short stature (finding)
C0349588|SS - Short stature
C0349588|Decreased body height
C0349588|Short stature (below 3rd percentile)
C0349588|Stature short
C0349588|short; stature
C0349588|stature; short
C0349588|Short;growth
C0017547|Gigantism
C0017547|gigantism (diagnosis)
C0017547|gigantism (physical finding)
C0017547|Giant -RETIRED-
C0017547|gigantism was noted
C0017547|Gigantism [Disease/Finding]
C0017547|Pituitary Gigantism
C0017547|Giant (disorder)
C0017547|Giant
C0017547|Genetic giant
C0017547|Normal giant
C0017547|Primordial giant
C0017547|Giantism
C0017547|Gigantism (disorder)
C0017547|gigantism; pituitary
C0017547|pituitary; gigantism
C0017547|Giant, NOS
C0017547|Giantism, NOS
C0017547|Gigantism, NOS
C0017547|Gigantism, Pituitary
C1844723|Short stature (males)
C1844723|Short stature (in males)
C2750631|Short stature (final adult height less than 152cm)
C2748450|Increased birth length
C2751301|Short stature (some)
C2751301|Short stature (in some patients)
C2751647|Growth retardation in childhood
C2749299|Short stature (postnatal onset) (97%)
C2749067|Short stature (female)
C2752046|Tall stature (>97th centile)
C2751023|Accelerated linear growth (in 1 of 2 patients)
C2751617|Short stature (if untreated)
C0424639|Height / growth measure
C0424639|Stature
C0424639|Height and growth
C0424639|Length and growth
C0424639|Observation of height and growth
C0424639|Height / growth measure (observable entity)
C3149920|Short stature, relative (in some patients)
C3150077|Short stature, mild
C3150077|Mild short stature
C3151876|Dwarfism, mild
C3148867|Short stature (3rd percentile)
C3149248|Dwarfism, mild short-limb
C3150094|Dwarfism, marked micromelic
C3148833|Short stature, disproportionate (short trunk), identifiable in childhood
C3148833|Disproportionate short stature (short trunk), identifiable in childhood
C3148833|Short-trunk dwarfism identifiable during childhood
C3148833|Childhood-onset short-trunk short stature
C3151646|Short stature, disproportionate (short trunk), identifiable late childhood-early puberty
C3149232|Short stature, mild to moderate
C3149908|Dwarfism, short-trunk, identifiable at birth
C3149908|Neonatal short-trunk short stature
C3149908|Short-trunk dwarfism identifiable at birth
C3151648|Short stature, disproportionate short-trunked (identifiable at birth)
C1855274|Short stature, disproportionate mesomelic
C1855274|Dwarfism, short limb mesomelic
C1855274|Short stature, mesomelic
C1855274|Mesomelic short stature
C1855274|Mesomelic dwarfism
C3150493|Short stature, pre- and postnatal
C3278794|Below 3rd percentile
C3280406|Increased stature
C3280830|Growth deficit affecting lower segment of body
C3276917|Short stature, prenatal and postnatal
C3277096|Short stature (deletion patients)
C3278061|Short stature, severe (in some patients)
C3276033|Less than tenth centile
C3279161|Increased height in females
C3280176|Short stature (1 patient)
C3277493|Short stature (postnatal onset) (81%)
C3275498|Less than third centile
C3280343|Adult height, average
C3279055|Tall stature (46%)
C1850171|Short-limbed dwarfism identifiable at birth
C1850171|Short-limb dwarfism identifiable neonatally
C1850171|Short-limb dwarfism identifiable at birth
C1850171|Dwarfism, neonatal short-limbed
C1850171|Short limb dwarfism recognizable at birth
C1850171|Dwarfism, short limbed, recognizable at birth
C1850171|Neonatal short-limb short stature
C1850171|Neonatal short-limbed dwarfism
C3275910|Short stature (13 of 23 patients)
C3278752|Postnatal growth delay
C3278027|Normal linear growth
C1859778|Postnatal growth failure
C1859778|Growth failure, postnatal
C1859778|Postnatal growth retardation
C1859778|Growth retardation as children
C1859778|Postnatal growth deficiency
C1859778|Postnatal growth deceleration
C1859778|Growth retardation, postnatal
C3553080|Height in third centile
C3553254|Short stature, mild (in some)
C3554766|Short stature (1 family)
C3551740|Short stature (of varying degrees)
C1853174|Short stature (adult)
C1853174|Short stature (adults)
C3553733|Short stature, disproportionate, prenatal onset
C3551528|Small birth length
C3551528|Low birth length
C3554671|less than 3rd centile (in one patient)
C3554440|Low weight (<3.5 SD below the mean)
C3550824|Short stature (in 2 of 3 siblings)
C3550931|Short stature (2/4 patients)
C3550970|Average height in adulthood
C3550969|Delayed growth spurt in puberty
C3550879|Short stature, mildly disproportionate
C3551144|Short stature (reported in 2 families)
C3553468|Low-normal height
C1857641|Marked growth retardation
C1857641|Postnatal growth retardation, severe
C1857641|Severe postnatal growth deficiency
C1857641|Severe postnatal growth retardation
C1857641|Severe postnatal growth failure
C3805986|Short stature (<25% centile)
C0024032|Birth Weight, Low
C0024032|Birth Weights, Low
C0024032|Low Birth Weights
C0024032|Low birth weight
C0024032|low birth weight (history)
C0024032|Low birthweight
C0024032|low birth weight (diagnosis)
C0024032|Subnormal birth weight
C0024032|Birth weight low
C0024032|Birth weight subnormal
C0024032|Birthweight low
C0024032|Birthweight subnormal
C0024032|Weight birth subnormal
C0024032|birthweight; low, for gestational age
C0024032|birthweight; low
C0024032|low; birthweight, for gestational age
C0024032|low; birthweight
C3806181|Birth length less than 38 cm
C1855165|Disproportionate dwarfism
C1855165|Dwarfism, disproportionate
C3806979|Short stature (rare)
C3808712|Short stature (fifth to tenth centile)
C3809260|Continued growth into adulthood (in male and female patients)
C3836210|recumbent height ___
C3836210|recumbent height
C3836210|recumbent height (physical finding)
C3836390|pre-operative height (physical finding)
C3836390|pre-operative height
C3835668|stated height
C3835668|stated height (symptom)
C0424645|standing height
C0424645|standing height ___
C0424645|Standing height (physical finding)
C0424645|Standing height (observable entity)
C0241240|Tall stature
C0241240|Increased linear growth
C0241240|Accelerated linear growth
C0241240|tall stature (physical finding)
C0241240|Increased body height
C0241240|Stature tall
C0241240|Large stature
C0241240|Tall stature (finding)
C0241240|stature; tall
C0241240|tall; stature
C3550852|Long limbs
C3550852|long limbs (physical finding)
C0424646|sitting height ___
C0424646|sitting height ___ (physical finding)
C0424646|Sitting height
C0424646|Sitting height (observable entity)
C4014547|Tall stature (+3 S.D)
C4011875|Short trunk, not evident at birth
C4012355|Long birth length (in some patients)
C4014677|Short stature (-3.8 to -5.2 SD)
C3150281|Fetal overgrowth
C4015717|Birth length >97th percentile
C4011876|Reduced upper- to lower-body segment ratio
C4012406|Increased height velocity (+6.1 SD)
C4015086|Short stature (in 1 of 2 sibs)
C4012405|Tall stature (+3.4 SD)
C4014716|Poor linear growth
C4014065|Postnatal growth failure (in some patients)
C4012972|Proportionate short stature at birth
C4014691|Tall stature (+2 to +4 SD, present at birth)
C3808925|Growth retardation (in some patients)
C4015568|Short stature (79%)
C4028803|long slender trunk (physical finding)
C4028803|long slender trunk
C1849934|Birth length < 3rd percentile (63%)
C1843420|Short stature (less common)
C1842215|Adult male height 142-169 cm
C1850172|Adult height 92-108 cm
C1850289|Dwarfism, identifiable at birth
C1866224|Normal to increased birth length
C0878660|Proportionate small stature
C0878660|Proportionate short stature
C0878660|Short stature, proportionate
C1854709|Birth length 1.5-2 S.D. below mean
C1854762|Adult height 110-140 cm
C1854812|Adult height 82 to 115 cm
C1854812|Adult height 82-115 cm
C1851058|Short stature (-4 to -6 S.D. below mean)
C1860171|Average adult male height, 100.5cm
C1854922|Birth length less than normal
C0013336|Dwarfism
C0013336|Nanism
C0013336|Constitutional dwarfism
C0013336|Physiologic dwarfism
C0013336|Constitutional short stature
C0013336|Constitutional short stature (disorder)
C0013336|[D]Short stature, constitutional (context-dependent category)
C0013336|Short stature, severe
C0013336|Proportionate dwarfism
C0013336|dwarfism (diagnosis)
C0013336|Pure dwarf
C0013336|Normal dwarf
C0013336|Normal dwarfism
C0013336|True dwarf
C0013336|Nanosomia
C0013336|Pure dwarfism
C0013336|True dwarfism
C0013336|constitutional dwarfism (diagnosis)
C0013336|Runting
C0013336|Short stature disorder
C0013336|Dwarf
C0013336|Dwarfism [Disease/Finding]
C0013336|Short stature
C0013336|Little person
C0013336|Dwarfism (disorder)
C0013336|[D]Short stature, hereditary
C0013336|[D]Short stature, constitutional
C0013336|[D]Short stature, constitutional (situation)
C0013336|Primordial dwarfism
C0013336|Primordial dwarf
C0013336|Nanosoma
C0013336|Severe short stature
C0013336|Dwarfism NOS
C0013336|Primordial dwarfism (disorder)
C0013336|Short stature disorder (disorder)
C0013336|constitutional; dwarfism
C0013336|dwarfism; constitutional
C0013336|short; stature, constitutional
C0013336|stature; short, constitutional
C0013336|Dwarf, NOS
C0013336|Dwarfism, NOS
C0013336|Dwarfism (disorder) [Ambiguous]
C1849359|Birth length less than 40cm
C1855198|Average adult height, 107 to 143 cm
C1856225|Average male height 155-157 cm
C1856226|Average female height 152 cm
C1834972|Adult height 130-160cm
C1867868|Length deceleration in first few months
C1867871|Steady childhood growth
C1865835|Adult female height 152-167cm
C1854706|Short stature, prenatal onset
C1854706|Prenatal onset of short stature
C1860407|Short stature (in patients with childhood-onset)
C1859418|Average adult female height 144cm
C1835758|Short stature (less than tenth percentile)
C1861928|Birth length 35-49 cm
C1855724|Height in childhood <5th percentile
C1851729|Growth parallels curve at or above 95%
C1845249|Short stature (less than 3rd percentile)
C1849337|Short stature (postnatal onset)
C1849337|Short stature, postnatal onset
C1849527|Average adult male height 142 cm (4'8")
C0587053|Normal height
C0587053|Normal height (finding)
C1846797|Short stature, severe disproportionate
C1846797|Severely disproportionate short stature
C1832820|Short stature (adult height <152cm)
C1835111|Mean adult height 191.3 +/- 9 cm for males
C1839504|Short stature (<10th percentile for age)
C1839635|Increased birth length (>90th percentile)
C1859880|Height loss secondary to spinal changes
C1855650|Birth length <3rd percentile
C1855650|Birth length less than 3rd percentile
C1855650|Birth length < 3rd percentile
C1834319|Short stature (in some cases)
C1857259|Adult height 100-140cm
C1851539|Final adult height 145-170cm
C1857399|Short stature in first year of life
C1864856|Tall stature (male mean adult height 195.6cm, female mean adult height 177.8cm)
C1846844|Normal stature
C1836592|Short trunk short stature (<3rd - 50th percentile)
C1846435|Short stature, disproportionate (short trunk)
C1846435|Short-trunked dwarfism
C1846435|Disproportionate short-trunk short stature
C1846435|Disproportionate short-trunked short stature
C1846435|Disproportionate short-trunked dwarfism
C1858451|Height 2 S.D. below expected height
C1854708|Adult female height 126-151 cm
C1835465|Short stature, postnatal
C1835465|Postnatal short stature
C1861720|Length at or greater than 97th percentile through early adolescence
C1861845|Normal in majority of cases
C1866730|Symmetrical rhizomelic limb shortening
C1866730|Rhizomelic limb shortening
C1866730|Rhizomelic dwarfism
C1866730|Rhizomelia
C1866730|Short stature, rhizomelic
C1866730|Rhizomelic shortening
C1866730|Rhizomelic short stature
C1866730|Rhizomelic short limbs
C1859417|Average adult male height 151cm
C1856284|Final adult height normal
C1856284|Normal final adult height
C1833749|Short stature, often below 5th percentile
C1863420|Mean male adult height, 131 cm
C1833775|Height often shorter than unaffected family members
C1840336|Final height, 125 to 160 cm
C1856995|Average adult height, 109 to 152 cm
C1860148|Short stature (<25th percentile)
C1857258|Mean birth length 42cm, specific growth curve available
C1866709|Dwarfism, short-trunk, short-limbed
C1866721|Final adult height, 84-128cm
C1851987|Adult height 135cm to normal
C1834951|Final adult height 106-145cm
C1867125|Average adult female height 147 cm
C1849528|Average adult female height 135 (4'5")
C1836324|Short stature (<3rd percentile)
C1836875|Short stature, disproportionate short-limbed (dwarfism)
C1864359|Final adult height 38-49 inches
C1864360|Small-normal birth length
C1865834|Adult male height 167-173cm
C1867487|Short-limb dwarfism identifiable during childhood
C1867487|Childhood onset short-limb short stature
C1835113|Disproportionate tall stature, upper to lower segment ratio less than 0.85
C1861719|Mean full term birth length 55.2cm
C1861721|Adult height often normal
C1861723|Mean female adult height 172.9cm
C1839692|Adult height 120-150cm
C1839712|Short stature (3rd-10th percentile)
C1863421|Mean female height, 124 cm
C1857182|Adult height 98-127 cm
C1857200|Average birth length 44cm
C1851416|Short stature in less than 50%
C1867106|Average adult male height, 149.5 cm
C1837662|Length <3rd percentile by 6 months
C1837663|Adult height 110-130cm
C1842150|Short stature, proportionate (<5th percentile)
C1861137|Short stature (20% of adults)
C1866225|Postnatal deceleration of length
C1854707|Adult male height 136-161 cm
C1867488|Adult height, 82-130 cm
C1848504|Increased prenatal/postnatal length
C1846061|Short-trunk dwarfism, identifiable in infancy
C1846061|Infancy onset short-trunk short stature
C1855609|Stature below 25th percentile
C1833774|Normal to near normal stature
C1839811|Short to normal stature
C1860105|Severe short-limb dwarfism
C1834731|Short stature (3rd-25th percentile)
C1844832|Short stature (<5-15th percentile)
C1855748|Adult female height 107-143 cm
C1856085|Normal to tall stature
C1849526|Short stature from birth
C1867107|Average female adult height, 138 cm
C0521527|Short trunk
C0521527|Shortened appearance of trunk
C0521527|Shortened trunk
C0521527|Shortened trunk (disorder)
C1867869|Mean adult male height, 155 cm
C1867872|Fall-off in adolescent growth
C1849936|Adult female height 128-151cm
C0878659|Short stature, disproportionate
C0878659|Disproportionate short stature
C1832113|Short stature (<5th-10th percentile)
C1835109|Mean length at birth 53 +/- 4.4 cm for males
C1835110|Mean length at birth 52.5 +/- 3.5 cm for females
C1848489|Normal adult height
C1835580|Postnatal onset of mild growth retardation
C1835580|Mild postnatal growth retardation
C1856467|Normal upper/lower segment ratio
C1863393|Deceleration of linear growth during childhood
C1856919|Short stature (3rd-90th centile, infrequent finding)
C1860172|Average adult female height, 99.5cm
C1855747|Adult male height 136-157 cm
C1851728|Average birth length, 52.6cm
C1849264|Gigantism, mild-moderate
C1867124|Average adult male height 153 cm
C1839249|Final adult height 131-156 cm
C1839271|Birth length greater than 97th percentile
C1834991|Severe short stature, postnatal onset
C1834992|Average adult height 125cm
C1849935|Adult male height 141-155cm
C1842216|Adult female height 130-157 cm
C1848098|Severe short-trunked dwarfism (identifiable in early childhood)
C1835112|Mean adult height 175.4 +/- 8.2 cm for females
C1835114|Arm span to height > 1.05
C1848183|Tall for females (mean height 171.5cm)
C1861722|Mean male adult height 184.3cm
C1848394|Birth length > 90th percentile
C1855764|Below the third percentile
C1863345|Brachymelic dwarfism (upper limbs greater than lower limbs)
C1866694|Adult height 130-150 cm
C1854923|Deceleration of linear growth during first year
C1834760|Height >90th percentile
C1832445|Short stature (5th-10th percentile)
C1855200|Specific growth curves are available
C1855060|Short stature, most below 3rd percentile for height
C1855189|Short stature, disproportionate (short lower limbs)
C1855199|Weak or absent pubertal growth spurt
C1849535|Adult height less than 150 cm
C1867870|Mean adult female height, 147 cm
C1968810|Height less than 5th percentile
C1836996|Reduced upper-lower segment ratio
C1836996|Marfanoid habitus
C1836996|Marfanoid body habitus
C1836996|Reduced upper to lower segment ratio
C1836996|Disproportionate tall stature
C1969400|Stature (<10th percentile)
C1970082|Decreased height compared to unaffected siblings
C1970823|Tall, thin habitus
C0456070|Delayed growth
C0456070|Growth deficiency
C0456070|Delayed;growth
C0456070|Growth delay
C0456070|Growth delay (disorder)
C1970694|Normal stature (+1 SD to +2 SD)
C0015934|Fetal Growth Retardation
C0015934|Growth Retardation, Fetal
C0015934|Retardation, Fetal Growth
C0015934|Retardation, Intrauterine Growth
C0015934|intrauterine growth retardation
C0015934|Slow fetal growth, unspecified
C0015934|prenatal growth disorder
C0015934|Fetal growth restriction
C0015934|Intrauterine growth retardation (IUGR)
C0015934|intrauterine growth retardation (diagnosis)
C0015934|Intrauterine growth restriction
C0015934|Fet growth retard wtNOS
C0015934|IUGR
C0015934|Fetal Growth Retardation [Disease/Finding]
C0015934|Growth Retardation, Intrauterine
C0015934|Foetal growth restriction
C0015934|Microsomia
C0015934|Fetal growth retardation, unspecified, unspecified [weight]
C0015934|Fetal growth retardation, unspecified [weight]
C0015934|Poor prenatal growth
C0015934|(Fetal growth retardation NOS) or (intrauterine growth retardation)
C0015934|Insufficiency - placental
C0015934|(Fetal growth retardation NOS) or (intrauterine growth retardation) (disorder)
C0015934|Intrauterine growth retardatn.
C0015934|Fetal growth retardation NOS
C0015934|Fetal growth retardation NOS (disorder)
C0015934|Poor foetal growth state
C0015934|FGR - Foetal growth retardation
C0015934|Poor foetal growth
C0015934|Foetal growth retardation
C0015934|Intrauterine growth retardation (IUGR
C0015934|Foetal growth retardation, unspecified {weight}
C0015934|Fetal growth retardation, unspecified
C0015934|Growth intrauterine retard
C0015934|Foetal growth retardation, unspecified
C0015934|Fetal growth retardation, unspecified {weight}
C0015934|Intrauterine growth retard
C0015934|Poor fetal growth state
C0015934|Microsomic baby
C0015934|IUGR - Intrauterine growth retardation
C0015934|Poor fetal growth
C0015934|FGR - Fetal growth retardation
C0015934|Fetal growth retardation (disorder)
C0015934|fetal; growth retardation
C0015934|fetal; poor growth
C0015934|fetal; slow growth
C0015934|poor; fetal growth
C0015934|slow; fetal growth
C0015934|Fetal growth retardation, NOS
C0015934|Intrauterine growth retardation, NOS
C0015934|Foetal growth retardation, NOS
C0015934|Fetal growth retardation, unspecified weight
C0015934|Intrauterine growth retardatio
C1968917|Adult height (<100cm)
C0151686|Growth retardation
C0151686|Retarded growth
C0151686|Growth retardation (disorder)
C0151686|Retardation;growth
C0151686|Growth suppression
C0151686|Growth retarded
C0151686|Decreased growth
C0151686|Growth retardation (morphologic abnormality)
C0151686|growth; retardation
C0151686|retardation; growth
C0151686|Decreased growth, NOS
C0151686|Growth retardation, NOS
C0151686|Growth suppression, NOS
C1970743|Relative short stature (compared to unaffected males in family)
C1855652|Intrauterine growth failure
C1855652|Prenatal onset growth retardation
C1855652|Prenatal growth retardation
C1855652|Prenatal growth deficiency
C1855652|Prenatal-onset growth retardation
C1855652|Prenatal growth failure
C1855652|Fetus Small for Gestational Age
C1855652|Fetal SGA
C1855652|Fetal Small for Gestational Age
C1855652|Fetal Growth Restriction
C1855652|Intrauterine Growth Restriction
C1855652|IUGR
C1855652|In utero growth retardation
C1855652|Intrauterine growth retardation
C1855652|Intrauterine growth retardation (IUGR)
C1855652|Intrauterine growth retardation, IUGR
C0221097|Total Body Length
C0221097|Body Length
C0221097|BODLNGTH
C0221097|Length of body
C0221097|Length of body (observable entity)
C0005890|Body Height
C0005890|Body Heights
C0005890|Height, Body
C0005890|Heights, Body
C0005890|Stature
C0005890|Body height measure (observable entity)
C0005890|Body height measure
C0005890|Body height, NOS
C0005890|Body length
C0005890|Body length, NOS
C0005890|Height (Body)
C0242789|Crown Rump Length
C0242789|Crown-Rump Length
C0242789|Crown-Rump Lengths
C0242789|Length, Crown-Rump
C0242789|Lengths, Crown-Rump
C0242789|Length.crown rump
C0242789|CRL - Crown rump length
C0242789|Crown rump length (observable entity)
C0424648|Height from demispan
C0424648|Height from demispan (observable entity)
C0424647|Pubis to ground height
C0424647|Pubis to ground height (observable entity)
C0455805|Subischial leg length
C0455805|Subischial leg length (observable entity)
C1827986|Method for measuring height
C1827986|Method for measuring height (observable entity)
C0487985|Body height:Length:Point in time:^Patient:Quantitative
C0487985|Body height
C0487985|Body height:Len:Pt:^Patient:Qn
C0424651|Growth velocity centile
C0424651|Growth velocity centile (observable entity)
C0424649|Height centile
C0424649|Length centile
C0424649|Height centile (observable entity)
C0419485|Child height centiles
C0419485|Height centiles - child
C0419485|Child height centiles NOS
C0419485|Child height centiles NOS (finding)
C0419485|Child height centiles NOS (observable entity)
C0419485|Child height centile (observable entity)
C0419485|Child height centile
C1156245|Growth pattern (observable entity)
C1156245|Growth pattern
C0424638|Height and weight
C0424638|Height and Weight (observable entity)
C0424638|Height & weight
