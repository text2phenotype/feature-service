C0205177|T169|Active|
C0205177|T169|Active (qualifier value)|
C1446392|T033|Problem resolved (finding)|
C1446392|T033|Problem resolved|
C0277786|T033|Complaint|
C0277786|T033|Complaint (finding)|
C0205177|T169|Active|
C0205177|T169|Active (qualifier value)|
C0001779|T032|Age, function|
C0001779|T032|Age (observable entity)|
C0001779|T032|Age|
C0001779|T032|Has age|
C0001779|T032|Age, function (observable entity)|
C0012634|T047|Diseases|
C0012634|T047|Disease|
C0039082|T047|Syndrome|
C0012634|T047|Disorders|
C0012634|T047|Clinical disease AND/OR syndrome present|
C0012634|T047|Clinical disease AND/OR syndrome|
C0012634|T047|Disease (disorder)|
C0012634|T047|Disease AND/OR syndrome present|
C0012634|T047|Disorder|
C0012634|T047|Clinical disease or syndrome present, NOS|
C0012634|T047|Clinical disease or syndrome, NOS|
C0012634|T047|Disease or syndrome present, NOS|
C0012634|T047|Disease, NOS|
C0012634|T047|Disorder, NOS|
C0039082|T047|Syndrome, NOS|
C3495595|T203|Acetaminophen 325mg, Dextromethorphan Hydrobromide 10mg, Phenylephrine Hydrochloride 5mg Oral capsule, liquid filled, Acetaminophen 325mg, Dextromethorphan Hydrobromide 15mg, Doxylamine Succinate 6.25mg Oral capsule, liquid filled|
C2061888|T033|echocardiogram Pap muscles mitral transected posteromedial|
C2061888|T033|echocardiography: posteromedial mitral papillary muscles transected|
C2061888|T033|echocardiography: posteromedial mitral papillary muscles transected (procedure)|
C2935436|T116|ado-trastuzumab emtansine|
C2935436|T129|ado-trastuzumab emtansine|
C2935436|T121|ado-trastuzumab emtansine|
C1093123|T007|Streptomyces tenjimariensis|