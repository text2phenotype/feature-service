C0003873|Rheumatoid Arthritis
C1306838|Proliferative arthritis
C0003873|Rheumatoid arthritis
C0157913|Rheumatoid arthritis and other inflammatory polyarthropathies
C0015773|Feltys syndrome
C0015773|Feltys syndrome, unspecified site
C0015773|Rheumatoid arthritis with splenoadenomegaly and leukopenia
C0162323|Inflammatory polyarthropathies
C0162323|Inflammatory polyarthropathies (M05-M14)
C0240903|Rheumatoid vasculitis
C0264747|Rheumatoid pericarditis
C0392469|Rheumatoid carditis
C0409651|Seropositive rheumatoid arthritis
C0409651|Seropositive rheumatoid arthritis, unspecified
C0477541|Other seropositive rheumatoid arthritis
C0489959|Rheumatoid myocarditis
C0494896|Rheumatoid arthritis with involvement of other organs and systems
C0837507|Feltys syndrome, multiple sites
C0837511|Feltys syndrome, hand
C0837511|Feltys syndrome, unspecified hand
C0837514|Feltys syndrome, ankle and foot
C0837537|Rheu arthritis mult site w involv of organs and systems
C0837537|Rheumatoid arthritis of multiple sites with involvement of other organs and systems
C0837541|Rheumatoid arthritis of hand with involvement of other organs and systems
C0837544|Rheumatoid arthritis of ankle and foot with involvement of other organs and systems
C0837546|Rheu arthritis of unsp site w involv of organs and systems
C0837546|Rheumatoid arthritis of unspecified site with involvement of other organs and systems
C0994344|Rheumatoid lung disease
C2889108|Feltys syndrome, right shoulder
C2889109|Feltys syndrome, left shoulder
C2889110|Feltys syndrome, unspecified shoulder
C2889112|Feltys syndrome, right elbow
C2889113|Feltys syndrome, left elbow
C2889114|Feltys syndrome, carpal bones
C2889116|Feltys syndrome, right wrist
C2889117|Feltys syndrome, left wrist
C2889118|Feltys syndrome, unspecified wrist
C2889119|Feltys syndrome, metacarpus and phalanges
C2889120|Feltys syndrome, right hand
C2889121|Feltys syndrome, left hand
C2889122|Feltys syndrome, right hip
C2889123|Feltys syndrome, left hip
C2889126|Feltys syndrome, right knee
C2889127|Feltys syndrome, left knee
C2889128|Feltys syndrome, tarsus, metatarsus and phalanges
C2889129|Feltys syndrome, right ankle and foot
C2889130|Feltys syndrome, left ankle and foot
C2889131|Feltys syndrome, unspecified ankle and foot
C2889132|Rheumatoid lung disease with rheumatoid arthritis
C2889133|Rheumatoid lung disease w rheumatoid arthritis of unsp site
C2889133|Rheumatoid lung disease with rheumatoid arthritis of unspecified site
C2889134|Rheumatoid lung disease with rheumatoid arthritis of shoulder
C2889135|Rheumatoid lung disease w rheumatoid arthritis of r shoulder
C2889135|Rheumatoid lung disease with rheumatoid arthritis of right shoulder
C2889136|Rheumatoid lung disease w rheumatoid arthritis of l shoulder
C2889136|Rheumatoid lung disease with rheumatoid arthritis of left shoulder
C2889137|Rheu lung disease w rheumatoid arthritis of unsp shoulder
C2889137|Rheumatoid lung disease with rheumatoid arthritis of unspecified shoulder
C2889138|Rheumatoid lung disease with rheumatoid arthritis of elbow
C2889139|Rheumatoid lung disease w rheumatoid arthritis of r elbow
C2889139|Rheumatoid lung disease with rheumatoid arthritis of right elbow
C2889140|Rheumatoid lung disease w rheumatoid arthritis of left elbow
C2889140|Rheumatoid lung disease with rheumatoid arthritis of left elbow
C2889141|Rheumatoid lung disease w rheumatoid arthritis of unsp elbow
C2889141|Rheumatoid lung disease with rheumatoid arthritis of unspecified elbow
C2889142|Rheumatoid lung disease with rheumatoid arthritis, carpal bones
C2889143|Rheumatoid lung disease with rheumatoid arthritis of wrist
C2889144|Rheumatoid lung disease w rheumatoid arthritis of r wrist
C2889144|Rheumatoid lung disease with rheumatoid arthritis of right wrist
C2889145|Rheumatoid lung disease w rheumatoid arthritis of left wrist
C2889145|Rheumatoid lung disease with rheumatoid arthritis of left wrist
C2889146|Rheumatoid lung disease w rheumatoid arthritis of unsp wrist
C2889146|Rheumatoid lung disease with rheumatoid arthritis of unspecified wrist
C2889147|Rheumatoid lung disease with rheumatoid arthritis, metacarpus and phalanges
C2889148|Rheumatoid lung disease with rheumatoid arthritis of hand
C2889149|Rheumatoid lung disease w rheumatoid arthritis of right hand
C2889149|Rheumatoid lung disease with rheumatoid arthritis of right hand
C2889150|Rheumatoid lung disease w rheumatoid arthritis of left hand
C2889150|Rheumatoid lung disease with rheumatoid arthritis of left hand
C2889151|Rheumatoid lung disease w rheumatoid arthritis of unsp hand
C2889151|Rheumatoid lung disease with rheumatoid arthritis of unspecified hand
C2889152|Rheumatoid lung disease w rheumatoid arthritis of unsp hip
C2889152|Rheumatoid lung disease with rheumatoid arthritis of hip
C2889152|Rheumatoid lung disease with rheumatoid arthritis of unspecified hip
C2889153|Rheumatoid lung disease w rheumatoid arthritis of right hip
C2889153|Rheumatoid lung disease with rheumatoid arthritis of right hip
C2889154|Rheumatoid lung disease w rheumatoid arthritis of left hip
C2889154|Rheumatoid lung disease with rheumatoid arthritis of left hip
C2889155|Rheumatoid lung disease with rheumatoid arthritis of knee
C2889156|Rheumatoid lung disease w rheumatoid arthritis of right knee
C2889156|Rheumatoid lung disease with rheumatoid arthritis of right knee
C2889157|Rheumatoid lung disease w rheumatoid arthritis of left knee
C2889157|Rheumatoid lung disease with rheumatoid arthritis of left knee
C2889158|Rheumatoid lung disease w rheumatoid arthritis of unsp knee
C2889158|Rheumatoid lung disease with rheumatoid arthritis of unspecified knee
C2889159|Rheumatoid lung disease with rheumatoid arthritis, tarsus, metatarsus and phalanges
C2889160|Rheumatoid lung disease with rheumatoid arthritis of ankle and foot
C2889161|Rheu lung disease w rheumatoid arthritis of right ank/ft
C2889161|Rheumatoid lung disease with rheumatoid arthritis of right ankle and foot
C2889162|Rheu lung disease w rheumatoid arthritis of left ank/ft
C2889162|Rheumatoid lung disease with rheumatoid arthritis of left ankle and foot
C2889163|Rheu lung disease w rheumatoid arthritis of unsp ank/ft
C2889163|Rheumatoid lung disease with rheumatoid arthritis of unspecified ankle and foot
C2889164|Rheumatoid lung disease w rheumatoid arthritis mult site
C2889164|Rheumatoid lung disease with rheumatoid arthritis of multiple sites
C2889165|Rheumatoid vasculitis with rheumatoid arthritis
C2889165|Rheumatoid vasculitis with rheumatoid arthritis of unsp site
C2889165|Rheumatoid vasculitis with rheumatoid arthritis of unspecified site
C2889166|Rheumatoid vasculitis w rheumatoid arthritis of r shoulder
C2889166|Rheumatoid vasculitis with rheumatoid arthritis of right shoulder
C2889167|Rheumatoid vasculitis w rheumatoid arthritis of l shoulder
C2889167|Rheumatoid vasculitis with rheumatoid arthritis of left shoulder
C2889168|Rheu vasculitis w rheumatoid arthritis of unsp shoulder
C2889168|Rheumatoid vasculitis with rheumatoid arthritis of shoulder
C2889168|Rheumatoid vasculitis with rheumatoid arthritis of unspecified shoulder
C2889169|Rheumatoid vasculitis with rheumatoid arthritis of elbow
C2889170|Rheumatoid vasculitis w rheumatoid arthritis of right elbow
C2889170|Rheumatoid vasculitis with rheumatoid arthritis of right elbow
C2889171|Rheumatoid vasculitis w rheumatoid arthritis of left elbow
C2889171|Rheumatoid vasculitis with rheumatoid arthritis of left elbow
C2889172|Rheumatoid vasculitis w rheumatoid arthritis of unsp elbow
C2889172|Rheumatoid vasculitis with rheumatoid arthritis of unspecified elbow
C2889173|Rheumatoid vasculitis with rheumatoid arthritis, carpal bones
C2889174|Rheumatoid vasculitis with rheumatoid arthritis of wrist
C2889175|Rheumatoid vasculitis w rheumatoid arthritis of right wrist
C2889175|Rheumatoid vasculitis with rheumatoid arthritis of right wrist
C2889176|Rheumatoid vasculitis w rheumatoid arthritis of left wrist
C2889176|Rheumatoid vasculitis with rheumatoid arthritis of left wrist
C2889177|Rheumatoid vasculitis w rheumatoid arthritis of unsp wrist
C2889177|Rheumatoid vasculitis with rheumatoid arthritis of unspecified wrist
C2889178|Rheumatoid vasculitis with rheumatoid arthritis, metacarpus and phalanges
C2889179|Rheumatoid vasculitis with rheumatoid arthritis of hand
C2889179|Rheumatoid vasculitis with rheumatoid arthritis of unsp hand
C2889179|Rheumatoid vasculitis with rheumatoid arthritis of unspecified hand
C2889180|Rheumatoid vasculitis w rheumatoid arthritis of right hand
C2889180|Rheumatoid vasculitis with rheumatoid arthritis of right hand
C2889181|Rheumatoid vasculitis with rheumatoid arthritis of left hand
C2889182|Rheumatoid vasculitis with rheumatoid arthritis of hip
C2889183|Rheumatoid vasculitis with rheumatoid arthritis of right hip
C2889184|Rheumatoid vasculitis with rheumatoid arthritis of left hip
C2889185|Rheumatoid vasculitis with rheumatoid arthritis of unsp hip
C2889185|Rheumatoid vasculitis with rheumatoid arthritis of unspecified hip
C2889186|Rheumatoid vasculitis with rheumatoid arthritis of knee
C2889187|Rheumatoid vasculitis w rheumatoid arthritis of right knee
C2889187|Rheumatoid vasculitis with rheumatoid arthritis of right knee
C2889188|Rheumatoid vasculitis with rheumatoid arthritis of left knee
C2889189|Rheumatoid vasculitis with rheumatoid arthritis of unsp knee
C2889189|Rheumatoid vasculitis with rheumatoid arthritis of unspecified knee
C2889190|Rheumatoid vasculitis with rheumatoid arthritis, tarsus, metatarsus and phalanges
C2889191|Rheumatoid vasculitis with rheumatoid arthritis of ankle and foot
C2889192|Rheumatoid vasculitis w rheumatoid arthritis of right ank/ft
C2889192|Rheumatoid vasculitis with rheumatoid arthritis of right ankle and foot
C2889193|Rheumatoid vasculitis w rheumatoid arthritis of left ank/ft
C2889193|Rheumatoid vasculitis with rheumatoid arthritis of left ankle and foot
C2889194|Rheumatoid vasculitis w rheumatoid arthritis of unsp ank/ft
C2889194|Rheumatoid vasculitis with rheumatoid arthritis of unspecified ankle and foot
C2889195|Rheumatoid vasculitis w rheumatoid arthritis mult site
C2889195|Rheumatoid vasculitis with rheumatoid arthritis of multiple sites
C2889196|Rheumatoid endocarditis
C2889197|Rheumatoid heart disease with rheumatoid arthritis
C2889198|Rheumatoid heart disease w rheumatoid arthritis of unsp site
C2889198|Rheumatoid heart disease with rheumatoid arthritis of unspecified site
C2889199|Rheumatoid heart disease with rheumatoid arthritis of shoulder
C2889200|Rheu heart disease w rheumatoid arthritis of r shoulder
C2889200|Rheumatoid heart disease with rheumatoid arthritis of right shoulder
C2889201|Rheu heart disease w rheumatoid arthritis of l shoulder
C2889201|Rheumatoid heart disease with rheumatoid arthritis of left shoulder
C2889202|Rheu heart disease w rheumatoid arthritis of unsp shoulder
C2889202|Rheumatoid heart disease with rheumatoid arthritis of unspecified shoulder
C2889203|Rheumatoid heart disease with rheumatoid arthritis of elbow
C2889204|Rheumatoid heart disease w rheumatoid arthritis of r elbow
C2889204|Rheumatoid heart disease with rheumatoid arthritis of right elbow
C2889205|Rheumatoid heart disease w rheumatoid arthritis of l elbow
C2889205|Rheumatoid heart disease with rheumatoid arthritis of left elbow
C2889206|Rheu heart disease w rheumatoid arthritis of unsp elbow
C2889206|Rheumatoid heart disease with rheumatoid arthritis of unspecified elbow
C2889207|Rheumatoid heart disease with rheumatoid arthritis, carpal bones
C2889208|Rheumatoid heart disease with rheumatoid arthritis of wrist
C2889209|Rheumatoid heart disease w rheumatoid arthritis of r wrist
C2889209|Rheumatoid heart disease with rheumatoid arthritis of right wrist
C2889210|Rheumatoid heart disease w rheumatoid arthritis of l wrist
C2889210|Rheumatoid heart disease with rheumatoid arthritis of left wrist
C2889211|Rheu heart disease w rheumatoid arthritis of unsp wrist
C2889211|Rheumatoid heart disease with rheumatoid arthritis of unspecified wrist
C2889212|Rheumatoid heart disease with rheumatoid arthritis, metacarpus and phalanges
C2889213|Rheumatoid heart disease with rheumatoid arthritis of hand
C2889214|Rheu heart disease w rheumatoid arthritis of right hand
C2889214|Rheumatoid heart disease with rheumatoid arthritis of right hand
C2889215|Rheumatoid heart disease w rheumatoid arthritis of left hand
C2889215|Rheumatoid heart disease with rheumatoid arthritis of left hand
C2889216|Rheumatoid heart disease w rheumatoid arthritis of unsp hand
C2889216|Rheumatoid heart disease with rheumatoid arthritis of unspecified hand
C2889217|Rheumatoid heart disease w rheumatoid arthritis of unsp hip
C2889217|Rheumatoid heart disease with rheumatoid arthritis of hip
C2889217|Rheumatoid heart disease with rheumatoid arthritis of unspecified hip
C2889218|Rheumatoid heart disease w rheumatoid arthritis of right hip
C2889218|Rheumatoid heart disease with rheumatoid arthritis of right hip
C2889219|Rheumatoid heart disease w rheumatoid arthritis of left hip
C2889219|Rheumatoid heart disease with rheumatoid arthritis of left hip
C2889220|Rheumatoid heart disease with rheumatoid arthritis of knee
C2889221|Rheu heart disease w rheumatoid arthritis of right knee
C2889221|Rheumatoid heart disease with rheumatoid arthritis of right knee
C2889222|Rheumatoid heart disease w rheumatoid arthritis of left knee
C2889222|Rheumatoid heart disease with rheumatoid arthritis of left knee
C2889223|Rheumatoid heart disease w rheumatoid arthritis of unsp knee
C2889223|Rheumatoid heart disease with rheumatoid arthritis of unspecified knee
C2889224|Rheumatoid heart disease with rheumatoid arthritis, tarsus, metatarsus and phalanges
C2889225|Rheumatoid heart disease with rheumatoid arthritis of ankle and foot
C2889226|Rheu heart disease w rheumatoid arthritis of right ank/ft
C2889226|Rheumatoid heart disease with rheumatoid arthritis of right ankle and foot
C2889227|Rheu heart disease w rheumatoid arthritis of left ank/ft
C2889227|Rheumatoid heart disease with rheumatoid arthritis of left ankle and foot
C2889228|Rheu heart disease w rheumatoid arthritis of unsp ank/ft
C2889228|Rheumatoid heart disease with rheumatoid arthritis of unspecified ankle and foot
C2889229|Rheumatoid heart disease w rheumatoid arthritis mult site
C2889229|Rheumatoid heart disease with rheumatoid arthritis of multiple sites
C2889230|Rheumatoid myopathy with rheumatoid arthritis
C2889231|Rheumatoid myopathy with rheumatoid arthritis of unsp site
C2889231|Rheumatoid myopathy with rheumatoid arthritis of unspecified site
C2889232|Rheumatoid myopathy with rheumatoid arthritis of shoulder
C2889233|Rheumatoid myopathy w rheumatoid arthritis of right shoulder
C2889233|Rheumatoid myopathy with rheumatoid arthritis of right shoulder
C2889234|Rheumatoid myopathy w rheumatoid arthritis of left shoulder
C2889234|Rheumatoid myopathy with rheumatoid arthritis of left shoulder
C2889235|Rheumatoid myopathy w rheumatoid arthritis of unsp shoulder
C2889235|Rheumatoid myopathy with rheumatoid arthritis of unspecified shoulder
C2889236|Rheumatoid myopathy with rheumatoid arthritis of elbow
C2889237|Rheumatoid myopathy with rheumatoid arthritis of right elbow
C2889238|Rheumatoid myopathy with rheumatoid arthritis of left elbow
C2889239|Rheumatoid myopathy with rheumatoid arthritis of unsp elbow
C2889239|Rheumatoid myopathy with rheumatoid arthritis of unspecified elbow
C2889240|Rheumatoid myopathy with rheumatoid arthritis, carpal bones
C2889241|Rheumatoid myopathy with rheumatoid arthritis of wrist
C2889242|Rheumatoid myopathy with rheumatoid arthritis of right wrist
C2889243|Rheumatoid myopathy with rheumatoid arthritis of left wrist
C2889244|Rheumatoid myopathy with rheumatoid arthritis of unsp wrist
C2889244|Rheumatoid myopathy with rheumatoid arthritis of unspecified wrist
C2889245|Rheumatoid myopathy with rheumatoid arthritis, metacarpus and phalanges
C2889246|Rheumatoid myopathy with rheumatoid arthritis of hand
C2889246|Rheumatoid myopathy with rheumatoid arthritis of unsp hand
C2889246|Rheumatoid myopathy with rheumatoid arthritis of unspecified hand
C2889247|Rheumatoid myopathy with rheumatoid arthritis of right hand
C2889248|Rheumatoid myopathy with rheumatoid arthritis of left hand
C2889249|Rheumatoid myopathy with rheumatoid arthritis of hip
C2889250|Rheumatoid myopathy with rheumatoid arthritis of right hip
C2889251|Rheumatoid myopathy with rheumatoid arthritis of left hip
C2889252|Rheumatoid myopathy with rheumatoid arthritis of unsp hip
C2889252|Rheumatoid myopathy with rheumatoid arthritis of unspecified hip
C2889253|Rheumatoid myopathy with rheumatoid arthritis of knee
C2889254|Rheumatoid myopathy with rheumatoid arthritis of right knee
C2889255|Rheumatoid myopathy with rheumatoid arthritis of left knee
C2889256|Rheumatoid myopathy with rheumatoid arthritis of unsp knee
C2889256|Rheumatoid myopathy with rheumatoid arthritis of unspecified knee
C2889257|Rheumatoid myopathy with rheumatoid arthritis, tarsus, metatarsus and phalanges
C2889258|Rheumatoid myopathy with rheumatoid arthritis of ankle and foot
C2889259|Rheumatoid myopathy w rheumatoid arthritis of right ank/ft
C2889259|Rheumatoid myopathy with rheumatoid arthritis of right ankle and foot
C2889260|Rheumatoid myopathy w rheumatoid arthritis of left ank/ft
C2889260|Rheumatoid myopathy with rheumatoid arthritis of left ankle and foot
C2889261|Rheumatoid myopathy w rheumatoid arthritis of unsp ank/ft
C2889261|Rheumatoid myopathy with rheumatoid arthritis of unspecified ankle and foot
C2889262|Rheumatoid myopathy w rheumatoid arthritis of multiple sites
C2889262|Rheumatoid myopathy with rheumatoid arthritis of multiple sites
C2889263|Rheumatoid polyneuropathy with rheumatoid arthritis
C2889264|Rheumatoid polyneurop w rheumatoid arthritis of unsp site
C2889264|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified site
C2889265|Rheumatoid polyneuropathy with rheumatoid arthritis of shoulder
C2889266|Rheumatoid polyneurop w rheumatoid arthritis of r shoulder
C2889266|Rheumatoid polyneuropathy with rheumatoid arthritis of right shoulder
C2889267|Rheumatoid polyneurop w rheumatoid arthritis of l shoulder
C2889267|Rheumatoid polyneuropathy with rheumatoid arthritis of left shoulder
C2889268|Rheu polyneurop w rheumatoid arthritis of unsp shoulder
C2889268|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified shoulder
C2889269|Rheumatoid polyneurop w rheumatoid arthritis of right elbow
C2889269|Rheumatoid polyneuropathy with rheumatoid arthritis of right elbow
C2889270|Rheumatoid polyneurop w rheumatoid arthritis of left elbow
C2889270|Rheumatoid polyneuropathy with rheumatoid arthritis of left elbow
C2889271|Rheumatoid polyneurop w rheumatoid arthritis of unsp elbow
C2889271|Rheumatoid polyneuropathy with rheumatoid arthritis of elbow
C2889271|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified elbow
C2889272|Rheumatoid polyneuropathy with rheumatoid arthritis, carpal bones
C2889273|Rheumatoid polyneuropathy with rheumatoid arthritis of wrist
C2889274|Rheumatoid polyneurop w rheumatoid arthritis of right wrist
C2889274|Rheumatoid polyneuropathy with rheumatoid arthritis of right wrist
C2889275|Rheumatoid polyneurop w rheumatoid arthritis of left wrist
C2889275|Rheumatoid polyneuropathy with rheumatoid arthritis of left wrist
C2889276|Rheumatoid polyneurop w rheumatoid arthritis of unsp wrist
C2889276|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified wrist
C2889277|Rheumatoid polyneuropathy with rheumatoid arthritis, metacarpus and phalanges
C2889278|Rheumatoid polyneuropathy with rheumatoid arthritis of hand
C2889279|Rheumatoid polyneurop w rheumatoid arthritis of right hand
C2889279|Rheumatoid polyneuropathy with rheumatoid arthritis of right hand
C2889280|Rheumatoid polyneurop w rheumatoid arthritis of left hand
C2889280|Rheumatoid polyneuropathy with rheumatoid arthritis of left hand
C2889281|Rheumatoid polyneurop w rheumatoid arthritis of unsp hand
C2889281|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified hand
C2889282|Rheumatoid polyneuropathy with rheumatoid arthritis of hip
C2889283|Rheumatoid polyneurop w rheumatoid arthritis of right hip
C2889283|Rheumatoid polyneuropathy with rheumatoid arthritis of right hip
C2889284|Rheumatoid polyneuropathy w rheumatoid arthritis of left hip
C2889284|Rheumatoid polyneuropathy with rheumatoid arthritis of left hip
C2889285|Rheumatoid polyneuropathy w rheumatoid arthritis of unsp hip
C2889285|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified hip
C2889286|Rheumatoid polyneuropathy with rheumatoid arthritis of knee
C2889287|Rheumatoid polyneurop w rheumatoid arthritis of right knee
C2889287|Rheumatoid polyneuropathy with rheumatoid arthritis of right knee
C2889288|Rheumatoid polyneurop w rheumatoid arthritis of left knee
C2889288|Rheumatoid polyneuropathy with rheumatoid arthritis of left knee
C2889289|Rheumatoid polyneurop w rheumatoid arthritis of unsp knee
C2889289|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified knee
C2889290|Rheumatoid polyneuropathy with rheumatoid arthritis, tarsus, metatarsus and phalanges
C2889291|Rheumatoid polyneuropathy with rheumatoid arthritis of ankle and foot
C2889292|Rheumatoid polyneurop w rheumatoid arthritis of right ank/ft
C2889292|Rheumatoid polyneuropathy with rheumatoid arthritis of right ankle and foot
C2889293|Rheumatoid polyneurop w rheumatoid arthritis of left ank/ft
C2889293|Rheumatoid polyneuropathy with rheumatoid arthritis of left ankle and foot
C2889294|Rheumatoid polyneurop w rheumatoid arthritis of unsp ank/ft
C2889294|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified ankle and foot
C2889295|Rheumatoid polyneuropathy w rheumatoid arthritis mult site
C2889295|Rheumatoid polyneuropathy with rheumatoid arthritis of multiple sites
C2889296|Rheumatoid arthritis of shoulder with involvement of other organs and systems
C2889297|Rheu arthritis of r shoulder w involv of organs and systems
C2889297|Rheumatoid arthritis of right shoulder with involvement of other organs and systems
C2889298|Rheu arthritis of l shoulder w involv of organs and systems
C2889298|Rheumatoid arthritis of left shoulder with involvement of other organs and systems
C2889299|Rheu arthrit of unsp shoulder w involv of organs and systems
C2889299|Rheumatoid arthritis of unspecified shoulder with involvement of other organs and systems
C2889300|Rheumatoid arthritis of elbow with involvement of other organs and systems
C2889301|Rheu arthritis of r elbow w involv of organs and systems
C2889301|Rheumatoid arthritis of right elbow with involvement of other organs and systems
C2889302|Rheu arthritis of l elbow w involv of organs and systems
C2889302|Rheumatoid arthritis of left elbow with involvement of other organs and systems
C2889303|Rheu arthritis of unsp elbow w involv of organs and systems
C2889303|Rheumatoid arthritis of unspecified elbow with involvement of other organs and systems
C2889304|Rheumatoid arthritis of carpal bones with involvement of other organs and systems
C2889305|Rheumatoid arthritis of wrist with involvement of other organs and systems
C2889306|Rheu arthritis of r wrist w involv of organs and systems
C2889306|Rheumatoid arthritis of right wrist with involvement of other organs and systems
C2889307|Rheu arthritis of l wrist w involv of organs and systems
C2889307|Rheumatoid arthritis of left wrist with involvement of other organs and systems
C2889308|Rheu arthritis of unsp wrist w involv of organs and systems
C2889308|Rheumatoid arthritis of unspecified wrist with involvement of other organs and systems
C2889309|Rheumatoid arthritis of metacarpus and phalanges with involvement of other organs and systems
C2889310|Rheu arthritis of right hand w involv of organs and systems
C2889310|Rheumatoid arthritis of right hand with involvement of other organs and systems
C2889311|Rheu arthritis of left hand w involv of organs and systems
C2889311|Rheumatoid arthritis of left hand with involvement of other organs and systems
C2889312|Rheu arthritis of unsp hand w involv of organs and systems
C2889312|Rheumatoid arthritis of unspecified hand with involvement of other organs and systems
C2889313|Rheumatoid arthritis of hip with involvement of other organs and systems
C2889314|Rheu arthritis of right hip w involv of organs and systems
C2889314|Rheumatoid arthritis of right hip with involvement of other organs and systems
C2889315|Rheu arthritis of left hip w involv of organs and systems
C2889315|Rheumatoid arthritis of left hip with involvement of other organs and systems
C2889316|Rheu arthritis of unsp hip w involv of organs and systems
C2889316|Rheumatoid arthritis of unspecified hip with involvement of other organs and systems
C2889317|Rheumatoid arthritis of knee with involvement of other organs and systems
C2889318|Rheu arthritis of right knee w involv of organs and systems
C2889318|Rheumatoid arthritis of right knee with involvement of other organs and systems
C2889319|Rheu arthritis of left knee w involv of organs and systems
C2889319|Rheumatoid arthritis of left knee with involvement of other organs and systems
C2889320|Rheu arthritis of unsp knee w involv of organs and systems
C2889320|Rheumatoid arthritis of unspecified knee with involvement of other organs and systems
C2889321|Rheumatoid arthritis of tarsus, metatarsus and phalanges with involvement of other organs and systems
C2889322|Rheu arthrit of right ank/ft w involv of organs and systems
C2889322|Rheumatoid arthritis of right ankle and foot with involvement of other organs and systems
C2889323|Rheu arthritis of left ank/ft w involv of organs and systems
C2889323|Rheumatoid arthritis of left ankle and foot with involvement of other organs and systems
C2889324|Rheu arthritis of unsp ank/ft w involv of organs and systems
C2889324|Rheumatoid arthritis of unspecified ankle and foot with involvement of other organs and systems
C2889325|Rheumatoid arthritis with rheumatoid factor without organ or systems involvement
C2889326|Rheu arthritis w rheu factor of unsp site w/o org/sys involv
C2889326|Rheumatoid arthritis with rheumatoid factor of unspecified site without organ or systems involvement
C2889327|Rheumatoid arthritis with rheumatoid factor of shoulder without organ or systems involvement
C2889328|Rheu arthrit w rheu factor of r shoulder w/o org/sys involv
C2889328|Rheumatoid arthritis with rheumatoid factor of right shoulder without organ or systems involvement
C2889329|Rheu arthrit w rheu factor of l shoulder w/o org/sys involv
C2889329|Rheumatoid arthritis with rheumatoid factor of left shoulder without organ or systems involvement
C2889330|Rheu arthrit w rheu factor of unsp shldr w/o org/sys involv
C2889330|Rheumatoid arthritis with rheumatoid factor of unspecified shoulder without organ or systems involvement
C2889331|Rheumatoid arthritis with rheumatoid factor of elbow without organ or systems involvement
C2889332|Rheu arthritis w rheu factor of r elbow w/o org/sys involv
C2889332|Rheumatoid arthritis with rheumatoid factor of right elbow without organ or systems involvement
C2889333|Rheu arthritis w rheu factor of l elbow w/o org/sys involv
C2889333|Rheumatoid arthritis with rheumatoid factor of left elbow without organ or systems involvement
C2889334|Rheu arthrit w rheu factor of unsp elbow w/o org/sys involv
C2889334|Rheumatoid arthritis with rheumatoid factor of unspecified elbow without organ or systems involvement
C2889335|Rheumatoid arthritis with rheumatoid factor of wrist without organ or systems involvement
C2889336|Rheu arthritis w rheu factor of r wrist w/o org/sys involv
C2889336|Rheumatoid arthritis with rheumatoid factor of right wrist without organ or systems involvement
C2889337|Rheu arthritis w rheu factor of l wrist w/o org/sys involv
C2889337|Rheumatoid arthritis with rheumatoid factor of left wrist without organ or systems involvement
C2889338|Rheu arthrit w rheu factor of unsp wrist w/o org/sys involv
C2889338|Rheumatoid arthritis with rheumatoid factor of unspecified wrist without organ or systems involvement
C2889339|Rheumatoid arthritis with rheumatoid factor of hand without organ or systems involvement
C2889340|Rheu arthritis w rheu factor of r hand w/o org/sys involv
C2889340|Rheumatoid arthritis with rheumatoid factor of right hand without organ or systems involvement
C2889341|Rheu arthritis w rheu factor of left hand w/o org/sys involv
C2889341|Rheumatoid arthritis with rheumatoid factor of left hand without organ or systems involvement
C2889342|Rheu arthritis w rheu factor of unsp hand w/o org/sys involv
C2889342|Rheumatoid arthritis with rheumatoid factor of unspecified hand without organ or systems involvement
C2889343|Rheumatoid arthritis with rheumatoid factor of hip without organ or systems involvement
C2889344|Rheu arthritis w rheu factor of right hip w/o org/sys involv
C2889344|Rheumatoid arthritis with rheumatoid factor of right hip without organ or systems involvement
C2889345|Rheu arthritis w rheu factor of left hip w/o org/sys involv
C2889345|Rheumatoid arthritis with rheumatoid factor of left hip without organ or systems involvement
C2889346|Rheu arthritis w rheu factor of unsp hip w/o org/sys involv
C2889346|Rheumatoid arthritis with rheumatoid factor of unspecified hip without organ or systems involvement
C2889347|Rheumatoid arthritis with rheumatoid factor of knee without organ or systems involvement
C2889348|Rheu arthritis w rheu factor of r knee w/o org/sys involv
C2889348|Rheumatoid arthritis with rheumatoid factor of right knee without organ or systems involvement
C2889349|Rheu arthritis w rheu factor of left knee w/o org/sys involv
C2889349|Rheumatoid arthritis with rheumatoid factor of left knee without organ or systems involvement
C2889350|Rheu arthritis w rheu factor of unsp knee w/o org/sys involv
C2889350|Rheumatoid arthritis with rheumatoid factor of unspecified knee without organ or systems involvement
C2889351|Rheumatoid arthritis with rheumatoid factor of ankle and foot without organ or systems involvement
C2889352|Rheu arthrit w rheu fctr of right ank/ft w/o org/sys involv
C2889352|Rheumatoid arthritis with rheumatoid factor of right ankle and foot without organ or systems involvement
C2889353|Rheu arthrit w rheu factor of left ank/ft w/o org/sys involv
C2889353|Rheumatoid arthritis with rheumatoid factor of left ankle and foot without organ or systems involvement
C2889354|Rheu arthrit w rheu factor of unsp ank/ft w/o org/sys involv
C2889354|Rheumatoid arthritis with rheumatoid factor of unspecified ankle and foot without organ or systems involvement
C2889355|Rheu arthritis w rheu factor mult site w/o org/sys involv
C2889355|Rheumatoid arthritis with rheumatoid factor of multiple sites without organ or systems involvement
C2889356|Oth rheumatoid arthritis with rheumatoid factor of unsp site
C2889356|Other rheumatoid arthritis with rheumatoid factor
C2889356|Other rheumatoid arthritis with rheumatoid factor of unspecified site
C2889357|Other rheumatoid arthritis with rheumatoid factor of shoulder
C2889358|Oth rheumatoid arthritis w rheumatoid factor of r shoulder
C2889358|Other rheumatoid arthritis with rheumatoid factor of right shoulder
C2889359|Oth rheumatoid arthritis w rheumatoid factor of l shoulder
C2889359|Other rheumatoid arthritis with rheumatoid factor of left shoulder
C2889360|Oth rheu arthritis w rheumatoid factor of unsp shoulder
C2889360|Other rheumatoid arthritis with rheumatoid factor of unspecified shoulder
C2889361|Other rheumatoid arthritis with rheumatoid factor of elbow
C2889362|Oth rheumatoid arthritis w rheumatoid factor of right elbow
C2889362|Other rheumatoid arthritis with rheumatoid factor of right elbow
C2889363|Oth rheumatoid arthritis w rheumatoid factor of left elbow
C2889363|Other rheumatoid arthritis with rheumatoid factor of left elbow
C2889364|Oth rheumatoid arthritis w rheumatoid factor of unsp elbow
C2889364|Other rheumatoid arthritis with rheumatoid factor of unspecified elbow
C2889365|Other rheumatoid arthritis with rheumatoid factor of wrist
C2889366|Oth rheumatoid arthritis w rheumatoid factor of right wrist
C2889366|Other rheumatoid arthritis with rheumatoid factor of right wrist
C2889367|Oth rheumatoid arthritis w rheumatoid factor of left wrist
C2889367|Other rheumatoid arthritis with rheumatoid factor of left wrist
C2889368|Oth rheumatoid arthritis w rheumatoid factor of unsp wrist
C2889368|Other rheumatoid arthritis with rheumatoid factor of unspecified wrist
C2889369|Oth rheumatoid arthritis w rheumatoid factor of right hand
C2889369|Other rheumatoid arthritis with rheumatoid factor of right hand
C2889370|Oth rheumatoid arthritis with rheumatoid factor of left hand
C2889370|Other rheumatoid arthritis with rheumatoid factor of left hand
C2889371|Oth rheumatoid arthritis with rheumatoid factor of unsp hand
C2889371|Other rheumatoid arthritis with rheumatoid factor of hand
C2889371|Other rheumatoid arthritis with rheumatoid factor of unspecified hand
C2889372|Other rheumatoid arthritis with rheumatoid factor of hip
C2889373|Oth rheumatoid arthritis with rheumatoid factor of right hip
C2889373|Other rheumatoid arthritis with rheumatoid factor of right hip
C2889374|Oth rheumatoid arthritis with rheumatoid factor of left hip
C2889374|Other rheumatoid arthritis with rheumatoid factor of left hip
C2889375|Oth rheumatoid arthritis with rheumatoid factor of unsp hip
C2889375|Other rheumatoid arthritis with rheumatoid factor of unspecified hip
C2889376|Other rheumatoid arthritis with rheumatoid factor of knee
C2889377|Oth rheumatoid arthritis w rheumatoid factor of right knee
C2889377|Other rheumatoid arthritis with rheumatoid factor of right knee
C2889378|Oth rheumatoid arthritis with rheumatoid factor of left knee
C2889378|Other rheumatoid arthritis with rheumatoid factor of left knee
C2889379|Oth rheumatoid arthritis with rheumatoid factor of unsp knee
C2889379|Other rheumatoid arthritis with rheumatoid factor of unspecified knee
C2889380|Other rheumatoid arthritis with rheumatoid factor of ankle and foot
C2889381|Oth rheumatoid arthritis w rheumatoid factor of right ank/ft
C2889381|Other rheumatoid arthritis with rheumatoid factor of right ankle and foot
C2889382|Oth rheumatoid arthritis w rheumatoid factor of left ank/ft
C2889382|Other rheumatoid arthritis with rheumatoid factor of left ankle and foot
C2889383|Oth rheumatoid arthritis w rheumatoid factor of unsp ank/ft
C2889383|Other rheumatoid arthritis with rheumatoid factor of unspecified ankle and foot
C2889384|Oth rheumatoid arthritis w rheumatoid factor mult site
C2889384|Other rheumatoid arthritis with rheumatoid factor of multiple sites
C2889385|Rheumatoid arthritis with rheumatoid factor
C2889385|Rheumatoid arthritis with rheumatoid factor, unspecified
C3469320|Feltys syndrome, elbow
C3469320|Feltys syndrome, unspecified elbow
C3469322|Feltys syndrome, hip
C3469322|Feltys syndrome, unspecified hip
C3469323|Feltys syndrome, knee
C3469323|Feltys syndrome, unspecified knee
C3469325|Feltys syndrome, shoulder
C3469326|Feltys syndrome, wrist
C3714757|juvenile rheumatoid arthritis
C3714757|Rheumatoid arthritis, juvenile
C3714757|Unspecified juvenile rheumatoid arthritis
C3714757|JRA
C3714757|Childhood arthritis
C3714757|Juvenile idiopathic arthritis
C3714757|Juvenile rheumatoid arthritis (disorder)
C3714757|JRA - Juvenile rheumatoid arthritis
C3714757|Juvenile rheumatoid arthritis NOS (disorder)
C3714757|Juvenile rheumatoid arthritis NOS
C3714757|Juvenile rheumatoid a.
C3714757|Juvenile seropositive arthritis
C3714757|Rheumatoid arthritis in children
C3714757|Juvenile RA
C3714757|Juvenile Arthritis
C3714757|Juvenile Rheumatoid Arthritis (AQ)
C3714757|juvenile idiopathic arthritis (diagnosis)
C3714757|juvenile; arthritis, rheumatoid
C3714757|arthritis; juvenile, rheumatoid
C3714757|arthritis; rheumatoid, juvenile
C3714757|Juvenile rheumatoid arthritis, NOS
C0038013|Ankylosing spondylitis
C0038013|Bechterews Disease
C0038013|Marie Struempell Disease
C0038013|Spondylitis, Ankylosing
C0038013|Spondylitis, Rheumatoid
C0038013|BECHTEREW DIS
C0038013|MARIE STRUEMPELL DIS
C0038013|BECHTEREWS DIS
C0038013|ankylosing spondylitis (diagnosis)
C0038013|Ank spond
C0038013|Spondyloarthritides, Ankylosing
C0038013|Ankylosing Spondyloarthritides
C0038013|Spondylarthritides, Ankylosing
C0038013|Spondylarthritis, Ankylosing
C0038013|Spondyloarthritis, Ankylosing
C0038013|Ankylosing Spondylarthritides
C0038013|Rheumatoid arthritis of spine
C0038013|Rheumatoid Spondylitis
C0038013|Spondylarthritis Ankylopoietica
C0038013|Bechterew's Disease
C0038013|Bechterew Disease
C0038013|Marie-Struempell Disease
C0038013|Spondylitis, Ankylosing [Disease/Finding]
C0038013|Ankylosing Spondylarthritis
C0038013|Ankylosing Spondyloarthritis
C0038013|Disease;Bechterews
C0038013|Ankylosing spondylitis (disorder)
C0038013|Spondylitis Ankylopoietica
C0038013|Spondyloarthritis Ankylopoietica
C0038013|Spondylitis ankylosing
C0038013|Bekhterev's disease
C0038013|AS - Ankylosing spondylitis
C0038013|Idiopathic ankylosing spondylitis
C0038013|Marie-Strumpell spondylitis
C0038013|Marie Strümpell spondylitis
C0038013|arthritis; spine or vertebra, Marie-Strümpell
C0038013|arthritis; spine or vertebra, ankylosing
C0038013|Marie-Strümpell; spondylitis
C0038013|Marie-Strümpell
C0038013|Strümpell-Marie
C0038013|Von Bechterew
C0038013|Bechterew
C0038013|rheumatoid; arthritis, spine
C0038013|rheumatoid; spondylitis
C0038013|spine or vertebra; arthritis, Marie-Strümpell
C0038013|spine or vertebra; arthritis, ankylosing
C0038013|spondylitis; Marie-Strümpell
C0038013|spondylitis; ankylopoietica
C0038013|spondylitis; ankylosing
C0038013|spondylitis; rheumatoid
C0038013|ankylopoietica; spondylitis
C0038013|ankylosing; spondylitis
C0038013|arthritis; rheumatoid, spine
C0038013|Ankylosing spondylitis, NOS
C0038013|Rheumatoid arthritis of spine, NOS
C0038013|Spondylitis, Marie-Strumpell
C0038013|Rheumatioid arthritis of spine NOS
C0409628|Other rheumatoid arthropathy with visceral or systemic involvement (disorder)
C0409628|Other rheumatoid arthropathy with visceral or systemic involvement
C0409629|Rheumatoid arthritis of interphalangeal joint of toe
C0409629|Rheumatoid arthritis of interphalangeal joint of toe (disorder)
C0409630|Rheumatoid arthritis of lesser metatarsophalangeal joint
C0409630|Rheumatoid arthritis of lesser metatarsophalangeal joint (disorder)
C0409631|Rheumatoid arthritis of 1st metatarsophalangeal joint
C0409631|Rheumatoid arthritis of first metatarsophalangeal joint
C0409631|Rheumatoid arthritis of first metatarsophalangeal joint (disorder)
C0409632|Rheumatoid arthritis of other tarsal joint
C0409632|Rheumatoid arthritis of other tarsal joint (disorder)
C0409633|Rheumatoid arthritis of talonavicular joint
C0409633|Rheumatoid arthritis of talonavicular joint (disorder)
C0409634|Rheumatoid arthritis of subtalar joint
C0409634|Rheumatoid arthritis of subtalar joint (disorder)
C0409635|rheumatoid arthritis of ankle (diagnosis)
C0409635|rheumatoid arthritis of ankle
C0409635|Rheumatoid arthritis of ankle (disorder)
C0409637|rheumatoid arthritis of knee
C0409637|rheumatoid arthritis of knee (diagnosis)
C0409637|Rheumatoid arthritis of knee (disorder)
C0409639|Rheumatoid arthritis of hip
C0409639|rheumatoid arthritis of hip (diagnosis)
C0409639|Rheumatoid arthritis of hip (disorder)
C0409640|Rheumatoid arthritis of distal interphalangeal joint of finger
C0409640|Rheumatoid arthritis of distal interphalangeal joint of finger (disorder)
C0409641|Rheumatoid arthritis of proximal interphalangeal joint of finger
C0409641|Rheumatoid arthritis of proximal interphalangeal joint of finger (disorder)
C0409642|Rheumatoid arthritis of metacarpophalangeal joint
C0409642|Rheumatoid arthritis of metacarpophalangeal joint (disorder)
C0409643|rheumatoid arthritis of wrist
C0409643|rheumatoid arthritis of wrist (diagnosis)
C0409643|Rheumatoid arthritis of wrist (disorder)
C0409645|rheumatoid arthritis of elbow (diagnosis)
C0409645|Rheumatoid arthritis of elbow
C0409645|Rheumatoid arthritis of elbow (disorder)
C0409646|Rheumatoid arthritis of acromioclavicular joint
C0409646|Rheumatoid arthritis of acromioclavicular joint (disorder)
C0409647|Rheumatoid arthritis of sternoclavicular joint
C0409647|Rheumatoid arthritis of sternoclavicular joint (disorder)
C0409648|rheumatoid arthritis shoulder (diagnosis)
C0409648|rheumatoid arthritis shoulder
C0409648|Rheumatoid arthritis of shoulder
C0409648|Rheumatoid arthritis of shoulder (disorder)
C0409650|Rheumatoid arthritis of cervical spine
C0409650|Rheumatoid arthritis of cervical spine (disorder)
C0409651|Seropositive rheumatoid arthritis
C0409651|Seropositive rheumatoid arthritis, unspecified
C0409651|rheumatoid factor positive (diagnosis)
C0409651|rheumatoid factor positive
C0409651|[X]Seropositive rheumatoid arthritis, unspecified (disorder)
C0409651|[X]Seropositive rheumatoid arthritis, unspecified
C0409651|Seropositive RA
C0409651|Seropositive rheumatoid arthritis (disorder)
C0409651|rheumatoid; arthritis, seropositive
C0409651|arthritis; rheumatoid, seropositive
C0409652|Seronegative rheumatoid arthritis
C0409652|Seronegative rheumatoid arthritis (disorder)
C0409652|rheumatoid; arthritis, seronegative
C0409652|arthritis; rheumatoid, seronegative
C0409657|Rheumatoid arthritis with multisystem involvement
C0409657|Rheumatoid arthritis with multisystem involvement (disorder)
C0856832|Monoarthritic rheumatoid arthritis
C0477541|Other seropositive rheumatoid arthritis
C0477541|[X]Other seropositive rheumatoid arthritis
C0477541|[X]Other seropositive rheumatoid arthritis (disorder)
C0494896|Rheumatoid arthritis with involvement of other organs and systems
C0494896|rheumatoid; arthritis, with systemic involvement
C0494896|arthritis; rheumatoid, with systemic involvement
C0235762|Arthritis rheumatoid aggravated
C0235762|Rheumatoid arthritis aggravated
C0837691|Juv rheum arthritis NOS
C0837691|Polyarticular juvenile rheumatoid arthritis, chronic or unspecified
C0837691|juvenile idiopathic arthritis of multiple sites
C0837691|juvenile idiopathic arthritis multiple sites
C0837691|juvenile idiopathic arthritis of multiple sites (diagnosis)
C0263737|Uveitis-rheumatoid arthritis syndrome
C0263737|Uveitis-rheumatoid arthritis syndrome (disorder)
C0157914|Other rheumatoid arthritis with visceral or systemic involvement
C0157914|Rheumatoid arthritis with other visceral or systemic involvement -RETIRED-
C0157914|Syst rheum arthritis NEC
C0157914|Rheumatoid arthritis with other visceral or systemic involvement (disorder)
C0157914|Rheumatoid arthritis with other visceral or systemic involvement
C0157917|Pauciarticular juvenile arthritis
C0157917|Oligoarticular Still Disease
C0157917|Oligoarticular Still's Disease
C0157917|Pauciart juv rheum arthr
C0157917|Pauciarticular juvenile rheumatoid arthritis
C0157917|Pauciarticular juvenile rheumatoid arthritis, unspecified site
C0157917|Pauciarticular juvenile rheumatoid arthritis, unsp site
C0157917|Pauciarticular onset juvenile chronic arthritis (disorder)
C0157917|Pauciarticular onset juvenile chronic arthritis
C0157917|Pauciarticular JRA
C0157917|Pauciarticular juvenile chronic RA
C0157917|Pauciarticular Juvenile Rheumatoid Arthritis (AQ)
C0157917|Oligoarticular JRA
C0157917|Oligoarticular Juvenile Rheumatoid Arthritis
C0157917|JCA - Pauciarticular onset juvenile chronic arthritis
C0157917|Pauciarticular onset juvenile arthritis
C0157917|Pauciarticular juvenile rheumatoid arthritis (disorder)
C0157917|juvenile; arthritis, pauciarticular
C0157917|arthritis; juvenile, pauciarticular
C0409636|Rheumatoid arthritis of tibiofibular joint
C0409636|Rheumatoid arthritis of tibiofibular joint (disorder)
C0409644|Rheumatoid arthritis of distal radioulnar joint
C0409644|Rheumatoid arthritis of distal radioulnar joint (disorder)
C0409638|Rheumatoid arthritis of sacroiliac joint
C0409638|Rheumatoid arthritis of sacroiliac joint (disorder)
C0006915|Caplans Syndrome
C0006915|Caplan's syndrome
C0006915|Caplan's syndrome (diagnosis)
C0006915|Caplan Syndrome
C0006915|Caplan Syndromes
C0006915|Caplan Syndrome [Disease/Finding]
C0006915|Rheumatoid pneumoconiosis (disorder)
C0006915|Rheumatoid pneumoconiosis
C0006915|Caplan (etiology)
C0006915|Caplan (manifestation)
C0015773|Feltys Syndrome
C0015773|Syndrome, Felty's
C0015773|Felty's syndrome
C0015773|FELTY SYNDROME
C0015773|Felty's syndrome (diagnosis)
C0015773|Rheumatoid arthritis with splenoadenomegaly and leukopenia
C0015773|Felty's syndrome, unspecified site
C0015773|Syndrome, Felty
C0015773|Felty Syndrome [Disease/Finding]
C0015773|Felty's syndrome (disorder)
C0015773|Rheumatoid arthritis, leucopenia AND splenomegaly
C0015773|Rheumatoid arthritis, leukopenia AND splenomegaly
C0015773|Felty
C0015773|rheumatoid; arthritis, with splenoadenomegaly and leukopenia
C0015773|arthritis; rheumatoid, with splenoadenomegaly and leukopenia
C0015773|Rheumatoid arthritis, leukopenia and splenadenomegaly
C0035450|Nodule, Rheumatoid
C0035450|Nodules, Rheumatoid
C0035450|Rheumatoid Nodule
C0035450|Rheumatoid Nodules
C0035450|RHEUMATOID NODULOSIS
C0035450|Rheumatoid Nodule [Disease/Finding]
C0035450|Rheumatoid Noduloses
C0035450|Rheumatoid nodule (disorder)
C0035450|Subcutaneous rheumatoid nodule
C0035450|Rheumatoid nodule (morphologic abnormality)
C0035450|Rheumatoid nodulosis (disorder)
C0035450|Subcutaneous rheumatoid nodule (disorder)
C0035450|node; rheumatoid
C0035450|nodule; rheumatoid
C0035450|rheumatoid; node
C0035450|rheumatoid; nodule
C0035450|Rheumatoid nodule, NOS
C1527336|Sjogren's Syndrome
C1527336|Syndrome, Sjogren's
C1527336|Sjogrens Syndrome
C1527336|Sicca syndrome [Sjogren]
C1527336|Sjogren's disease
C1527336|SJOGREN SYNDROME
C1527336|Sjogren's Syndrome [Disease/Finding]
C1527336|Sicca (Sjogren's) syndrome
C1527336|Sjogren syndrome (diagnosis)
C1527336|Sjogren's
C1527336|Gougerot-Mulock-Houwer syndrome
C1527336|Syndrome Sjogren's
C1527336|Sjoegren's syndrome
C1527336|Sjögren's syndrome (disorder)
C1527336|Sjögren
C0085253|Adult Onset Still Disease
C0085253|Adult Onset Still's Disease
C0085253|Adult-Onset Stills Disease
C0085253|Still Disease, Adult Onset
C0085253|Still's Disease, Adult Onset
C0085253|Still's Disease, Adult-Onset
C0085253|Stills Disease, Adult-Onset
C0085253|Adult-onset Still's disease
C0085253|Adult-Onset Still Disease
C0085253|ADULT ONSET STILL DIS
C0085253|STILLS DIS ADULT ONSET
C0085253|ADULT ONSET STILLS DIS
C0085253|STILL DIS ADULT ONSET
C0085253|Still's disease adult onset
C0085253|adult onset Still's disease (diagnosis)
C0085253|AOSD (adult onset Still's disease)
C0085253|adult Still's disease
C0085253|Still's Disease, Adult-Onset [Disease/Finding]
C0085253|Still Disease, Adult-Onset
C0085253|Adult onset Still's disease (disorder)
C0085253|disease; Still's adult onset
C0085253|Still's adult onset; disease
C0085253|Still; adult-onset
C0085253|adult-onset; Still
C0003873|Rheumatoid arthritis
C0003873|Arthritis, Rheumatoid
C0003873|Rheumatoid arthritis, unspecified
C0003873|RA
C0003873|RA (rheumatoid arthritis)
C0003873|rheumatoid arthritis (diagnosis)
C0003873|R arthritis
C0003873|Rh arthritis
C0003873|Arthritis, Rheumatoid [Disease/Finding]
C0003873|Rheumatoid arthritis NOS (disorder)
C0003873|Rheumatoid arthritis NOS
C0003873|Rheumatoid arthritis (disorder)
C0003873|Arthritis rheumatoid
C0003873|Atrophic arthritis
C0003873|Systemic rheumatoid arthritis
C0003873|Chronic rheumatic arthritis
C0003873|Rheumatic gout
C0003873|RA - Rheumatoid arthritis
C0003873|RhA - Rheumatoid arthritis
C0003873|Rheumatoid disease
C0003873|atrophic; arthritis
C0003873|rheumatoid; arthritis
C0003873|arthritis; atrophic
C0003873|arthritis; rheumatoid
C0003873|Arthritis or polyarthritis, atrophic
C0003873|Arthritis or polyarthritis, rheumatic
C3495559|Chronic Arthritis, Juvenile
C3495559|Rheumatoid Arthritis, Juvenile
C3495559|Juvenile arthritis
C3495559|Juvenile arthritis, unspecified
C3495559|Arthritis, Juvenile Chronic
C3495559|Juvenile Idiopathic Arthritis
C3495559|Juvenile Chronic Arthritis
C3495559|Juvenile Rheumatoid Arthritis
C3495559|Arthritis, Juvenile Idiopathic
C3495559|juvenile arthritis (diagnosis)
C3495559|Arthritis, Juvenile
C3495559|Enthesitis Related Arthritis, Juvenile
C3495559|Juvenile Oligoarthritis
C3495559|Arthritis, Juvenile Systemic
C3495559|Juvenile Enthesitis-Related Arthritis
C3495559|Juvenile Systemic Arthritis
C3495559|Arthritis, Juvenile Psoriatic
C3495559|Juvenile Psoriatic Arthritis
C3495559|Arthritis, Juvenile Enthesitis-Related
C3495559|Oligoarthritis, Juvenile
C3495559|Arthritis, Juvenile Rheumatoid
C3495559|Enthesitis-Related Arthritis, Juvenile
C3495559|Psoriatic Arthritis, Juvenile
C3495559|Systemic Arthritis, Juvenile
C3495559|Arthritis, Juvenile [Disease/Finding]
C3495559|JIA
C3495559|Polyarthritis, Juvenile, Rheumatoid Factor Positive
C3495559|Polyarthritis, Juvenile, Rheumatoid Factor Negative
C3495559|JCA - Juvenile chronic arthritis
C3495559|Juvenile chronic arthritis (disorder)
C3495559|juvenile; arthritis
C3495559|arthritis; juvenile
C3495559|Juvenile chronic arthritis, polyarticular seropositive
C3495559|Juvenile idiopathic arthritis (disorder)
C3495559|Juvenile idiopathic arthritis, polyarthritis, rheumatoid factor positive
C3495559|Idiopathic Arthritis, Juvenile
C3495559|Arthritis;juvenile
C0409679|Seronegative arthritis
C0409679|Seronegative arthritis (disorder)
C0409679|Seronegative polyarthritis
C0409679|Sero negative arthropathy
C0409679|Seronegative arthritis NOS
C0409679|Seronegative arthropathy
C0409679|Seronegative arthritis [Ambiguous]
C0240903|Rheumatoid vasculitis
C0240903|rheumatoid vasculitis (diagnosis)
C0240903|Vasculitides, Rheumatoid
C0240903|Vasculitis, Rheumatoid
C0240903|Rheumatoid Vasculitides
C0240903|Rheumatoid Vasculitis [Disease/Finding]
C0240903|Rheumatoid vasculitis (disorder)
C0240903|rheumatoid; arthritis, with vasculitis
C0240903|rheumatoid; vasculitis
C0240903|vasculitis; rheumatoid
C0240903|arthritis; rheumatoid, with vasculitis
C2200410|rheumatoid arthritis of fingers
C2200410|rheumatoid arthritis of fingers (diagnosis)
C2200418|rheumatoid arthritis of toes (diagnosis)
C2200418|rheumatoid arthritis of toes
C0427391|Rheumatoid factor negative
C0427391|Negative rheumatoid factor
C0427391|rheumatoid factor negative (diagnosis)
C0427391|Rheumatiod factor negative
C0427391|Rheumatoid factor negative (finding)
C2200417|rheumatoid arthritis Steinbrocker classification (___0-IV)
C2200417|rheumatoid arthritis Steinbrocker classification (___0-IV) (diagnosis)
C2062580|rheumatoid arthritis with atlantoaxial subluxation (diagnosis)
C2062580|rheumatoid arthritis with atlantoaxial subluxation
C2931281|Sjogren-Mikulicz syndrome
C0085574|Palindromic rheumatism
C0085574|Palindrom rheum-unspec
C0085574|Palindromic rheumatism, unspecified site
C0085574|Palindromic rheumatism syndrome
C0085574|Palindromic rheumatism NOS (disorder)
C0085574|Palindromic rheumatism NOS
C0085574|Palindromic rheumatism of unspecified site (disorder)
C0085574|Hench - Rosenberg syndrome
C0085574|Palindromic rheumatism of unspecified site
C0085574|Palindromic rheumatism, site unspecified
C0085574|Hench-Rosenberg syndrome
C0085574|Palindromic rheumatism (disorder)
C0085574|palindromic; rheumatism
C0085574|rheumatism; palindromic
C3469328|rheumatoid arthritis nodule
C3469328|rheumatoid arthritis nodule (diagnosis)
C0451843|Rheumatoid bursitis
C0451843|Rheumatoid bursitis, unspecified site
C0451843|rheumatoid bursitis (diagnosis)
C0451843|Rheumatoid bursitis (disorder)
C0451843|bursitis; rheumatoid
C0451843|rheumatoid; bursitis
C2889134|Rheumatoid lung disease with rheumatoid arthritis of shoulder
C2889134|rheumatoid lung disease with rheumatoid arthritis of shoulder (diagnosis)
C2889138|Rheumatoid lung disease with rheumatoid arthritis of elbow
C2889138|rheumatoid lung disease with rheumatoid arthritis of elbow (diagnosis)
C2889143|Rheumatoid lung disease with rheumatoid arthritis of wrist
C2889143|rheumatoid lung disease with rheumatoid arthritis of wrist (diagnosis)
C2889148|Rheumatoid lung disease with rheumatoid arthritis of hand
C2889148|rheumatoid lung disease with rheumatoid arthritis of hand (diagnosis)
C2889152|Rheumatoid lung disease with rheumatoid arthritis of unspecified hip
C2889152|Rheumatoid lung disease with rheumatoid arthritis of hip
C2889152|Rheumatoid lung disease w rheumatoid arthritis of unsp hip
C2889152|rheumatoid lung disease with rheumatoid arthritis of hip (diagnosis)
C2889155|Rheumatoid lung disease with rheumatoid arthritis of knee
C2889155|rheumatoid lung disease with rheumatoid arthritis of knee (diagnosis)
C2889160|Rheumatoid lung disease with rheumatoid arthritis of ankle and foot
C2889160|rheumatoid lung disease with rheumatoid arthritis of ankle and foot (diagnosis)
C2889168|Rheumatoid vasculitis with rheumatoid arthritis of shoulder
C2889168|Rheumatoid vasculitis with rheumatoid arthritis of unspecified shoulder
C2889168|Rheu vasculitis w rheumatoid arthritis of unsp shoulder
C2889168|rheumatoid vasculitis with rheumatoid arthritis of shoulder (diagnosis)
C2889169|Rheumatoid vasculitis with rheumatoid arthritis of elbow
C2889169|rheumatoid vasculitis with rheumatoid arthritis of elbow (diagnosis)
C2889174|Rheumatoid vasculitis with rheumatoid arthritis of wrist
C2889174|rheumatoid vasculitis with rheumatoid arthritis of wrist (diagnosis)
C0564785|Rheumatoid arthritis of hand joint
C0564785|Rheumatoid arthritis - hand joint (disorder)
C0564785|Rheumatoid arthritis of hand joint (disorder)
C0564785|rheumatoid arthritis of hand (diagnosis)
C0564785|rheumatoid arthritis of hand
C0564785|Rheumatoid arthritis - hand joint
C0564786|Rheumatoid arthritis of ankle and/or foot
C0564786|Rheumatoid arthritis - ankle and/or foot (disorder)
C0564786|Rheumatoid arthritis of ankle and/or foot (disorder)
C0564786|rheumatoid arthritis of ankle and foot (diagnosis)
C0564786|rheumatoid arthritis of ankle and foot
C0564786|rheumatoid arthritis ankle and foot
C0564786|Rheumatoid arthritis - ankle/foot (disorder)
C0564786|Rheumatoid arthritis - ankle/foot
C0564786|Rheumatoid arthritis - ankle and/or foot
C3508970|rheumatoid arthritis vertebrae
C3508970|rheumatoid arthritis vertebrae (diagnosis)
C3508971|rheumatoid arthritis multiple sites
C3508971|rheumatoid arthritis multiple sites (diagnosis)
C0265176|Pericarditis secondary to rheumatoid arthritis
C0265176|Pericarditis secondary to rheumatoid arthritis (disorder)
C0265176|pericarditis; rheumatoid arthritis (etiology)
C0265176|pericarditis; rheumatoid arthritis (manifestation)
C0265176|rheumatoid arthritis; pericarditis (etiology)
C0265176|rheumatoid arthritis; pericarditis (manifestation)
C0265176|rheumatoid; arthritis, with pericarditis (etiology)
C0265176|rheumatoid; arthritis, with pericarditis (manifestation)
C0265176|arthritis; rheumatoid, with pericarditis (etiology)
C0265176|arthritis; rheumatoid, with pericarditis (manifestation)
C0564787|Rheumatoid arthritis - other joint
C0564787|Rheumatoid arthritis - other joint (disorder)
C0409649|Other rheumatoid arthritis of spine
C0409649|Other rheumatoid arthritis of spine (disorder)
C3836171|rheumatoid arthritis rf positive without involvement of other organs and systems
C3836171|rheumatoid arthritis rf positive without involvement of other organs and systems (diagnosis)
C3899278|Early Rheumatoid Arthritis
C0702102|Arthritis mutilans
C0702102|Psoriatic arthritis - destructive type
C0702102|Psoriatic arthritis - destructive type (disorder)
C0702102|Arthritis mutilans (disorder)
C0702102|mutilans; arthritis (etiology)
C0702102|mutilans; arthritis (manifestation)
C0702102|arthritis; mutilans (etiology)
C0702102|arthritis; mutilans (manifestation)
C0409653|Rheumatoid arthritis with organ / system involvement
C0409653|Rheumatoid arthritis with organ / system involvement (disorder)
C0477542|Other specified rheumatoid arthritis
C0477542|Other specified rheumatoid arthritis, unspecified site
C0477542|[X]Other specified rheumatoid arthritis
C0477542|[X]Other specified rheumatoid arthritis (disorder)
C0581345|Flare of rheumatoid arthritis
C0581345|Flare of rheumatoid arthritis (disorder)
C0564784|Rheumatoid arthritis of multiple joints
C0564784|Rheumatoid arthritis of multiple joints (disorder)
C0564784|Rheumatoid arthritis - multiple joint (disorder)
C0564784|Rheumatoid arthritis - multiple joint
C0263741|Extra-articular rheumatoid process (disorder)
C0263741|Extra-articular rheumatoid process
C0263741|Extra-articular rheumatoid process, NOS
C0866632|Arthritis or polyarthitis, chronic rheumatic
C1405320|polyarthritis; rheumatoid
C1405320|rheumatoid; polyarthritis
C1406307|rheumatoid\\see also condition
C0087031|Still's disease
C0087031|Juvenile Onset Still Disease
C0087031|Juvenile Onset Stills Disease
C0087031|Juvenile-Onset Still's Disease
C0087031|Still Disease, Juvenile Onset
C0087031|Still's Disease, Juvenile Onset
C0087031|Stills Disease, Juvenile-Onset
C0087031|Juvenile-Onset Still Disease
C0087031|STILL DISEASE JUVENILE ONSET
C0087031|JUVENILE ONSET STILL DIS
C0087031|JUVENILE ONSET STILLS DIS
C0087031|STILLS DIS JUVENILE ONSET
C0087031|Still's disease -RETIRED-
C0087031|juvenile onset Still's disease (diagnosis)
C0087031|juvenile Still's disease
C0087031|juvenile onset Still's disease
C0087031|Still Disease
C0087031|Still's disease NOS
C0087031|Still's disease - juvenile R.A
C0087031|Still's disease (disorder)
C0087031|Still's disease - juvenile rheumatoid arthritis (disorder)
C0087031|Still's disease - juvenile rheumatoid arthritis
C0087031|Systemic Onset Juvenile Rheumatoid Arthritis
C0087031|Systemic JRA
C0087031|sJRA
C0087031|Systemic Juvenile Rheumatoid Arthritis (AQ)
C0087031|Juvenile-Onset Stills Disease
C0087031|Still Disease, Juvenile-Onset
C0087031|Still's Disease, Juvenile-Onset
C0421288|Rheumatology disorder - joints affected (disorder)
C0421288|Rheumatology disorder - joints affected
C0421288|Rheumatology disorder - joints affected (finding)
C1998379|Rheumatoid arthritis of temporomandibular joint (disorder)
C1998379|Rheumatoid arthritis of temporomandibular joint
C1998063|Rheumatic arthritis of temporomandibular joint (disorder)
C1998063|Rheumatic arthritis of temporomandibular joint
C0585962|Seropositive errosive rheumatoid arthritis (disorder)
C0585962|Seropositive errosive rheumatoid arthritis
C1304220|Cutaneous complication of rheumatoid disease (disorder)
C1304220|Cutaneous complication of rheumatoid disease
C0409579|Articular rheumatic fever
C0409579|Rheumatic joint disease
C0409579|Arthritis due to rheumatic fever
C0409579|Rheumatic joint disease (disorder)
C0409579|Articular rheumatic fever, NOS
C0409579|Rheumatic joint disease, NOS
C1304215|Accelerated rheumatoid nodulosis (disorder)
C1304215|Accelerated rheumatoid nodulosis
C1997893|Rheumatoid arthritis of foot
C1997893|Rheumatoid arthritis of foot (disorder)
C0029408|Arthritides, Degenerative
C0029408|Degenerative Arthritides
C0029408|Osteoarthritides
C0029408|Osteoarthritis
C0029408|Osteoarthroses
C0029408|Degenerative Arthritis
C0029408|hypertrophic arthritis
C0029408|degenerative joint disease
C0029408|Osteoarthrosis
C0029408|OA
C0029408|DJD
C0029408|osteoarthrosis (diagnosis)
C0029408|osteoarthritis (diagnosis)
C0029408|Osteoarthritis NOS
C0029408|Osteoarthritis, unspecified site
C0029408|Arthritis, Degenerative
C0029408|Osteoarthritis [Disease/Finding]
C0029408|O/A
C0029408|Arthritis;degenerative
C0029408|Osteoarthritis;degenerative
C0029408|Osteoarthritis (M15-M19)
C0029408|Degenerative polyarthritis
C0029408|Degenerative joint disease (disorder)
C0029408|Degenerative arthropathy
C0029408|Joint degeneration
C0029408|Degenerative arthropathy (disorder)
C0029408|Osteoarthritis (& [allied disorders])
C0029408|Osteoarthritis (disorder)
C0029408|Osteoarthritis NOS (disorder)
C0029408|Hypertrophic polyarthritis
C0029408|[Joint degeneration] or [osteoarthritis NOS] (disorder)
C0029408|Osteoarthritis NOS, of unspecified site (disorder)
C0029408|Osteoarthritis and allied disorders
C0029408|OA - Osteoarthritis
C0029408|Osteoarthritis NOS, of unspecified site
C0029408|[Joint degeneration] or [osteoarthritis NOS]
C0029408|OA - Osteoarthrosis
C0029408|Osteoarthrosis, unspecified whether generalized or localized
C0029408|Degenerative polyarthritis (disorder)
C0029408|hypertrophy; arthritis
C0029408|arthritis; hypertrophy
C0029408|Degenerative arthritis, NOS
C0029408|Degenerative arthropathy, NOS
C0029408|Degenerative joint disease, NOS
C0029408|Degenerative polyarthritis, NOS
C0029408|Hypertrophic arthritis, NOS
C0029408|Hypertrophic polyarthritis, NOS
C0029408|Osteoarthritis, NOS
C0029408|degenerative osteoarthritis
C0029408|joint(s) degeneration
C0029408|Degeneration;joint(s)
C1306838|Proliferative arthritis
C1306838|Proliferative arthritis (disorder)
C1306838|Proliferative arthritis, NOS
C0157913|Rheumatoid arthritis and other inflammatory polyarthropathies
C0157913|Rheumatoid arthritis and other inflammatory polyarthropathies (disorder)
C0157919|Other specified inflammatory polyarthropathies
C0157919|Other specified inflammatory polyarthropathy
C0157919|Inflamm polyarthrop NEC
C0157919|Other specified inflammatory polyarthropathy (disorder)
C0157919|Other specified inflammatory polyarthropathy NOS (disorder)
C0157919|Other specified inflammatory polyarthropathy NOS
C0162323|Polyarthritis
C0162323|Polyarthritides
C0162323|Inflammatory polyarthropathy
C0162323|Inflammatory polyarthropathies
C0162323|Polyarthritis, unspecified
C0162323|polyarthritis (diagnosis)
C0162323|Inflamm polyarthrop NOS
C0162323|Inflammatory polyarthropathies (M05-M14)
C0162323|Inflammatory polyarthropathy NOS
C0162323|Inflammatory polyarthropathy NOS (disorder)
C0162323|Polyarthritis (disorder)
C0162323|Polyarthritis NOS
C0162323|[X]Inflammatory polyarthropathies (disorder)
C0162323|Inflammatory polyarthropathy (disorder)
C0162323|Polyarthropathy NOS -inflammat
C0162323|[X]Inflammatory polyarthropathies
C0162323|Polyarticular arthritis
C0162323|Inflammatory arthritis of multiple joints
C0162323|Unspecified inflammatory polyarthropathy
C0162323|Inflammatory polyarthropathy, NOS
C0162323|Polyarthritis, NOS
C0162323|Inflammatory polyarthropathy or polyarthritis NOS
C0409667|Juvenile Chronic Polyarthritis
C0409667|Polyarticular onset juvenile chronic arthritis (disorder)
C0409667|Juvenile chronic polyarthritis (disorder)
C0409667|Polyarticular onset juvenile chronic arthritis
C0409667|Polyarticular juvenile arthritis
C0409667|Juvenile chronic polyarthritis, NOS
C0152084|Chronic postrheumatic arthropathy
C0152084|Chronic postrheumatic arthropathy [Jaccoud]
C0152084|chronic postrheumatic arthropathy (diagnosis)
C0152084|Chronic postrheumatic arthropathy -RETIRED-
C0152084|Chr postrheum arthritis
C0152084|Jaccoud syndrome
C0152084|Chronic postrheumatic arthropathy [Jaccoud], unspecified site
C0152084|Chronic postrheumatic arthropathy, unspecified site
C0152084|Chronic postrheumatic arthropathy (disorder)
C0152084|Non-deforming erosive arthropathy
C0152084|Chronic post rheumatic arthropathy
C0152084|Jaccoud's arthropathy
C0152084|Jaccoud's syndrome
C0152084|Jaccoud's disease
C0152084|Jaccoud's arthritis
C0152084|Chronic post - rheumatic arthropathy
C0152084|Jaccoud's syndrome (disorder)
C0152084|arthropathy; Jaccoud
C0152084|Jaccoud; arthropathy
C0152084|Jaccoud
C3469325|Felty's syndrome, shoulder
C3469325|rheumatoid arthritis felty's syndrome shoulder
C3469325|Felty's syndrome of shoulder (diagnosis)
C3469325|Felty's syndrome of shoulder
C3469320|Felty's syndrome, elbow
C3469320|Felty's syndrome, unspecified elbow
C3469320|Felty's syndrome of elbow
C3469320|Felty's syndrome of elbow (diagnosis)
C3469320|rheumatoid arthritis felty's syndrome elbow
C3469326|Felty's syndrome, wrist
C3469326|Felty's syndrome of wrist
C3469326|Felty's syndrome of wrist (diagnosis)
C3469326|rheumatoid arthritis felty's syndrome wrist
C0837511|Felty's syndrome, hand
C0837511|Felty's syndrome, unspecified hand
C0837511|rheumatoid arthritis felty's syndrome hand
C0837511|Felty's syndrome of hand (diagnosis)
C0837511|Felty's syndrome of hand
C3469322|Felty's syndrome, hip
C3469322|Felty's syndrome, unspecified hip
C3469322|Felty's syndrome of hip (diagnosis)
C3469322|rheumatoid arthritis felty's syndrome hip
C3469322|Felty's syndrome of hip
C3469323|Felty's syndrome, unspecified knee
C3469323|Felty's syndrome, knee
C3469323|Felty's syndrome of knee
C3469323|Felty's syndrome of knee (diagnosis)
C3469323|rheumatoid arthritis felty's syndrome knee
C0837514|Felty's syndrome, ankle and foot
C0837514|rheumatoid arthritis felty's syndrome ankle and foot
C0837514|Felty's syndrome of ankle and foot
C0837514|Felty's syndrome of ankle and foot (diagnosis)
C0837507|Felty's syndrome, multiple sites
C0837507|Felty's syndrome of multiple sites (diagnosis)
C0837507|rheumatoid arthritis felty's syndrome multiple sites
C0837507|Felty's syndrome of multiple sites
C2936659|Familial Feltys Syndrome
C2936659|Felty's Syndrome, Familial
C2936659|Syndrome, Familial Felty's
C2936659|Syndrome, Familial Felty
C2936659|Felty Syndrome, Familial
C2936659|Familial Felty's Syndrome
C2936659|Rheumatoid Arthritis, Splenomegaly and Neutropenia
C2936659|Familial Felty Syndrome
C0234948|Polyarthritis generalized
C0234948|Polyarthritis generalised
C0520533|Polyarthritis acute
C0520533|Acute polyarthritis
C0520533|Acute polyarthritis (disorder)
C0158017|Unspecified polyarthropathy or polyarthritis involving shoulder region
C0158017|Polyarthritis NOS-shlder
C0158017|Unspecified polyarthropathy or polyarthritis, shoulder region
C0158018|Unspecified polyarthropathy or polyarthritis involving upper arm
C0158018|Polyarthritis NOS-up/arm
C0158018|Unspecified polyarthropathy or polyarthritis, upper arm
C0158019|Unspecified polyarthropathy or polyarthritis involving forearm
C0158019|Polyarthrit NOS-forearm
C0158019|Unspecified polyarthropathy or polyarthritis, forearm
C0158020|Unspecified polyarthropathy or polyarthritis involving hand
C0158020|Polyarthritis NOS-hand
C0158020|Unspecified polyarthropathy or polyarthritis, hand
C0158021|Unspecified polyarthropathy or polyarthritis involving pelvic region and thigh
C0158021|Polyarthritis NOS-pelvis
C0158021|Unspecified polyarthropathy or polyarthritis, pelvic region and thigh
C0158022|Unspecified polyarthropathy or polyarthritis involving lower leg
C0158022|Polyarthritis NOS-l/leg
C0158022|Unspecified polyarthropathy or polyarthritis, lower leg
C0158023|Unspecified polyarthropathy or polyarthritis involving ankle and foot
C0158023|Polyarthritis NOS-ankle
C0158023|Unspecified polyarthropathy or polyarthritis, ankle and foot
C0158024|Unspecified polyarthropathy or polyarthritis involving other specified sites
C0158024|Polyarthrit NOS-oth site
C0158024|Unspecified polyarthropathy or polyarthritis, other specified sites
C0856585|Polyarthropathy (excl rheumatoid arthritis)
C0856585|Polyarthropathy (excluding rheumatoid arthritis)
C0018099|Gout
C0018099|Gout, unspecified
C0018099|gout (diagnosis)
C0018099|Gout NOS
C0018099|Gout [Disease/Finding]
C0018099|Gouts
C0018099|Gout NOS (disorder)
C0018099|Gout (disorder)
C0018099|gout; in
C0018099|Gout, NOS
C0494904|Other arthritis
C0409848|Other crystal arthropathies
C0409848|Other crystal arthropathy NOS (disorder)
C0409848|Other crystal arthropathies (disorder)
C0409848|Other crystal arthropathies of unspecified site (disorder)
C0409848|Other crystal arthropathy NOS
C0409848|Other crystal arthropathies of unspecified site
C0494897|Other rheumatoid arthritis
C0029746|Other specified arthropathy
C0029746|Other specified disorders of joint
C0029746|Other specified arthropathy, site unspecified
C0029746|Other specified disorders of joint, site unspecified
C0029746|Other specified joint disorders
C0029746|Other specific arthropathies
C0029746|Arthropathy, other specified
C0029746|[X]Other specified joint disorders
C0029746|[X]Other specified joint disorders (disorder)
C0029746|Other specified arthropathies
C0029746|Other specified arthropathy of unspecified site (disorder)
C0029746|Other specified arthropathy NOS (disorder)
C0029746|Other specified arthropathy (disorder)
C0029746|Other specified arthropathy NOS
C0029746|Other specified arthropathy of unspecified site
C0029746|Other specified joint disorders of unspecified site (disorder)
C0029746|Other specified joint disorders of unspecified site
C0029746|Other specified joint disorders NOS (disorder)
C0029746|Other specified joint disorders (disorder)
C0029746|Other specified joint disorders NOS
C0029746|Other specified arthropathies (disorder)
C0694515|Psoriatic and enteropathic arthropathies
C0694516|Juvenile arthritis in diseases classified elsewhere
C0694517|Arthropathies in other diseases classified elsewhere
C2889385|Rheumatoid arthritis with rheumatoid factor, unspecified
C2889385|Rheumatoid arthritis with rheumatoid factor
C2889493|Enteropathic arthropathies
C2889493|enteropathic arthropathy (diagnosis)
C2889493|enteropathic arthropathy
C1442831|Other and unspecified arthropathies
C1442831|Other and unspecified disorders of joint
C1442831|Other joint disorders
C1442831|Other disorder of joint, NOS
C1442831|Other disorder of joint -RETIRED-
C1442831|Other and unspecified arthropathy
C1442831|Other joint disorders (M20-M25)
C1442831|[X]Other joint disorders
C1442831|Other disorder of joint (disorder)
C1442831|Other and unspecified joint disorders
C1442831|Other disorder of joint
C1442831|Other and unspecified joint disorders (disorder)
C1442831|[X]Other joint disorders (disorder)
C1442831|Other and unspecified arthropathies (disorder)
C2919482|RS3PE - Remitting seronegative symmetric synovitis with pitting edema
C2919482|Remitting seronegative symmetrical synovitis with pitting edema (disorder)
C2919482|Relapsing seronegative symmetrical synovitis with pitting oedema
C2919482|RS3PE - Remitting seronegative symmetric synovitis with pitting oedema
C2919482|Remitting seronegative symmetrical synovitis with pitting edema
C2919482|Remitting seronegative symmetrical synovitis with pitting oedema
C2919482|Relapsing seronegative symmetrical synovitis with pitting edema
C2111765|polyarthritis of shoulder (diagnosis)
C2111765|polyarthritis of shoulder
C2111767|polyarthritis of upper arm (diagnosis)
C2111767|polyarthritis of upper arm
C2083206|polyarthritis of forearm
C2083206|polyarthritis of forearm (diagnosis)
C2239149|polyarthritis hand
C2239149|polyarthritis of hand
C2239149|polyarthritis of hand (diagnosis)
C2083209|polyarthritis of pelvic region
C2083209|polyarthritis of pelvic region (diagnosis)
C2111766|polyarthritis of thigh (diagnosis)
C2111766|polyarthritis of thigh
C2083207|polyarthritis of lower leg (diagnosis)
C2083207|polyarthritis of lower leg
C2083204|polyarthritis ankle
C2083204|polyarthritis of ankle
C2083204|polyarthritis of ankle (diagnosis)
C2083205|polyarthritis of foot
C2083205|polyarthritis of foot (diagnosis)
C2083208|polyarthritis of multiple sites (diagnosis)
C2083208|polyarthritis of multiple sites
C0268108|Chronic gout
C0268108|gouty arthropathy chronic (diagnosis)
C0268108|gouty arthropathy chronic
C0268108|chronic gout (diagnosis)
C0268108|gout chronic
C0268108|Chronic gouty arthritis
C0268108|Chronic gouty arthritis (disorder)
C2103075|axial polyarticular inflammation (diagnosis)
C2103075|axial polyarticular inflammation
C3495373|arthritis of multiple sites
C3495373|arthritis multiple sites
C3495373|arthritis multiple sites (diagnosis)
C1260913|Pneumococcal arthritis and polyarthritis
C1260913|Pneumococcal arthritis and polyarthritis (disorder)
C1260913|Arthritis or Polyarthritis due to Pneumococcus
C1260913|Pneumococcal arthritis or polyarthritis
C0263721|Polyarthritis associated with disorder classified elsewhere
C0263721|Polyarthritis associated with another disorder (disorder)
C0263721|Polyarthritis associated with another disorder
C0275601|Nonsuppurative polyarthritis in lambs
C0275601|Nonsuppurative polyarthritis in lambs (disorder)
C0263735|Polyarthritis in Greyhounds
C0263735|Polyarthritis in Greyhounds (disorder)
C1290689|Arthritis of temporomandibular joint as part of polyarthritis (disorder)
C1290689|Arthritis of temporomandibular joint as part of polyarthritis
C1290689|Systemic arthritis including temporomandibular joint
C0263734|Progressive feline polyarthritis
C0263734|Progressive feline polyarthritis (disorder)
C0276035|Infectious polyarthritis
C0276035|Porcine polyserositis
C0276035|Glasser's disease (disorder)
C0276035|Glasser's disease
C0409668|Early onset polyarticular juvenile chronic arthritis
C0409668|Early onset polyarticular juvenile chronic arthritis (disorder)
C0263739|Polyarticular JCA
C0263739|Polyarticular juvenile chronic RA
C0263739|Chronic polyarticular juvenile rheumatoid arthritis
C0263739|Chronic polyarticular juvenile rheumatoid arthritis (disorder)
C0409510|Infective arthritis of multiple sites
C0409510|Infective polyarthritis
C0409510|Infective arthritis NOS, of multiple sites
C0409510|Infective arthritis NOS, of multiple sites (disorder)
C0409510|Infective polyarthritis (disorder)
C0409510|Infective polyarthritis, NOS
C0477535|Arthritis and polyarthritis due to other specified bacterial agents
C0477535|[X]Arthritis and polyarthritis due to other specified bacterial agents
C0477535|[X]Arthritis and polyarthritis due to other specified bacterial agents (disorder)
C0276114|Chlamydial polyarthritis
C0276114|Transmissible serositis
C0276114|Chlamydial polyarthritis (disorder)
C0240344|Migratory polyarthritis (disorder)
C0240344|Migratory polyarthritis
C0240344|Migratory polyarthritis, NOS
C0409669|Late onset polyarticular juvenile chronic arthritis
C0409669|Late onset polyarticular juvenile chronic arthritis (disorder)
C0409702|Undifferentiated inflammatory oligoarthritis
C0409702|Undifferentiated inflammatory oligoarthritis (disorder)
C0263736|Enzootic polyarthritis in goats (disorder)
C0263736|Enzootic polyarthritis in goats
C0263733|Idiopathic polyarthritis
C0263733|Idiopathic polyarthritis (disorder)
C0311284|Lipoid dermatoarthritis
C0311284|lipoid metabolism disorder lipoid dermatoarthritis
C0311284|lipoid dermatoarthritis (diagnosis)
C0311284|Multicentric reticulohistiocytosis
C0311284|Multicentric reticulohistiocytosis (disorder)
C0311284|Nicolau-Balus syndrome
C0311284|Lipoid dermatoarthritis (disorder)
C1302753|Fibroblastic rheumatism (disorder)
C1302753|Fibroblastic rheumatism
C1535016|Polyarthropathy (& [inflammatory]) NOS (disorder)
C1535016|Polyarthropathy (& [inflammatory]) NOS
C3646092|spondylopathy inflammatory multiple sites spine
C3646092|spondylopathy inflammatory multiple sites spine (diagnosis)
C3687214|Immune mediated polyarthritis
C3687214|Immune mediated polyarthritis (disorder)
C0477553|Arthropathies in other endocrine, nutritional and metabolic disorders
C0477553|[X]Arthropathies in other endocrine, nutritional and metabolic disorders
C0477553|[X]Arthropathies in other endocrine, nutritional and metabolic disorders (disorder)
C0477554|Arthropathies in other specified diseases classified elsewhere
C0477554|[X]Arthropathies in other specified diseases classified elsewhere
C0477554|[X]Arthropathies in other specified diseases classified elsewhere (disorder)
C0477549|Other specific arthropathies, NEC in SNOMEDCT
C0477549|[X]Other specific arthropathies, not elsewhere classified
C0477549|[X]Other specific arthropathies, not elsewhere classified (disorder)
C0477550|Other specified arthritis
C0477550|Other specified arthritis, unspecified site
C0477550|[X]Other specified arthritis (disorder)
C0477550|[X]Other specified arthritis
C0003892|Neurogenic arthropathy
C0003892|Arthropathies, Neurogenic
C0003892|Arthropathy, Neurogenic
C0003892|Charcot Joint
C0003892|Charcots Joint
C0003892|Neurogenic Arthropathies
C0003892|Arthropathy associated with neurological disorders
C0003892|Joint, Charcot's
C0003892|Neuropathic arthropathy
C0003892|neuropathic joint disease (diagnosis)
C0003892|Charcot's arthropathy
C0003892|Charcot's arthropathy (diagnosis)
C0003892|neuropathic joint disease
C0003892|Charcot's joint was observed
C0003892|Charcot's joint (physical finding)
C0003892|Charcot's joint
C0003892|Arthropathy w nerve dis
C0003892|Charcot arthropathy
C0003892|Arthropathy, Neurogenic [Disease/Finding]
C0003892|Neuropathic arthropathy (& Charcot's) (disorder)
C0003892|Charcot's arthropathy (disorder)
C0003892|Neuropathic arthropathy (& Charcot's)
C0003892|Neurogenic arthropathy of Charcot
C0003892|Neurogenic arthropathy of Charcot (disorder)
C0003892|Charcot joints
C0003892|Arthropathy neurogenic
C0003892|Arthropathy associated with a neurological disorder
C0003892|Arthropathy associated with a neurological disorder (disorder)
C0003892|Charcot's joint disease
C0003892|Charcot's arthropathy (disorder) [Ambiguous]
C0003892|Neurogenic arthropathy of Charcot (disorder) [Ambiguous]
C1692871|Inflammatory polyarthritis
C1692871|inflammatory; polyarthritis
C1692871|polyarthritis; inflammatory
C1692871|Inflammatory polyarthritis, NOS
C1692872|Undifferentiated inflammatory polyarthritis
C1692872|Undifferentiated inflammatory polyarthritis (disorder)
C0409252|Allergic arthritis involving multiple sites
C0409252|allergic arthritis of multiple sites (diagnosis)
C0409252|allergic arthritis of multiple sites
C0409252|Allerg arthritis-mult
C0409252|Allergic arthritis, multiple sites
C0409252|Allergic arthritis of multiple sites (disorder)
C0157916|Acute polyarticular juvenile rheumatoid arthritis
C0157916|Polyart juv rheum arthr
C0157916|Acute polyarticular juvenile rheumatoid arthritis (disorder)
C0157916|Polyarticular juvenile rheumatoid arthritis, acute
C0157916|acute polyarticular juvenile idiopathic arthritis (diagnosis)
C0157916|juvenile idiopathic arthritis, polyarticular acute
C0157916|acute polyarticular juvenile idiopathic arthritis
C0157916|Acute juvenile rheumatoid arthritis
C0157916|Acute polyarticular juvenile rheumatoid arthritis [dup] (disorder)
C1827497|Post-infective polyarthritis
C1827497|Reactive arthritis of multiple sites
C1827497|Post-infective polyarthritis (disorder)
C0409703|Secondary inflammatory arthritis
C0409703|Secondary inflammatory arthritis (disorder)
C2889165|Rheumatoid vasculitis with rheumatoid arthritis
C2889165|Rheumatoid vasculitis with rheumatoid arthritis of unspecified site
C2889165|Rheumatoid vasculitis with rheumatoid arthritis of unsp site
C2889165|rheumatoid vasculitis with rheumatoid arthritis (diagnosis)
C2889179|Rheumatoid vasculitis with rheumatoid arthritis of unspecified hand
C2889179|Rheumatoid vasculitis with rheumatoid arthritis of hand
C2889179|Rheumatoid vasculitis with rheumatoid arthritis of unsp hand
C2889179|rheumatoid vasculitis with rheumatoid arthritis of hand (diagnosis)
C2889182|Rheumatoid vasculitis with rheumatoid arthritis of hip
C2889182|rheumatoid vasculitis with rheumatoid arthritis of hip (diagnosis)
C2889186|Rheumatoid vasculitis with rheumatoid arthritis of knee
C2889186|rheumatoid vasculitis with rheumatoid arthritis of knee (diagnosis)
C2889195|Rheumatoid vasculitis with rheumatoid arthritis of multiple sites
C2889195|Rheumatoid vasculitis w rheumatoid arthritis mult site
C2889195|rheumatoid vasculitis with rheumatoid arthritis of multiple sites (diagnosis)
C0264993|Rheumatoid arteritis
C0264993|Rheumatoid arteritis (disorder)
C0343204|Necrotizing rheumatoid vasculitis
C0343204|necrotizing rheumatoid vasculitis (diagnosis)
C0343204|Necrotising rheumatoid vasculitis
C0343204|Necrotizing rheumatoid vasculitis (disorder)
C0343202|Nailfold rheumatoid vasculitis
C0343202|Nailfold rheumatoid vasculitis (disorder)
C0343203|Systemic rheumatoid vasculitis
C0343203|Systemic rheumatoid vasculitis (disorder)
C1276120|Bywater lesions
C1276120|Nailfold/finger-pulp infarcts in rheumatoid disease (disorder)
C1276120|Nailfold/finger-pulp infarcts in rheumatoid disease
C0155555|Acute rheumatic pericarditis
C0155555|acute rheumatic pericarditis (diagnosis)
C0155555|Acute rheumatic pericard
C0155555|Rheumatic pericarditis (acute)
C0155555|Pericarditis;rheumatic;acute
C0155555|Acute rheumatic pericarditis (disorder)
C0155555|Active rheumatic fever with pericarditis
C0155555|Acute rheumatic fever with pericarditis
C0155555|acute; pericarditis, rheumatic
C0155555|pericarditis; acute, rheumatic
C0155555|pericarditis; with rheumatic fever, active
C0155555|rheumatic fever; in pericarditis, active
C0155555|Rheumatic pericarditis, acute
C0155561|Chronic rheumatic pericarditis
C0155561|chronic rheumatic pericarditis (diagnosis)
C0155561|Chr rheumatic pericard
C0155561|Pericarditis;rheumatic;chronic
C0155561|Chronic rheumatic pericarditis NOS
C0155561|Chronic rheumatic pericarditis (disorder)
C0155561|Chronic rheumatic pericarditis NOS (disorder)
C0264747|rheumatic pericarditis (diagnosis)
C0264747|rheumatic pericarditis
C0264747|Pericarditis rheumatic
C0264747|Rheumatoid pericarditis
C0264747|Rheumatic pericarditis (disorder)
C0264747|pericarditis; rheumatic fever
C0264747|pericarditis; rheumatic
C0264747|rheumatic fever; pericarditis
C0264747|rheumatic; pericarditis
C0264747|Rheumatic pericarditis, NOS
C0264747|Rheumatic fever with pericarditis
C0392469|Rheumatoid carditis
C0392469|Rheumatoid carditis (disorder)
C0994344|Rheumatoid lung
C0994344|Rheumatoid lung disease
C0994344|Rheumatoid lung (disorder)
C0994344|Rheumatoid lung disease (disorder)
C0994344|lung; rheumatoid (etiology)
C0994344|lung; rheumatoid (manifestation)
C0994344|rheumatoid; arthritis, with lung involvement (etiology)
C0994344|rheumatoid; arthritis, with lung involvement (manifestation)
C0994344|rheumatoid; lung (etiology)
C0994344|rheumatoid; lung (manifestation)
C0994344|arthritis; rheumatoid, with lung involvement (etiology)
C0994344|arthritis; rheumatoid, with lung involvement (manifestation)
C0151379|Rheumatoid factor positive
C0151379|Rheumatoid factor positive (finding)
C3508972|rheumatoid arthritis rf positive of shoulder
C3508972|rheumatoid arthritis rf positive of shoulder (diagnosis)
C3508973|rheumatoid arthritis rf positive of elbow
C3508973|rheumatoid arthritis rf positive of elbow (diagnosis)
C3508974|rheumatoid arthritis rf positive of wrist
C3508974|rheumatoid arthritis rf positive of wrist (diagnosis)
C3508975|rheumatoid arthritis rf positive of hand
C3508975|rheumatoid arthritis rf positive of hand (diagnosis)
C3508976|rheumatoid arthritis rf positive of hip (diagnosis)
C3508976|rheumatoid arthritis rf positive of hip
C3508977|rheumatoid arthritis rf positive of knee (diagnosis)
C3508977|rheumatoid arthritis rf positive of knee
C3508978|rheumatoid arthritis rf positive of ankle and foot
C3508978|rheumatoid arthritis rf positive of ankle and foot (diagnosis)
C3508979|rheumatoid arthritis rf positive of multiple sites
C3508979|rheumatoid arthritis rf positive of multiple sites (diagnosis)
C3507373|rheumatoid arthritis rf positive with involvement of other organs and systems (diagnosis)
C3507373|rheumatoid arthritis rf positive with involvement of other organs and systems
C0848642|Sacroilitis
C0489959|Rheumatic myocarditis
C0489959|Rheumatoid myocarditis
C0489959|Myocarditis rheumatic
C0489959|Rheumatic degeneration of myocardium
C0489959|Rheumatic myocarditis (disorder)
C0489959|Rheumatoid myocarditis (disorder)
C0489959|myocarditis; rheumatic
C0489959|rheumatic; myocarditis
C1563314|Rheumatic myocarditis (& [chronic])
C1563314|Rheumatic myocarditis (& [chronic]) (disorder)
C0155557|Acute rheumatic myocarditis
C0155557|acute rheumatic myocarditis (diagnosis)
C0155557|Ac rheumatic myocarditis
C0155557|Myocarditis;rheumatic;acute
C0155557|Acute rheumatic myocarditis (disorder)
C0155557|Active rheumatic fever with myocarditis
C0155557|Acute rheumatic fever with myocarditis
C0155557|acute; myocarditis, rheumatic
C0155557|myocarditis; rheumatic fever, active or acute
C0155557|myocarditis; rheumatic fever
C0155557|myocarditis; rheumatic, active or acute
C0155557|rheumatic fever; myocarditis, active or acute
C0155557|rheumatic; myocarditis, active or acute
C0155557|Acute rheumatic myocarditis (disorder) [Ambiguous]
C0155557|Rheumatic fever with myocarditis
C0264752|chronic rheumatic myocarditis
C0264752|chronic rheumatic myocarditis (diagnosis)
C0264752|Myocarditis;rheumatic;chronic
C0264752|Myocarditis-RH chronic
C0264752|Chronic rheumatic heart disease with myocarditis
C0264752|Chronic rheumatic heart disease with myocarditis (disorder)
C0264756|chronic rheumatic myopericarditis
C0264756|chronic rheumatic myopericarditis (diagnosis)
C0264756|Chronic rheumatic myopericarditis (disorder)
C0264756|chronic; rheumatic myopericarditis
C0264756|myopericarditis; chronic rheumatic
C0264756|Chronic rheumatic, myopericarditis
C1386193|rheumatic fever; inactive or quiescent with myocarditis, myocardial degeneration, myocardial degeneration
C1386196|rheumatic fever; myocarditis, inactive or chronic
C0003960|Bodies, Aschoff
C0003960|Aschoff body
C0003960|Aschoff nodule
C0003960|Aschoff body (morphologic abnormality)
C0003960|Aschoff's bodies
C0003960|bodies; Aschoff
C0003960|Aschoff; bodies
C0003960|Aschoff Bodies
C1391999|cardiomyopathy; rheumatic
C1391999|rheumatic; cardiomyopathy
C1395016|degeneration; myocardial, with rheumatic fever
C1395019|degeneration; myocardial, with rheumatic fever, inactive
C1404473|insufficiency; myocardial, with rheumatic fever
C1404473|myocardium; insufficiency, with rheumatic fever
C1404476|insufficiency; myocardial, with rheumatic fever, inactive or quiescent (with chorea)
C1404476|myocardium; insufficiency, with rheumatic fever, inactive or quiescent (with chorea)
C1404477|insufficiency; myocardial, rheumatic
C1404477|myocardium; insufficiency, rheumatic
C1404480|insufficiency; myocardial, rheumatic, inactive or quiescent (with chorea)
C1404480|myocardium; insufficiency, rheumatic, inactive or quiescent (with chorea)
C0837546|Rheumatoid arthritis of unspecified site with involvement of other organs and systems
C0837546|Rheu arthritis of unsp site w involv of organs and systems
C2889296|Rheumatoid arthritis of shoulder with involvement of other organs and systems
C2889300|Rheumatoid arthritis of elbow with involvement of other organs and systems
C2889305|Rheumatoid arthritis of wrist with involvement of other organs and systems
C0837541|Rheumatoid arthritis of hand with involvement of other organs and systems
C2889313|Rheumatoid arthritis of hip with involvement of other organs and systems
C2889317|Rheumatoid arthritis of knee with involvement of other organs and systems
C0837544|Rheumatoid arthritis of ankle and foot with involvement of other organs and systems
C0837537|Rheumatoid arthritis of multiple sites with involvement of other organs and systems
C0837537|Rheu arthritis mult site w involv of organs and systems
C1384964|disease (or disorder); heart, in rheumatoid arthritis (etiology)
C1384964|disease (or disorder); heart, in rheumatoid arthritis (manifestation)
C1388626|rheumatoid; arthritis, with involvement of organs
C1388626|arthritis; rheumatoid, with involvement of organs
C1388627|rheumatoid; arthritis, with carditis (etiology)
C1388627|rheumatoid; arthritis, with carditis (manifestation)
C1388627|arthritis; rheumatoid, with carditis (etiology)
C1388627|arthritis; rheumatoid, with carditis (manifestation)
C1388628|endocarditis; rheumatoid arthritis (etiology)
C1388628|endocarditis; rheumatoid arthritis (manifestation)
C1388628|rheumatoid arthritis; endocarditis (etiology)
C1388628|rheumatoid arthritis; endocarditis (manifestation)
C1388628|rheumatoid; arthritis, with endocarditis (etiology)
C1388628|rheumatoid; arthritis, with endocarditis (manifestation)
C1388628|arthritis; rheumatoid, with endocarditis (etiology)
C1388628|arthritis; rheumatoid, with endocarditis (manifestation)
C1388629|rheumatoid; arthritis, with heart involvement (etiology)
C1388629|rheumatoid; arthritis, with heart involvement (manifestation)
C1388629|arthritis; rheumatoid, with heart involvement (etiology)
C1388629|arthritis; rheumatoid, with heart involvement (manifestation)
C1388630|myocarditis; rheumatoid arthritis (etiology)
C1388630|myocarditis; rheumatoid arthritis (manifestation)
C1388630|rheumatoid arthritis; myocarditis (etiology)
C1388630|rheumatoid arthritis; myocarditis (manifestation)
C1388630|rheumatoid; arthritis, with myocarditis (etiology)
C1388630|rheumatoid; arthritis, with myocarditis (manifestation)
C1388630|arthritis; rheumatoid, with myocarditis (etiology)
C1388630|arthritis; rheumatoid, with myocarditis (manifestation)
C0343237|Myopathy due to rheumatoid arthritis
C0343237|Myopathy due to rheumatoid arthritis (disorder)
C0343237|myopathy; rheumatoid arthritis (etiology)
C0343237|myopathy; rheumatoid arthritis (manifestation)
C0343237|rheumatoid arthritis; myopathy (etiology)
C0343237|rheumatoid arthritis; myopathy (manifestation)
C0343237|rheumatoid; arthritis, with myopathy (etiology)
C0343237|rheumatoid; arthritis, with myopathy (manifestation)
C0343237|arthritis; rheumatoid, with myopathy (etiology)
C0343237|arthritis; rheumatoid, with myopathy (manifestation)
C0338555|Polyneuropathy in rheumatoid arthritis
C0338555|Polyneuropathy in rheumatoid arthritis (disorder)
C0338555|polyneuropathy; rheumatoid arthritis (etiology)
C0338555|polyneuropathy; rheumatoid arthritis (manifestation)
C0338555|rheumatoid arthritis; polyneuropathy (etiology)
C0338555|rheumatoid arthritis; polyneuropathy (manifestation)
C0338555|rheumatoid; arthritis, with polyneuropathy (etiology)
C0338555|rheumatoid; arthritis, with polyneuropathy (manifestation)
C0338555|arthritis; rheumatoid, with polyneuropathy (etiology)
C0338555|arthritis; rheumatoid, with polyneuropathy (manifestation)
C1388632|rheumatoid; arthritis, with visceral involvement
C1388632|arthritis; rheumatoid, with visceral involvement
C1392056|carditis; rheumatoid (etiology)
C1392056|carditis; rheumatoid (manifestation)
C1392056|rheumatoid; carditis (etiology)
C1392056|rheumatoid; carditis (manifestation)
C1399132|heart; disease, in rheumatoid arthritis (etiology)
C1399132|heart; disease, in rheumatoid arthritis (manifestation)
C1404498|myocarditis; rheumatoid (etiology)
C1404498|myocarditis; rheumatoid (manifestation)
C1404498|rheumatoid; myocarditis (etiology)
C1404498|rheumatoid; myocarditis (manifestation)
C1406303|pericarditis; rheumatoid (etiology)
C1406303|pericarditis; rheumatoid (manifestation)
C1406303|rheumatoid; pericarditis (etiology)
C1406303|rheumatoid; pericarditis (manifestation)
C2889120|Felty's syndrome, right hand
C2889121|Felty's syndrome, left hand
C2889129|Felty's syndrome, right ankle and foot
C2889130|Felty's syndrome, left ankle and foot
C2889131|Felty's syndrome, unspecified ankle and foot
C2889310|Rheumatoid arthritis of right hand with involvement of other organs and systems
C2889310|Rheu arthritis of right hand w involv of organs and systems
C2889311|Rheumatoid arthritis of left hand with involvement of other organs and systems
C2889311|Rheu arthritis of left hand w involv of organs and systems
C2889312|Rheumatoid arthritis of unspecified hand with involvement of other organs and systems
C2889312|Rheu arthritis of unsp hand w involv of organs and systems
C2889322|Rheumatoid arthritis of right ankle and foot with involvement of other organs and systems
C2889322|Rheu arthrit of right ank/ft w involv of organs and systems
C2889323|Rheumatoid arthritis of left ankle and foot with involvement of other organs and systems
C2889323|Rheu arthritis of left ank/ft w involv of organs and systems
C2889324|Rheumatoid arthritis of unspecified ankle and foot with involvement of other organs and systems
C2889324|Rheu arthritis of unsp ank/ft w involv of organs and systems
C2889132|Rheumatoid lung disease with rheumatoid arthritis
C2889132|rheumatoid lung disease with rheumatoid arthritis (diagnosis)
C1385071|disease (or disorder); lung, rheumatoid (diffuse) (interstitial) (etiology)
C1385071|disease (or disorder); lung, rheumatoid (diffuse) (interstitial) (manifestation)
C1385071|lung; disease, rheumatoid (diffuse) (interstitial) (etiology)
C1385071|lung; disease, rheumatoid (diffuse) (interstitial) (manifestation)
C1385163|disease (or disorder); respiratory, in rheumatoid arthritis (etiology)
C1385163|disease (or disorder); respiratory, in rheumatoid arthritis (manifestation)
C1405189|pneumoconiosis; rheumatoid (etiology)
C1405189|pneumoconiosis; rheumatoid (manifestation)
C1405189|rheumatoid; pneumoconiosis (etiology)
C1405189|rheumatoid; pneumoconiosis (manifestation)
C1406187|respiratory; disorder, in rheumatoid arthritis (etiology)
C1406187|respiratory; disorder, in rheumatoid arthritis (manifestation)
C3505955|rheumatoid necrobiotic nodule (diagnosis)
C3505955|rheumatoid necrobiotic nodule
C3505955|rheumatoid nodule
C3505955|rheumatoid arthritis - necrobiotic nodule
C2889108|Felty's syndrome, right shoulder
C2889109|Felty's syndrome, left shoulder
C2889110|Felty's syndrome, unspecified shoulder
C2889112|Felty's syndrome, right elbow
C2889113|Felty's syndrome, left elbow
C2889116|Felty's syndrome, right wrist
C2889117|Felty's syndrome, left wrist
C2889118|Felty's syndrome, unspecified wrist
C2889122|Felty's syndrome, right hip
C2889123|Felty's syndrome, left hip
C2889126|Felty's syndrome, right knee
C2889127|Felty's syndrome, left knee
C2889133|Rheumatoid lung disease with rheumatoid arthritis of unspecified site
C2889133|Rheumatoid lung disease w rheumatoid arthritis of unsp site
C2889164|Rheumatoid lung disease with rheumatoid arthritis of multiple sites
C2889164|Rheumatoid lung disease w rheumatoid arthritis mult site
C2889164|rheumatoid lung disease with rheumatoid arthritis of multiple sites (diagnosis)
C2889135|Rheumatoid lung disease with rheumatoid arthritis of right shoulder
C2889135|Rheumatoid lung disease w rheumatoid arthritis of r shoulder
C2889136|Rheumatoid lung disease with rheumatoid arthritis of left shoulder
C2889136|Rheumatoid lung disease w rheumatoid arthritis of l shoulder
C2889137|Rheumatoid lung disease with rheumatoid arthritis of unspecified shoulder
C2889137|Rheu lung disease w rheumatoid arthritis of unsp shoulder
C2889139|Rheumatoid lung disease with rheumatoid arthritis of right elbow
C2889139|Rheumatoid lung disease w rheumatoid arthritis of r elbow
C2889140|Rheumatoid lung disease with rheumatoid arthritis of left elbow
C2889140|Rheumatoid lung disease w rheumatoid arthritis of left elbow
C2889141|Rheumatoid lung disease with rheumatoid arthritis of unspecified elbow
C2889141|Rheumatoid lung disease w rheumatoid arthritis of unsp elbow
C2889144|Rheumatoid lung disease with rheumatoid arthritis of right wrist
C2889144|Rheumatoid lung disease w rheumatoid arthritis of r wrist
C2889145|Rheumatoid lung disease with rheumatoid arthritis of left wrist
C2889145|Rheumatoid lung disease w rheumatoid arthritis of left wrist
C2889146|Rheumatoid lung disease with rheumatoid arthritis of unspecified wrist
C2889146|Rheumatoid lung disease w rheumatoid arthritis of unsp wrist
C2889149|Rheumatoid lung disease with rheumatoid arthritis of right hand
C2889149|Rheumatoid lung disease w rheumatoid arthritis of right hand
C2889150|Rheumatoid lung disease with rheumatoid arthritis of left hand
C2889150|Rheumatoid lung disease w rheumatoid arthritis of left hand
C2889151|Rheumatoid lung disease with rheumatoid arthritis of unspecified hand
C2889151|Rheumatoid lung disease w rheumatoid arthritis of unsp hand
C2889153|Rheumatoid lung disease with rheumatoid arthritis of right hip
C2889153|Rheumatoid lung disease w rheumatoid arthritis of right hip
C2889154|Rheumatoid lung disease with rheumatoid arthritis of left hip
C2889154|Rheumatoid lung disease w rheumatoid arthritis of left hip
C2889156|Rheumatoid lung disease with rheumatoid arthritis of right knee
C2889156|Rheumatoid lung disease w rheumatoid arthritis of right knee
C2889157|Rheumatoid lung disease with rheumatoid arthritis of left knee
C2889157|Rheumatoid lung disease w rheumatoid arthritis of left knee
C2889158|Rheumatoid lung disease with rheumatoid arthritis of unspecified knee
C2889158|Rheumatoid lung disease w rheumatoid arthritis of unsp knee
C2889161|Rheumatoid lung disease with rheumatoid arthritis of right ankle and foot
C2889161|Rheu lung disease w rheumatoid arthritis of right ank/ft
C2889162|Rheumatoid lung disease with rheumatoid arthritis of left ankle and foot
C2889162|Rheu lung disease w rheumatoid arthritis of left ank/ft
C2889163|Rheumatoid lung disease with rheumatoid arthritis of unspecified ankle and foot
C2889163|Rheu lung disease w rheumatoid arthritis of unsp ank/ft
C2889191|Rheumatoid vasculitis with rheumatoid arthritis of ankle and foot
C2889191|rheumatoid vasculitis with rheumatoid arthritis of ankle and foot (diagnosis)
C2889166|Rheumatoid vasculitis with rheumatoid arthritis of right shoulder
C2889166|Rheumatoid vasculitis w rheumatoid arthritis of r shoulder
C2889167|Rheumatoid vasculitis with rheumatoid arthritis of left shoulder
C2889167|Rheumatoid vasculitis w rheumatoid arthritis of l shoulder
C2889170|Rheumatoid vasculitis with rheumatoid arthritis of right elbow
C2889170|Rheumatoid vasculitis w rheumatoid arthritis of right elbow
C2889171|Rheumatoid vasculitis with rheumatoid arthritis of left elbow
C2889171|Rheumatoid vasculitis w rheumatoid arthritis of left elbow
C2889172|Rheumatoid vasculitis with rheumatoid arthritis of unspecified elbow
C2889172|Rheumatoid vasculitis w rheumatoid arthritis of unsp elbow
C2889175|Rheumatoid vasculitis with rheumatoid arthritis of right wrist
C2889175|Rheumatoid vasculitis w rheumatoid arthritis of right wrist
C2889176|Rheumatoid vasculitis with rheumatoid arthritis of left wrist
C2889176|Rheumatoid vasculitis w rheumatoid arthritis of left wrist
C2889177|Rheumatoid vasculitis with rheumatoid arthritis of unspecified wrist
C2889177|Rheumatoid vasculitis w rheumatoid arthritis of unsp wrist
C2889180|Rheumatoid vasculitis with rheumatoid arthritis of right hand
C2889180|Rheumatoid vasculitis w rheumatoid arthritis of right hand
C2889181|Rheumatoid vasculitis with rheumatoid arthritis of left hand
C2889183|Rheumatoid vasculitis with rheumatoid arthritis of right hip
C2889184|Rheumatoid vasculitis with rheumatoid arthritis of left hip
C2889185|Rheumatoid vasculitis with rheumatoid arthritis of unspecified hip
C2889185|Rheumatoid vasculitis with rheumatoid arthritis of unsp hip
C2889187|Rheumatoid vasculitis with rheumatoid arthritis of right knee
C2889187|Rheumatoid vasculitis w rheumatoid arthritis of right knee
C2889188|Rheumatoid vasculitis with rheumatoid arthritis of left knee
C2889189|Rheumatoid vasculitis with rheumatoid arthritis of unspecified knee
C2889189|Rheumatoid vasculitis with rheumatoid arthritis of unsp knee
C2889192|Rheumatoid vasculitis with rheumatoid arthritis of right ankle and foot
C2889192|Rheumatoid vasculitis w rheumatoid arthritis of right ank/ft
C2889193|Rheumatoid vasculitis with rheumatoid arthritis of left ankle and foot
C2889193|Rheumatoid vasculitis w rheumatoid arthritis of left ank/ft
C2889194|Rheumatoid vasculitis with rheumatoid arthritis of unspecified ankle and foot
C2889194|Rheumatoid vasculitis w rheumatoid arthritis of unsp ank/ft
C2889198|Rheumatoid heart disease with rheumatoid arthritis of unspecified site
C2889198|Rheumatoid heart disease w rheumatoid arthritis of unsp site
C2889199|Rheumatoid heart disease with rheumatoid arthritis of shoulder
C2889199|rheumatoid heart disease with rheumatoid arthritis of shoulder (diagnosis)
C2889203|Rheumatoid heart disease with rheumatoid arthritis of elbow
C2889203|rheumatoid heart disease with rheumatoid arthritis of elbow (diagnosis)
C2889208|Rheumatoid heart disease with rheumatoid arthritis of wrist
C2889208|rheumatoid heart disease with rheumatoid arthritis of wrist (diagnosis)
C2889213|Rheumatoid heart disease with rheumatoid arthritis of hand
C2889213|rheumatoid heart disease with rheumatoid arthritis of hand (diagnosis)
C2889217|Rheumatoid heart disease with rheumatoid arthritis of hip
C2889217|Rheumatoid heart disease with rheumatoid arthritis of unspecified hip
C2889217|Rheumatoid heart disease w rheumatoid arthritis of unsp hip
C2889217|rheumatoid heart disease with rheumatoid arthritis of hip (diagnosis)
C2889220|Rheumatoid heart disease with rheumatoid arthritis of knee
C2889220|rheumatoid heart disease with rheumatoid arthritis of knee (diagnosis)
C2889225|Rheumatoid heart disease with rheumatoid arthritis of ankle and foot
C2889225|rheumatoid heart disease with rheumatoid arthritis of ankle and foot (diagnosis)
C2889229|Rheumatoid heart disease with rheumatoid arthritis of multiple sites
C2889229|Rheumatoid heart disease w rheumatoid arthritis mult site
C2889229|rheumatoid heart disease with rheumatoid arthritis of multiple sites (diagnosis)
C2889200|Rheumatoid heart disease with rheumatoid arthritis of right shoulder
C2889200|Rheu heart disease w rheumatoid arthritis of r shoulder
C2889201|Rheumatoid heart disease with rheumatoid arthritis of left shoulder
C2889201|Rheu heart disease w rheumatoid arthritis of l shoulder
C2889202|Rheumatoid heart disease with rheumatoid arthritis of unspecified shoulder
C2889202|Rheu heart disease w rheumatoid arthritis of unsp shoulder
C2889204|Rheumatoid heart disease with rheumatoid arthritis of right elbow
C2889204|Rheumatoid heart disease w rheumatoid arthritis of r elbow
C2889205|Rheumatoid heart disease with rheumatoid arthritis of left elbow
C2889205|Rheumatoid heart disease w rheumatoid arthritis of l elbow
C2889206|Rheumatoid heart disease with rheumatoid arthritis of unspecified elbow
C2889206|Rheu heart disease w rheumatoid arthritis of unsp elbow
C2889209|Rheumatoid heart disease with rheumatoid arthritis of right wrist
C2889209|Rheumatoid heart disease w rheumatoid arthritis of r wrist
C2889210|Rheumatoid heart disease with rheumatoid arthritis of left wrist
C2889210|Rheumatoid heart disease w rheumatoid arthritis of l wrist
C2889211|Rheumatoid heart disease with rheumatoid arthritis of unspecified wrist
C2889211|Rheu heart disease w rheumatoid arthritis of unsp wrist
C2889214|Rheumatoid heart disease with rheumatoid arthritis of right hand
C2889214|Rheu heart disease w rheumatoid arthritis of right hand
C2889215|Rheumatoid heart disease with rheumatoid arthritis of left hand
C2889215|Rheumatoid heart disease w rheumatoid arthritis of left hand
C2889216|Rheumatoid heart disease with rheumatoid arthritis of unspecified hand
C2889216|Rheumatoid heart disease w rheumatoid arthritis of unsp hand
C2889218|Rheumatoid heart disease with rheumatoid arthritis of right hip
C2889218|Rheumatoid heart disease w rheumatoid arthritis of right hip
C2889219|Rheumatoid heart disease with rheumatoid arthritis of left hip
C2889219|Rheumatoid heart disease w rheumatoid arthritis of left hip
C2889221|Rheumatoid heart disease with rheumatoid arthritis of right knee
C2889221|Rheu heart disease w rheumatoid arthritis of right knee
C2889222|Rheumatoid heart disease with rheumatoid arthritis of left knee
C2889222|Rheumatoid heart disease w rheumatoid arthritis of left knee
C2889223|Rheumatoid heart disease with rheumatoid arthritis of unspecified knee
C2889223|Rheumatoid heart disease w rheumatoid arthritis of unsp knee
C2889226|Rheumatoid heart disease with rheumatoid arthritis of right ankle and foot
C2889226|Rheu heart disease w rheumatoid arthritis of right ank/ft
C2889227|Rheumatoid heart disease with rheumatoid arthritis of left ankle and foot
C2889227|Rheu heart disease w rheumatoid arthritis of left ank/ft
C2889228|Rheumatoid heart disease with rheumatoid arthritis of unspecified ankle and foot
C2889228|Rheu heart disease w rheumatoid arthritis of unsp ank/ft
C2889231|Rheumatoid myopathy with rheumatoid arthritis of unspecified site
C2889231|Rheumatoid myopathy with rheumatoid arthritis of unsp site
C2889232|Rheumatoid myopathy with rheumatoid arthritis of shoulder
C2889236|Rheumatoid myopathy with rheumatoid arthritis of elbow
C2889241|Rheumatoid myopathy with rheumatoid arthritis of wrist
C2889246|Rheumatoid myopathy with rheumatoid arthritis of hand
C2889246|Rheumatoid myopathy with rheumatoid arthritis of unspecified hand
C2889246|Rheumatoid myopathy with rheumatoid arthritis of unsp hand
C2889249|Rheumatoid myopathy with rheumatoid arthritis of hip
C2889253|Rheumatoid myopathy with rheumatoid arthritis of knee
C2889258|Rheumatoid myopathy with rheumatoid arthritis of ankle and foot
C2889262|Rheumatoid myopathy with rheumatoid arthritis of multiple sites
C2889262|Rheumatoid myopathy w rheumatoid arthritis of multiple sites
C2889233|Rheumatoid myopathy with rheumatoid arthritis of right shoulder
C2889233|Rheumatoid myopathy w rheumatoid arthritis of right shoulder
C2889234|Rheumatoid myopathy with rheumatoid arthritis of left shoulder
C2889234|Rheumatoid myopathy w rheumatoid arthritis of left shoulder
C2889235|Rheumatoid myopathy with rheumatoid arthritis of unspecified shoulder
C2889235|Rheumatoid myopathy w rheumatoid arthritis of unsp shoulder
C2889237|Rheumatoid myopathy with rheumatoid arthritis of right elbow
C2889238|Rheumatoid myopathy with rheumatoid arthritis of left elbow
C2889239|Rheumatoid myopathy with rheumatoid arthritis of unspecified elbow
C2889239|Rheumatoid myopathy with rheumatoid arthritis of unsp elbow
C2889242|Rheumatoid myopathy with rheumatoid arthritis of right wrist
C2889243|Rheumatoid myopathy with rheumatoid arthritis of left wrist
C2889244|Rheumatoid myopathy with rheumatoid arthritis of unspecified wrist
C2889244|Rheumatoid myopathy with rheumatoid arthritis of unsp wrist
C2889247|Rheumatoid myopathy with rheumatoid arthritis of right hand
C2889248|Rheumatoid myopathy with rheumatoid arthritis of left hand
C2889250|Rheumatoid myopathy with rheumatoid arthritis of right hip
C2889251|Rheumatoid myopathy with rheumatoid arthritis of left hip
C2889252|Rheumatoid myopathy with rheumatoid arthritis of unspecified hip
C2889252|Rheumatoid myopathy with rheumatoid arthritis of unsp hip
C2889254|Rheumatoid myopathy with rheumatoid arthritis of right knee
C2889255|Rheumatoid myopathy with rheumatoid arthritis of left knee
C2889256|Rheumatoid myopathy with rheumatoid arthritis of unspecified knee
C2889256|Rheumatoid myopathy with rheumatoid arthritis of unsp knee
C2889259|Rheumatoid myopathy with rheumatoid arthritis of right ankle and foot
C2889259|Rheumatoid myopathy w rheumatoid arthritis of right ank/ft
C2889260|Rheumatoid myopathy with rheumatoid arthritis of left ankle and foot
C2889260|Rheumatoid myopathy w rheumatoid arthritis of left ank/ft
C2889261|Rheumatoid myopathy with rheumatoid arthritis of unspecified ankle and foot
C2889261|Rheumatoid myopathy w rheumatoid arthritis of unsp ank/ft
C2889264|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified site
C2889264|Rheumatoid polyneurop w rheumatoid arthritis of unsp site
C2889265|Rheumatoid polyneuropathy with rheumatoid arthritis of shoulder
C2889271|Rheumatoid polyneuropathy with rheumatoid arthritis of elbow
C2889271|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified elbow
C2889271|Rheumatoid polyneurop w rheumatoid arthritis of unsp elbow
C2889273|Rheumatoid polyneuropathy with rheumatoid arthritis of wrist
C2889278|Rheumatoid polyneuropathy with rheumatoid arthritis of hand
C2889282|Rheumatoid polyneuropathy with rheumatoid arthritis of hip
C2889286|Rheumatoid polyneuropathy with rheumatoid arthritis of knee
C2889291|Rheumatoid polyneuropathy with rheumatoid arthritis of ankle and foot
C2889295|Rheumatoid polyneuropathy with rheumatoid arthritis of multiple sites
C2889295|Rheumatoid polyneuropathy w rheumatoid arthritis mult site
C2889266|Rheumatoid polyneuropathy with rheumatoid arthritis of right shoulder
C2889266|Rheumatoid polyneurop w rheumatoid arthritis of r shoulder
C2889267|Rheumatoid polyneuropathy with rheumatoid arthritis of left shoulder
C2889267|Rheumatoid polyneurop w rheumatoid arthritis of l shoulder
C2889268|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified shoulder
C2889268|Rheu polyneurop w rheumatoid arthritis of unsp shoulder
C2889269|Rheumatoid polyneuropathy with rheumatoid arthritis of right elbow
C2889269|Rheumatoid polyneurop w rheumatoid arthritis of right elbow
C2889270|Rheumatoid polyneuropathy with rheumatoid arthritis of left elbow
C2889270|Rheumatoid polyneurop w rheumatoid arthritis of left elbow
C2889274|Rheumatoid polyneuropathy with rheumatoid arthritis of right wrist
C2889274|Rheumatoid polyneurop w rheumatoid arthritis of right wrist
C2889275|Rheumatoid polyneuropathy with rheumatoid arthritis of left wrist
C2889275|Rheumatoid polyneurop w rheumatoid arthritis of left wrist
C2889276|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified wrist
C2889276|Rheumatoid polyneurop w rheumatoid arthritis of unsp wrist
C2889279|Rheumatoid polyneuropathy with rheumatoid arthritis of right hand
C2889279|Rheumatoid polyneurop w rheumatoid arthritis of right hand
C2889280|Rheumatoid polyneuropathy with rheumatoid arthritis of left hand
C2889280|Rheumatoid polyneurop w rheumatoid arthritis of left hand
C2889281|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified hand
C2889281|Rheumatoid polyneurop w rheumatoid arthritis of unsp hand
C2889283|Rheumatoid polyneuropathy with rheumatoid arthritis of right hip
C2889283|Rheumatoid polyneurop w rheumatoid arthritis of right hip
C2889284|Rheumatoid polyneuropathy with rheumatoid arthritis of left hip
C2889284|Rheumatoid polyneuropathy w rheumatoid arthritis of left hip
C2889285|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified hip
C2889285|Rheumatoid polyneuropathy w rheumatoid arthritis of unsp hip
C2889287|Rheumatoid polyneuropathy with rheumatoid arthritis of right knee
C2889287|Rheumatoid polyneurop w rheumatoid arthritis of right knee
C2889288|Rheumatoid polyneuropathy with rheumatoid arthritis of left knee
C2889288|Rheumatoid polyneurop w rheumatoid arthritis of left knee
C2889289|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified knee
C2889289|Rheumatoid polyneurop w rheumatoid arthritis of unsp knee
C2889292|Rheumatoid polyneuropathy with rheumatoid arthritis of right ankle and foot
C2889292|Rheumatoid polyneurop w rheumatoid arthritis of right ank/ft
C2889293|Rheumatoid polyneuropathy with rheumatoid arthritis of left ankle and foot
C2889293|Rheumatoid polyneurop w rheumatoid arthritis of left ank/ft
C2889294|Rheumatoid polyneuropathy with rheumatoid arthritis of unspecified ankle and foot
C2889294|Rheumatoid polyneurop w rheumatoid arthritis of unsp ank/ft
C2889297|Rheumatoid arthritis of right shoulder with involvement of other organs and systems
C2889297|Rheu arthritis of r shoulder w involv of organs and systems
C2889298|Rheumatoid arthritis of left shoulder with involvement of other organs and systems
C2889298|Rheu arthritis of l shoulder w involv of organs and systems
C2889299|Rheumatoid arthritis of unspecified shoulder with involvement of other organs and systems
C2889299|Rheu arthrit of unsp shoulder w involv of organs and systems
C2889301|Rheumatoid arthritis of right elbow with involvement of other organs and systems
C2889301|Rheu arthritis of r elbow w involv of organs and systems
C2889302|Rheumatoid arthritis of left elbow with involvement of other organs and systems
C2889302|Rheu arthritis of l elbow w involv of organs and systems
C2889303|Rheumatoid arthritis of unspecified elbow with involvement of other organs and systems
C2889303|Rheu arthritis of unsp elbow w involv of organs and systems
C2889306|Rheumatoid arthritis of right wrist with involvement of other organs and systems
C2889306|Rheu arthritis of r wrist w involv of organs and systems
C2889307|Rheumatoid arthritis of left wrist with involvement of other organs and systems
C2889307|Rheu arthritis of l wrist w involv of organs and systems
C2889308|Rheumatoid arthritis of unspecified wrist with involvement of other organs and systems
C2889308|Rheu arthritis of unsp wrist w involv of organs and systems
C2889314|Rheumatoid arthritis of right hip with involvement of other organs and systems
C2889314|Rheu arthritis of right hip w involv of organs and systems
C2889315|Rheumatoid arthritis of left hip with involvement of other organs and systems
C2889315|Rheu arthritis of left hip w involv of organs and systems
C2889316|Rheumatoid arthritis of unspecified hip with involvement of other organs and systems
C2889316|Rheu arthritis of unsp hip w involv of organs and systems
C2889318|Rheumatoid arthritis of right knee with involvement of other organs and systems
C2889318|Rheu arthritis of right knee w involv of organs and systems
C2889319|Rheumatoid arthritis of left knee with involvement of other organs and systems
C2889319|Rheu arthritis of left knee w involv of organs and systems
C2889320|Rheumatoid arthritis of unspecified knee with involvement of other organs and systems
C2889320|Rheu arthritis of unsp knee w involv of organs and systems
C2889326|Rheumatoid arthritis with rheumatoid factor of unspecified site without organ or systems involvement
C2889326|Rheu arthritis w rheu factor of unsp site w/o org/sys involv
C2889327|Rheumatoid arthritis with rheumatoid factor of shoulder without organ or systems involvement
C2889331|Rheumatoid arthritis with rheumatoid factor of elbow without organ or systems involvement
C2889335|Rheumatoid arthritis with rheumatoid factor of wrist without organ or systems involvement
C2889339|Rheumatoid arthritis with rheumatoid factor of hand without organ or systems involvement
C2889343|Rheumatoid arthritis with rheumatoid factor of hip without organ or systems involvement
C2889347|Rheumatoid arthritis with rheumatoid factor of knee without organ or systems involvement
C2889351|Rheumatoid arthritis with rheumatoid factor of ankle and foot without organ or systems involvement
C2889355|Rheumatoid arthritis with rheumatoid factor of multiple sites without organ or systems involvement
C2889355|Rheu arthritis w rheu factor mult site w/o org/sys involv
C2889328|Rheumatoid arthritis with rheumatoid factor of right shoulder without organ or systems involvement
C2889328|Rheu arthrit w rheu factor of r shoulder w/o org/sys involv
C2889329|Rheumatoid arthritis with rheumatoid factor of left shoulder without organ or systems involvement
C2889329|Rheu arthrit w rheu factor of l shoulder w/o org/sys involv
C2889330|Rheumatoid arthritis with rheumatoid factor of unspecified shoulder without organ or systems involvement
C2889330|Rheu arthrit w rheu factor of unsp shldr w/o org/sys involv
C2889332|Rheumatoid arthritis with rheumatoid factor of right elbow without organ or systems involvement
C2889332|Rheu arthritis w rheu factor of r elbow w/o org/sys involv
C2889333|Rheumatoid arthritis with rheumatoid factor of left elbow without organ or systems involvement
C2889333|Rheu arthritis w rheu factor of l elbow w/o org/sys involv
C2889334|Rheumatoid arthritis with rheumatoid factor of unspecified elbow without organ or systems involvement
C2889334|Rheu arthrit w rheu factor of unsp elbow w/o org/sys involv
C2889336|Rheumatoid arthritis with rheumatoid factor of right wrist without organ or systems involvement
C2889336|Rheu arthritis w rheu factor of r wrist w/o org/sys involv
C2889337|Rheumatoid arthritis with rheumatoid factor of left wrist without organ or systems involvement
C2889337|Rheu arthritis w rheu factor of l wrist w/o org/sys involv
C2889338|Rheumatoid arthritis with rheumatoid factor of unspecified wrist without organ or systems involvement
C2889338|Rheu arthrit w rheu factor of unsp wrist w/o org/sys involv
C2889340|Rheumatoid arthritis with rheumatoid factor of right hand without organ or systems involvement
C2889340|Rheu arthritis w rheu factor of r hand w/o org/sys involv
C2889341|Rheumatoid arthritis with rheumatoid factor of left hand without organ or systems involvement
C2889341|Rheu arthritis w rheu factor of left hand w/o org/sys involv
C2889342|Rheumatoid arthritis with rheumatoid factor of unspecified hand without organ or systems involvement
C2889342|Rheu arthritis w rheu factor of unsp hand w/o org/sys involv
C2889344|Rheumatoid arthritis with rheumatoid factor of right hip without organ or systems involvement
C2889344|Rheu arthritis w rheu factor of right hip w/o org/sys involv
C2889345|Rheumatoid arthritis with rheumatoid factor of left hip without organ or systems involvement
C2889345|Rheu arthritis w rheu factor of left hip w/o org/sys involv
C2889346|Rheumatoid arthritis with rheumatoid factor of unspecified hip without organ or systems involvement
C2889346|Rheu arthritis w rheu factor of unsp hip w/o org/sys involv
C2889348|Rheumatoid arthritis with rheumatoid factor of right knee without organ or systems involvement
C2889348|Rheu arthritis w rheu factor of r knee w/o org/sys involv
C2889349|Rheumatoid arthritis with rheumatoid factor of left knee without organ or systems involvement
C2889349|Rheu arthritis w rheu factor of left knee w/o org/sys involv
C2889350|Rheumatoid arthritis with rheumatoid factor of unspecified knee without organ or systems involvement
C2889350|Rheu arthritis w rheu factor of unsp knee w/o org/sys involv
C2889352|Rheumatoid arthritis with rheumatoid factor of right ankle and foot without organ or systems involvement
C2889352|Rheu arthrit w rheu fctr of right ank/ft w/o org/sys involv
C2889353|Rheumatoid arthritis with rheumatoid factor of left ankle and foot without organ or systems involvement
C2889353|Rheu arthrit w rheu factor of left ank/ft w/o org/sys involv
C2889354|Rheumatoid arthritis with rheumatoid factor of unspecified ankle and foot without organ or systems involvement
C2889354|Rheu arthrit w rheu factor of unsp ank/ft w/o org/sys involv
C2889356|Other rheumatoid arthritis with rheumatoid factor
C2889356|Other rheumatoid arthritis with rheumatoid factor of unspecified site
C2889356|Oth rheumatoid arthritis with rheumatoid factor of unsp site
C2889357|Other rheumatoid arthritis with rheumatoid factor of shoulder
C2889361|Other rheumatoid arthritis with rheumatoid factor of elbow
C2889365|Other rheumatoid arthritis with rheumatoid factor of wrist
C2889371|Other rheumatoid arthritis with rheumatoid factor of hand
C2889371|Other rheumatoid arthritis with rheumatoid factor of unspecified hand
C2889371|Oth rheumatoid arthritis with rheumatoid factor of unsp hand
C2889372|Other rheumatoid arthritis with rheumatoid factor of hip
C2889376|Other rheumatoid arthritis with rheumatoid factor of knee
C2889380|Other rheumatoid arthritis with rheumatoid factor of ankle and foot
C2889384|Other rheumatoid arthritis with rheumatoid factor of multiple sites
C2889384|Oth rheumatoid arthritis w rheumatoid factor mult site
C2889358|Other rheumatoid arthritis with rheumatoid factor of right shoulder
C2889358|Oth rheumatoid arthritis w rheumatoid factor of r shoulder
C2889359|Other rheumatoid arthritis with rheumatoid factor of left shoulder
C2889359|Oth rheumatoid arthritis w rheumatoid factor of l shoulder
C2889360|Other rheumatoid arthritis with rheumatoid factor of unspecified shoulder
C2889360|Oth rheu arthritis w rheumatoid factor of unsp shoulder
C2889362|Other rheumatoid arthritis with rheumatoid factor of right elbow
C2889362|Oth rheumatoid arthritis w rheumatoid factor of right elbow
C2889363|Other rheumatoid arthritis with rheumatoid factor of left elbow
C2889363|Oth rheumatoid arthritis w rheumatoid factor of left elbow
C2889364|Other rheumatoid arthritis with rheumatoid factor of unspecified elbow
C2889364|Oth rheumatoid arthritis w rheumatoid factor of unsp elbow
C2889366|Other rheumatoid arthritis with rheumatoid factor of right wrist
C2889366|Oth rheumatoid arthritis w rheumatoid factor of right wrist
C2889367|Other rheumatoid arthritis with rheumatoid factor of left wrist
C2889367|Oth rheumatoid arthritis w rheumatoid factor of left wrist
C2889368|Other rheumatoid arthritis with rheumatoid factor of unspecified wrist
C2889368|Oth rheumatoid arthritis w rheumatoid factor of unsp wrist
C2889369|Other rheumatoid arthritis with rheumatoid factor of right hand
C2889369|Oth rheumatoid arthritis w rheumatoid factor of right hand
C2889370|Other rheumatoid arthritis with rheumatoid factor of left hand
C2889370|Oth rheumatoid arthritis with rheumatoid factor of left hand
C2889373|Other rheumatoid arthritis with rheumatoid factor of right hip
C2889373|Oth rheumatoid arthritis with rheumatoid factor of right hip
C2889374|Other rheumatoid arthritis with rheumatoid factor of left hip
C2889374|Oth rheumatoid arthritis with rheumatoid factor of left hip
C2889375|Other rheumatoid arthritis with rheumatoid factor of unspecified hip
C2889375|Oth rheumatoid arthritis with rheumatoid factor of unsp hip
C2889377|Other rheumatoid arthritis with rheumatoid factor of right knee
C2889377|Oth rheumatoid arthritis w rheumatoid factor of right knee
C2889378|Other rheumatoid arthritis with rheumatoid factor of left knee
C2889378|Oth rheumatoid arthritis with rheumatoid factor of left knee
C2889379|Other rheumatoid arthritis with rheumatoid factor of unspecified knee
C2889379|Oth rheumatoid arthritis with rheumatoid factor of unsp knee
C2889381|Other rheumatoid arthritis with rheumatoid factor of right ankle and foot
C2889381|Oth rheumatoid arthritis w rheumatoid factor of right ank/ft
C2889382|Other rheumatoid arthritis with rheumatoid factor of left ankle and foot
C2889382|Oth rheumatoid arthritis w rheumatoid factor of left ank/ft
C2889383|Other rheumatoid arthritis with rheumatoid factor of unspecified ankle and foot
C2889383|Oth rheumatoid arthritis w rheumatoid factor of unsp ank/ft
C2889197|Rheumatoid heart disease with rheumatoid arthritis
C2889197|rheumatoid heart disease with rheumatoid arthritis (diagnosis)
C2889230|Rheumatoid myopathy with rheumatoid arthritis
C2889263|Rheumatoid polyneuropathy with rheumatoid arthritis
C2889325|Rheumatoid arthritis with rheumatoid factor without organ or systems involvement
