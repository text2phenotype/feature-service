C0010403|Cryoglobulinemia
C0543697|Mixed cryoglobulinemia
C0543697|Mixed cryoglobulinaemia
C0010403|Cryoglobulinemia
C0010403|Cryoglobulinemias
C0010403|Cryoglobulinaemia
C0010403|cryoglobulinemia (diagnosis)
C0010403|Cryoglobulinemia [Disease/Finding]
C0010403|Cryoglobulinemia (disorder)
C0010403|Cryoimmunoglobulinaemia
C0010403|Cryoimmunoglobulinemia
C0010403|Cryoglobulinemia, NOS
C0010403|Cryoimmunoglobulinemia, NOS
C0010403|Cryoglobulinaemia, NOS
C0340992|cryoglobulinemic vasculitis (diagnosis)
C0340992|cryoglobulinemic vasculitis
C0340992|Cryoglobulinaemic vasculitis
C0340992|Cryoglobulinemic vasculitis (disorder)
C0340992|cryoglobulinemic; vasculitis
C0340992|vasculitis; cryoglobulinemic
C0340979|cryoglobulinemic purpura
C0340979|cryoglobulinemic purpura (diagnosis)
C0340979|Cryoglobulinaemic purpura
C0340979|Cryoglobulinemic purpura (disorder)
C0340979|cryoglobulinemic; purpura
C0340979|purpura; cryoglobulinemic
C0343208|mixed essential cryoglobulinemia (diagnosis)
C0343208|mixed essential cryoglobulinemia
C0343208|Essential mixed cryoglobulinemia
C0343208|Essential mixed cryoglobulinaemia
C0343208|Essential cryoglobulinaemic vasculitis
C0343208|Essential cryoglobulinemic vasculitis
C0343208|Essential mixed cryoglobulinemia (disorder)
C0272263|Cryofibrinogenemia
C0272263|Cryofibrinogenaemia
C0272263|Cryofibrinogenemia (disorder)
C0272263|Cryofibrinogenemia, NOS
C1852456|CRYOGLOBULINEMIA, FAMILIAL MIXED
C1852456|Meltzer Syndrome
C1852457|CRYOFIBRINOGENEMIA, FAMILIAL PRIMARY
C0272261|Mixed cryoimmunoglobulinemia with monoclonal component
C0272261|Mixed cryoimmunoglobulinaemia with monoclonal component
C0272261|Mixed cryoimmunoglobulinemia with monoclonal component (disorder)
C0272262|Mixed polyclonal cryoimmunoglobulinemia
C0272262|Mixed polyclonal cryoimmunoglobulinaemia
C0272262|Mixed polyclonal cryoimmunoglobulinemia (disorder)
C0272260|Monoclonal cryoimmunoglobulinemia
C0272260|Monoclonal cryoimmunoglobulinaemia
C0272260|Monoclonal cryoimmunoglobulinemia (disorder)
C0272258|Primary cryoglobulinemia
C0272258|Primary cryoglobulinaemia
C0272258|Primary cryoglobulinemia (disorder)
C0272259|Secondary cryoglobulinemia
C0272259|Secondary cryoglobulinaemia
C0272259|Secondary cryoglobulinemia (disorder)
C1384927|disease (or disorder); glomerular, in cryoglobulinemia (etiology)
C1384927|disease (or disorder); glomerular, in cryoglobulinemia (manifestation)
C1394252|cryoglobulinemia; with lung involvement (etiology)
C1394252|cryoglobulinemia; with lung involvement (manifestation)
C1394252|disease (or disorder); lung, in cryoglobulinemia (etiology)
C1394252|disease (or disorder); lung, in cryoglobulinemia (manifestation)
C1394252|lung; cryoglobulinemia (etiology)
C1394252|lung; cryoglobulinemia (manifestation)
C1394252|lung; disease, in cryoglobulinemia (manifestation)
C1385201|disease (or disorder); tubulo-interstitial, mixed cryoglobulinemia (etiology)
C1385201|disease (or disorder); tubulo-interstitial, mixed cryoglobulinemia (manifestation)
C1394251|cryoglobulinemia; glomerulonephritis (etiology)
C1394251|cryoglobulinemia; glomerulonephritis (manifestation)
C1394251|glomerulonephritis; cryoglobulinemia (etiology)
C1394251|glomerulonephritis; cryoglobulinemia (manifestation)
C1394253|cryoglobulinemia; pyelonephritis (etiology)
C1394253|cryoglobulinemia; pyelonephritis (manifestation)
C1394253|pyelonephritis; cryoglobulinemia (etiology)
C1394253|pyelonephritis; cryoglobulinemia (manifestation)
C1398770|glomerular; disease, in cryoglobulinemia (etiology)
C1398770|glomerular; disease, in cryoglobulinemia (manifestation)
C1407782|tubulo-interstitial; disease, mixed cryoglobulinemia (etiology)
C1407782|tubulo-interstitial; disease, mixed cryoglobulinemia (manifestation)
