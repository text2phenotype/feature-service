Quantity|equal|iso|||
Quantity|none|nulli|||none
Quantity|half|hemi||hemiplegia|half, partial
Quantity|half|semi||semilunar|half, partial
Quantity|one|primi||primigravida|first
Quantity|one|uni|||one
Quantity|one|mono||monocyte|one
Quantity|two|bi|||two
Quantity|two|di|||two
Quantity|two|diplo||diplopia|double
Quantity|two|dupli||duplication|double
Quantity|three|tri|||three
Quantity|four|quad||quadruple|four
Quantity|four|quadri||quadriplegia|four
Quantity|four|tetra||tetralogy|four
Quantity|poly|poly||polycystic|many, much, excessive, frequent
Quantity|all|pan|||all
Quantity|small|oligo||oligospermia|short
Quantity|small||icle|ventricle|small
Quantity|micro|micro||microscope|small, tiny
Quantity|milli|milli||millileter|thousandth
Quantity|large|macro||macroglossia|large
Quantity|large|mega||megacolon|big
Quantity|large|maxim||maximum|max
Quantity|ultra|ultra||ultrasound|beyond, excessive

