C0002210|alpha-Fetoproteins
C0201539|Alpha one fetoprotein measurement
C0002210|alpha Fetoprotein
C0002210|alpha Fetoproteins
C0002210|alpha-Fetoproteins
C0002210|fetuin
C0002210|alpha Foetoprotein
C0002210|alpha-Fetoprotein
C0002210|alpha-Fetoproteins [Chemical/Ingredient]
C0002210|Alpha-1-Fetoprotein
C0002210|AFP
C0002210|Alpha Fetal Protein
C0002210|AFP - Alpha-fetoprotein
C0002210|Fetuin (substance)
C0002210|alpha Fetoprotein (substance)
C0002210|Alpha-Fetoglobulin
C2717473|AFPep peptide
C2717473|TOVNO peptide
C2742043|alpha-fetoprotein related protein, mouse
C2742043|ARG protein, mouse
C2975076|growth inhibitory peptide-34, human
C2975076|GIP-34 peptide, human
C1863081|alpha-Fetoprotein Deficiency
C1863081|AFPD
C1981150|Alpha-1-fetoprotein &#x7C; amniotic fluid
C2600377|Alpha-1-Fetoprotein &#x7C; Blood cord
C1981155|Alpha-1-fetoprotein &#x7C; Peritoneal fluid
C1981152|Alpha-1-fetoprotein &#x7C; body fluid
C1981160|Alpha-1-fetoprotein L3 &#x7C; bld-ser-plas
C1981153|Alpha-1-fetoprotein &#x7C; cerebral spinal fluid
C1981151|Alpha-1-fetoprotein &#x7C; bld-ser-plas
C2600378|Alpha-1-Fetoprotein.tumor marker &#x7C; Bld-Ser-Plas
C1981156|Alpha-1-fetoprotein &#x7C; pleural fluid
C1648292|Alpha-1-Fetoprotein.L3
C1648292|alpha Fetoprotein, L3
C1648292|Alpha-fetoprotein, L3
C1648292|alpha Fetoprotein, L3 (substance)
C1648292|Alpha-1-fetoprotein, L3
C0612946|ALF-DTPA
C0612946|asialofetuin-DTPA complex
C0059058|embryonin
C0623170|Ep-459-AF
C0623170|Ep 459-asialofetuin conjugate
C0623170|asialofetuin-Ep 459
C0636374|Thr-Leu-His-N-methylamide
C0636374|threonyl-leucyl-histidine-N-methylamide
C0641482|asialofetuin-polylysine-5'-uridine monophosphate conjugate
C0641482|AsF-PL-UMP
C0655320|PEG modified asialofetuin
C0655320|PEG-asialofetuin
C0655320|polyethylene glycol-asialofetuin complex
C0251381|AsF12 peptide
C0251381|asialofetuin 12 peptide
C0251383|AsF 21-45 peptide
C0251383|asialofetuin 21-45 peptide
C0251385|AsF 69-28 peptide
C0251385|asialofetuin 69-28 peptide
C1435546|alpha-fetoprotein, rat
C1435546|Afp protein, rat
C1435546|alpha-fetospecific glycoprotein, rat
C1435546|AF glycoprotein, rat
C1569245|P149 protein, human
C1307640|AFP protein, human
C1307640|alpha-fetoprotein, human
C1307640|alpha-fetospecific glycoprotein, human
C1307640|alpha-glycoprotein, fetospecific, human
C1307640|glycosylated AFP protein, human
C1307640|AF glycoprotein, human
C0201539|AFP
C0201539|Alpha 1 foetoprotein
C0201539|AFP Alphafoetoprotein
C0201539|Alpha-fetoprotein Measurement
C0201539|Alpha-1-Foetoprotein measurement
C0201539|Alpha Foetoprotein measurement
C0201539|Alpha one fetoprotein measurement
C0201539|Test;alpha fetoprotein
C0201539|Alpha-fetoprotein NOS
C0201539|Alpha-fetoprotein NOS (procedure)
C0201539|Alpha-fetoprotein (AFP)
C0201539|Alpha Fetoprotein
C0201539|Alpha-1-Fetoprotein Measurement
C0201539|Alphafetoprotein
C0201539|Alpha 1 fetoprotein
C0201539|Alphafoetoprotein
C0201539|AFP measurement
C0201539|Alpha Fetoprotein measurement
C0201539|Alpha-1-Fetoprotein measurement (procedure)
C0201539|alpha fetoprotein test
C2711551|Measurement of alpha fetoprotein as marker for malignant neoplasm (procedure)
C2711551|Measurement of alpha fetoprotein as marker for malignant neoplasm
C2711939|Measurement of alpha fetoprotein in second trimester
C2711939|Measurement of alpha fetoprotein in second trimester (procedure)
C2368140|body fluid alpha-fetoprotein
C2368140|body fluid AFP
C2368140|body fluid alpha-fetoprotein measurement
C2368140|body fluid alpha-fetoprotein measurement (lab test)
C3272858|Alpha-fetoprotein Ratio Measurement
C3272862|Alpha Fetoprotein L1 Measurement
C3272862|Alpha Fetoprotein L1
C3272862|AFPL1
C3272863|Alpha Fetoprotein L2 Measurement
C3272863|Alpha Fetoprotein L2
C3272863|AFPL2
C3272864|Alpha Fetoprotein L3 Measurement
C3272864|Alpha Fetoprotein L3
C3272864|AFPL3
C2210854|alpha-fetoprotein tetra profile
C2210854|alpha-fetoprotein tetra profile (lab test)
C2210854|prenatal maternal AFP quad screen
C0546833|Alpha-fetoprotein (AFP); serum
C0546833|serum alpha-fetoprotein measurement (lab test)
C0546833|serum AFP
C0546833|serum alpha-fetoprotein
C0546833|serum alpha-fetoprotein measurement
C0546833|serum alpha-fetoprotein (AFP) measurement
C0546833|ALPHA-FETOPROTEIN SERUM
C0546833|Alpha-fetoprotein (AFP) level, serum
C0546833|Measurement of alpha-fetoprotein (AFP) in serum
C0546833|Alpha-fetoprotein (AFP) level, serum"
C1740749|Alpha-fetoprotein (AFP); AFP-L3 fraction isoform and total AFP (including ratio)
C1740749|ALPHA-FETOPROTEIN L3
C1740749|AFP-L3 FRACTION ISOFORM & TOTAL AFP W/RATIO
C1740749|Measurement of alpha fetoprotein-L3 fraction isoform and total alpha-fetoprotein with ratio
C3714538|Alpha-fetoprotein (AFP); amniotic fluid
C3714538|amniotic fluid alpha-fetoprotein
C3714538|amniotic fluid alpha-fetoprotein measurement (lab test)
C3714538|amniotic fluid alpha-fetoprotein measurement
C3714538|amniotic fluid AFP measurement
C3714538|ALPHA-FETOPROTEIN AMNIOTIC
C3714538|ALPHA-FETOPROTEIN AMNIOTIC FLUID
C3714538|Alpha-fetoprotein (AFP) level, amniotic fluid
C3714538|Measurement of alpha-fetoprotein (AFP) in amniotic fluid
C3714538|Amniotic fluid AFP NOS
C3714538|Amniotic fluid AFP NOS (procedure)
C3714538|Amniotic fluid AFP
C3714538|Amniotic fluid AFP (procedure)
C3714538|Alphafetoprotein amniotic fluid
C3714538|Alphafoetoprotein amniotic fluid
C3714538|AFP amniotic fluid
C0428145|Alpha 1 foetoprotein amniotic fluid
C0428145|Alpha-1-Foetoprotein measurement, amniotic fluid
C0428145|amniotic fluid alpha-1-fetoprotein (lab test)
C0428145|amniotic fluid alpha-1-fetoprotein
C0428145|Alpha 1 fetoprotein amniotic fluid
C0428145|Alpha-1-Fetoprotein measurement, amniotic fluid
C0428145|Alpha-1-Fetoprotein measurement, amniotic fluid (procedure)
C1446076|cerebrospinal fluid alpha fetoprotein measurement (lab test)
C1446076|CSF alpha fetoprotein measurement
C1446076|cerebrospinal fluid alpha fetoprotein measurement
C1446076|CSF AFP level
C1446076|Alpha-1-Foetoprotein measurement, spinal fluid
C1446076|ASV measurement
C1446076|Alpha-1-Fetoprotein measurement, spinal fluid
C1446076|Alpha-1-Fetoprotein measurement, spinal fluid (procedure)
C1446076|Cerebrospinal fluid alpha-fetoprotein measurement (procedure)
C1446076|Cerebrospinal fluid alpha-fetoprotein measurement
C0419584|Alpha-fetoprotein blood test
C0419584|Alpha-fetoprotein blood test (procedure)
C1271788|Fluid sample AFP level (procedure)
C1271788|Fluid sample alpha fetoprotein level
C1271788|Fluid sample alpha fetoprotein level (procedure)
C1271788|Fluid sample AFP level
C1271652|MS alpha-fetoprotein level (procedure)
C1271652|Maternal serum (MS) alpha-fetoprotein level
C1271652|Maternal serum alpha-fetoprotein level (procedure)
C1271652|Maternal serum alpha-fetoprotein level
C1271652|Maternal serum (MS) alpha-fetoprotein level (procedure)
C1271652|MS alpha-fetoprotein level
C1271652|MSAFP level
C1271652|Maternal serum alpha fetoprotein level
C1278027|Plasma alpha-fetoprotein multiple of median measurement (procedure)
C1278027|Plasma AFP mean of median measurement
C1278027|Plasma alpha-fetoprotein multiple of median measurement
C1278027|Plasma alpha-fetoprotein (AFP) multiple of median measurement
C1278027|Plasma AFP mean of median measurement (procedure)
C1278027|Plasma AFP MoM
C1278027|Plasma AFP MoM (procedure)
C0856296|Screening neural tube defect (maternal serum AFP)
