C0270611|Brain Injuries
C0347535|Intracranial injury
C0006109|Brain Damage, Chronic
C0019151|Hepatic Encephalopathy
C0006107|Concussion
C0006107|Brain Concussion
C0006107|Brain Concussions
C0006107|Concussion, Brain
C0006107|concussion (diagnosis)
C0006107|Cerebral Concussions
C0006107|Concussion, Cerebral
C0006107|Concussion NOS
C0006107|Commotio cerebri
C0006107|Brain Concussion [Disease/Finding]
C0006107|Cerebral Concussion
C0006107|Concussion (disorder)
C0006107|Concussion NOS (disorder)
C0006107|concussion injury of brain (diagnosis)
C0006107|Concussion injury of brain
C0006107|Brain--Concussion
C0006107|Mild traumatic brain injury
C0006107|MTBI - Mild traumatic brain injury
C0006107|Commotio
C0006107|Concussion, unspecified
C0006107|Neuro: Concussion
C0006107|Concussion injury of brain (disorder)
C0006107|brain; blast
C0006107|brain; commotio
C0006107|brain; concussion
C0006107|cerebral; concussion
C0006107|cerebri; commotio
C0006107|commotio; brain
C0006107|concussion; brain
C0006107|concussion; cerebral
C0006107|Concussion (Brain)
C0006107|Injury;concussion;head
C0852861|Brain damage (excluding perinatal)
C0852861|Brain damage (excl perinatal)
C0014557|Epilepsies, Post-Traumatic
C0014557|Epilepsies, Traumatic
C0014557|Epilepsy, Post Traumatic
C0014557|Epilepsy, Post-Traumatic
C0014557|Post-Traumatic Epilepsies
C0014557|Post-Traumatic Epilepsy
C0014557|Traumatic Epilepsies
C0014557|Traumatic Epilepsy
C0014557|SEIZURE DIS POST TRAUMATIC
C0014557|POST TRAUMATIC SEIZURE DIS
C0014557|Disorder, Post-Traumatic Seizure
C0014557|Disorders, Post-Traumatic Seizure
C0014557|Post Traumatic Seizure Disorder
C0014557|Post-Traumatic Seizure Disorders
C0014557|Seizure Disorder, Post Traumatic
C0014557|Seizure Disorders, Post-Traumatic
C0014557|Epilepsy, Post-Traumatic [Disease/Finding]
C0014557|Post-Traumatic Seizure Disorder
C0014557|Epilepsy, Traumatic
C0014557|Seizure Disorder, Post-Traumatic
C0014557|Traumatic epilepsy (disorder)
C0014557|PTE - Post-traumatic epilepsy
C0014557|Post-traumatic epilepsy (disorder)
C0014557|epilepsy; traumatic
C0014557|traumatic; epileptic
C0032268|Pneumocephalus
C0032268|Airocele, Cranial
C0032268|Airoceles, Cranial
C0032268|Cranial Airoceles
C0032268|Pneumocyst, Cranial
C0032268|Cranial Pneumocysts
C0032268|Pneumocysts, Cranial
C0032268|Gas, Intracranial
C0032268|Cranial Airocele
C0032268|Cranial Pneumocyst
C0032268|Pneumocephalus [Disease/Finding]
C0032268|Intracranial Gas
C0032268|Airocoele
C0032268|Airocele
C0032268|Pneumocephalus (disorder)
C0751799|Brain Hemorrhage, Traumatic
C0751799|Brain Hemorrhages, Traumatic
C0751799|Hemorrhage, Traumatic Brain
C0751799|Traumatic Brain Hemorrhages
C0751799|Brain Hemorrhage, Traumatic [Disease/Finding]
C0751799|Traumatic Brain Hemorrhage
C0751799|brain; hemorrhage, traumatic
C0751799|hemorrhage; brain, traumatic
C0751813|BRAIN INJ CHRONIC
C0751813|CHRONIC BRAIN INJ
C0751813|ENCEPHALOPATHY POSTTRAUMATIC CHRONIC
C0751813|TRAUMATIC ENCEPH CHRONIC
C0751813|INJ BRAIN CHRONIC
C0751813|ENCEPH POST TRAUMATIC CHRONIC
C0751813|CHRONIC POST TRAUMATIC ENCEPH
C0751813|Brain Injuries, Chronic
C0751813|Brain Injury, Chronic
C0751813|Chronic Brain Injuries
C0751813|Chronic Post Traumatic Encephalopathy
C0751813|Chronic Post-Traumatic Encephalopathies
C0751813|Encephalopathies, Chronic Post-Traumatic
C0751813|Encephalopathy, Chronic Post-Traumatic
C0751813|Post-Traumatic Encephalopathies, Chronic
C0751813|Post-Traumatic Encephalopathy, Chronic
C0751813|Chronic Traumatic Encephalopathy
C0751813|Encephalopathy, Chronic Traumatic
C0751813|Traumatic Encephalopathies, Chronic
C0751813|Brain Injury, Chronic [Disease/Finding]
C0751813|Chronic Brain Injury
C0751813|Traumatic Encephalopathy, Chronic
C0751813|Chronic Post-Traumatic Encephalopathy
C0751813|Encephalopathy, Post-Traumatic, Chronic
C0751813|Injury, Brain, Chronic
C0751813|chronic traumatic encephalopathy (diagnosis)
C0752219|Diffuse axonal injury
C0752219|DIFFUSE AXONAL INJ
C0752219|AXONAL INJ DIFFUSE
C0752219|Axonal Injuries, Diffuse
C0752219|Diffuse Axonal Injuries
C0752219|Injuries, Diffuse Axonal
C0752219|Injury, Diffuse Axonal
C0752219|DAI (Diffuse Axonal Injury)
C0752219|Axonal Injury, Diffuse
C0752219|Diffuse Axonal Injury [Disease/Finding]
C0752219|DAIs (Diffuse Axonal Injury)
C0686721|shaken infant syndrome (diagnosis)
C0686721|shaken infant syndrome
C0686721|Shaken Baby Syndrome
C0686721|Shaken Baby Syndrome [Disease/Finding]
C0686721|Shaken baby syndrome (finding)
C0686721|Shaken baby syndrome - non-accidental injury
C0686721|Shaken baby
C0270611|Brain Injuries
C0270611|Brain Injury
C0270611|Injury, Brain
C0270611|Damage, brain
C0270611|Brain Damage
C0270611|BRAIN INJ
C0270611|INJ BRAIN
C0270611|brain lesion (from injury)
C0270611|brain injury (diagnosis)
C0270611|Brain injury NOS
C0270611|Brain Injuries [Disease/Finding]
C0270611|Injuries, Brain
C0270611|Injury;cerebral
C0270611|Acquired brain injury
C0270611|Intracerebral injury
C0270611|Intracerebral injury NOS
C0270611|Brain injury NOS (disorder)
C0270611|Cerebral damage
C0270611|Acquired brain injury (disorder)
C0270611|Brain damage (disorder)
C0270611|Brain tissue injury
C0270611|brain; damage
C0270611|brain; injury
C0270611|cerebral; injury
C0270611|damage; brain
C0270611|injury; brain
C0270611|injury; cerebral
C0270611|Brain damage, NOS
C0270611|Injury;brain;acquired
C0270611|cerebral injury
C0876926|ENCEPH TRAUMATIC
C0876926|TRAUMATIC BRAIN INJ
C0876926|INJ BRAIN TRAUMATIC
C0876926|BRAIN INJ TRAUMATIC
C0876926|TRAUMATIC ENCEPH
C0876926|traumatic brain injury
C0876926|traumatic brain injury (diagnosis)
C0876926|brain injury due to trauma
C0876926|brain trauma
C0876926|Brain damage (traumatic)
C0876926|TBI
C0876926|Brain damage - traumatic
C0876926|Traumatic encephalopathy
C0876926|Traumatic encephalopathy (disorder)
C0876926|traumatic brain damage (diagnosis)
C0876926|traumatic brain damage
C0876926|brain damage traumatic
C0876926|Encephalopathy, Traumatic
C0876926|TBI (Traumatic Brain Injury)
C0876926|Trauma, Brain
C0876926|Injury, Brain, Traumatic
C0876926|Brain damage - traumatic (disorder)
C0876926|Traumatic brain injury (disorder)
C0876926|encephalopathy; traumatic
C0876926|traumatic; encephalopathy
C0876926|Traumatic encephalopathy (disorder) [Ambiguous]
C0876926|Brain Injury (Traumatic)
C0876926|Brain Injuries, Traumatic
C0876926|Brain Injury, Traumatic
C0876926|Injuries, Traumatic Brain
C0876926|Injury, Traumatic Brain
C0876926|Traumatic Brain Injuries
C0876926|Brain Traumas
C0876926|Traumas, Brain
C0876926|Encephalopathies, Traumatic
C0876926|Traumatic Encephalopathies
C0876926|TBIs (Traumatic Brain Injury)
C0876926|Injury;brain;traumatic
C1403070|brain injury cicatrix
C1403070|brain cicatrix
C1403070|cicatrix due to brain injury (diagnosis)
C1403070|cicatrix due to brain injury
C1403070|brain; cicatrix
C1403070|brain; scar
C1403070|scar; brain
C1399577|acquired brain deformity due to injury (diagnosis)
C1399577|brain injury acquired deformity
C1399577|acquired brain deformity due to injury
C1399577|acquired brain deformity
C1399577|brain; deformity, acquired
C1399577|deformity; brain, acquired
C2729127|cerebral granuloma due to injury
C2729127|cerebral granuloma due to injury (diagnosis)
C2729127|brain injury cerebral granuloma
C2729128|brain hypertrophy due to injury (diagnosis)
C2729128|brain hypertrophy due to injury
C2729128|brain injury hypertrophy
C2729129|brain induration due to injury (diagnosis)
C2729129|brain injury induration
C2729129|brain induration due to injury
C2729130|intracranial pneumatocele due to injury (diagnosis)
C2729130|intracranial pneumatocele due to injury
C2729130|brain injury intracranial pneumatocele
C2728325|medullary depression due to brain injury (diagnosis)
C2728325|medullary depression due to brain injury
C2728325|brain injury medullary depression
C2728507|Morel-Lavallee lesion due to brain injury
C2728507|Morel-Lavallee lesion due to brain injury (diagnosis)
C2728507|brain injury Morel-Lavallee lesion
C2729131|pneumocephalus due to brain injury (diagnosis)
C2729131|brain injury pneumocephalus
C2729131|pneumocephalus due to brain injury
C2728280|brain injury respiratory center depression
C2728280|respiratory center depression due to brain injury
C2728280|respiratory center depression due to brain injury (diagnosis)
C2728512|speech impediment due to brain injury
C2728512|brain injury speech impediment due to organic lesion
C2728512|speech impediment due to organic lesion
C2728512|speech impediment due to brain injury (diagnosis)
C0433845|Cortex laceration with open intracranial wound and prolonged loss of consciousness (more than 24 hours) without return to pre-existing conscious level
C0433845|Cortex (cerebral) lacer with open intcran wound, with prolonged loc, w/o rtrn to pecl
C0433845|Opn cortex lac-deep coma
C0433845|Cortex (cerebral) laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0433845|Cortex laceration with open intracranial wound AND prolonged loss of consciousness (more than 24 hours) without return to pre-existing conscious level (disorder)
C0433845|Cortex laceration with open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious level
C0433845|Cortex laceration with open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious level (disorder)
C0433845|Cerebral cortex laceration with open intracranial wound, with more than 24 hours loss of consciousness, without return to pre-existing conscious level
C0433845|Cortex laceration with open intracranial wound, with more than 24 hours loss of consciousness, without return to pre-existing conscious level
C0433845|Cerebral cortex laceration with open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C0433845|Cortex laceration with open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C3509561|birth trauma brain damage
C3509561|brain damage due to birth trauma
C3509561|brain damage due to birth trauma (diagnosis)
C0149844|Brain Contusions
C0149844|Contusion, Brain
C0149844|Contusions, Brain
C0149844|Brain contusion
C0149844|Contusion of brain
C0149844|Contusion of brain (diagnosis)
C0149844|head injury contusion of brain
C0149844|Contusional brain injury
C0149844|Contusion of brain (disorder)
C0149844|brain; contusion
C0149844|contusion; brain
C0149844|Contusion of brain, NOS
C0750973|ENCEPH POST TRAUMATIC
C0750973|POST TRAUMATIC ENCEPH
C0750973|Encephalopathies, Post-Traumatic
C0750973|Encephalopathy, Post Traumatic
C0750973|Post Traumatic Encephalopathy
C0750973|Post-Traumatic Encephalopathies
C0750973|Post-traumatic encephalopathy
C0750973|Encephalopathy, Post-Traumatic
C0750971|cerebral contusion
C0750971|cerebral contusion (diagnosis)
C0750971|Contusion, Cortical
C0750971|Contusions, Cortical
C0750971|Cortical Contusions
C0750971|Contusion;cerebral
C0750971|Cortical Contusion
C0750971|Contusion of cerebrum
C0750971|Contusion of cerebrum (disorder)
C0750971|cerebral; contusion
C0750971|contusion; cerebral
C0750971|Cerebral contusion, NOS
C0750972|POST CONCUSSIVE ENCEPH
C0750972|ENCEPH POST CONCUSSIVE
C0750972|Encephalopathies, Post-Concussive
C0750972|Encephalopathy, Post Concussive
C0750972|Post Concussive Encephalopathy
C0750972|Post-Concussive Encephalopathies
C0750972|Post-Concussive Encephalopathy
C0750972|Encephalopathy, Post-Concussive
C0452047|Focal brain injury
C0452047|FOCAL BRAIN INJ
C0452047|BRAIN INJ FOCAL
C0452047|Brain Injury, Focal
C0452047|Injuries, Focal Brain
C0452047|Injury, Focal Brain
C0452047|Brain Injuries, Focal
C0452047|Focal Brain Injuries
C0452047|Focal brain injury (disorder)
C0452047|brain; injury, focal
C0452047|injury; brain, focal
C0085742|Acute Brain Injury
C0085742|Brain Injury, Acute
C0085742|Injury, Acute Brain
C0085742|INJ ACUTE BRAIN
C0085742|ACUTE BRAIN INJ
C0085742|BRAIN INJ ACUTE
C0085742|Injuries, Acute Brain
C0085742|Acute Brain Injuries
C0085742|Brain Injuries, Acute
C0272945|Brain Laceration
C0272945|Laceration, Brain
C0272945|Lacerations, Brain
C0272945|Laceration of brain (disorder)
C0272945|Lacerating brain injury
C0272945|Laceration of brain
C0272945|Laceration of brain (diagnosis)
C0272945|brain; laceration
C0272945|laceration; brain
C0272945|Laceration of brain, NOS
C0272945|Brain Lacerations
C0433856|Diffuse brain injury
C0433856|BRAIN INJ DIFFUSE
C0433856|Brain Injury, Diffuse
C0433856|Diffuse Brain Injuries
C0433856|Injuries, Diffuse Brain
C0433856|Injury, Diffuse Brain
C0433856|Diffuse axonal brain injury
C0433856|Diffuse brain injury (disorder)
C0433856|Brain Injuries, Diffuse
C0433856|brain; injury, diffuse
C0433856|injury; brain, diffuse
C0003132|Anoxic Encephalopathy
C0003132|ANOXIC ENCEPH
C0003132|Brain Damage, Anoxic
C0003132|Damage, Anoxic Brain
C0003132|Anoxic Encephalopathies
C0003132|Encephalopathies, Anoxic
C0003132|Encephalopathy, Anoxic
C0003132|Anoxic brain damage
C0003132|Anoxic encephalopathy (disorder)
C0003132|Anoxic brain injury
C0003132|Anoxic brain damage, NOS
C0003132|Anoxic encephalopathy, NOS
C0003132|Anoxic encephalopathy [dup] (disorder)
C0242670|Persistent Vegetative State
C0242670|Persistent Vegetative States
C0242670|Vegetative States, Persistent
C0242670|persistent vegetative state (diagnosis)
C0242670|Persistent Unawareness States
C0242670|State, Persistent Unawareness
C0242670|States, Persistent Unawareness
C0242670|Unawareness State, Persistent
C0242670|Unawareness States, Persistent
C0242670|State, Persistent Vegetative
C0242670|States, Persistent Vegetative
C0242670|Persistent vegtv state
C0242670|Persistent Unawareness State
C0242670|Persistent Vegetative State [Disease/Finding]
C0242670|PVS (Persistent Vegetative State)
C0242670|Vegetative State, Persistent
C0242670|PVSs (Persistent Vegetative State)
C0242670|Persistent vegetative state (disorder)
C0242670|Chronic vegetative state
C0242670|Vegetative state chronic
C0242670|PVS - Persistent vegetative state
C0549117|Frontal lobe syndrome
C0549117|frontal lobe syndrome (diagnosis)
C0549117|Frontal lobe syndrome (disorder)
C0549117|[X]Frontal lobe syndrome
C0549117|frontal lobe; syndrome
C0549117|syndrome; frontal lobe
C0006110|Brain Death
C0006110|cerebral death
C0006110|Death, Brain
C0006110|brain death (diagnosis)
C0006110|Brain Deads
C0006110|Brain Death [Disease/Finding]
C0006110|Coma Depasse
C0006110|Brain Dead
C3508472|brain injury traumatic mild (diagnosis)
C3508472|brain injury traumatic mild
C3508472|Mild Traumatic Brain Injury
C3508472|Injury, Brain, Traumatic Mild
C0272927|Closed traumatic brain injury
C0272927|Brain injury without open intracranial wound
C0272927|brain injury without open intracranial wound (diagnosis)
C0272927|Brain injury without open intracranial wound (disorder)
C0272927|Brain injury without open intracranial wound, NOS
C0021879|Brain injury NEC
C0021879|Intcran inj of oth and unspec nature, w/o ment of open intcran wound, with state of cons unspec
C0021879|Intracranial injury of other and unspecified nature without mention of open intracranial wound, unspecified state of consciousness
C1140716|HYPOXIC ENCEPH
C1140716|ENCEPH HYPOXIC
C1140716|Brain disorder resulting from a period of impaired oxygen delivery to the brain
C1140716|Brain Damage, Hypoxic
C1140716|Damage, Hypoxic Brain
C1140716|Encephalopathies, Hypoxic
C1140716|Hypoxic Encephalopathies
C1140716|Hypoxic brain damage
C1140716|Brain damage due to hypoxia
C1140716|Hypoxic brain injury
C1140716|Hypoxic-ischemic brain injury
C1140716|Hypoxic-ischaemic brain injury
C1140716|Hypoxic encephalopathy
C1140716|Encephalopathy, Hypoxic
C1140716|Brain disorder resulting from a period of impaired oxygen delivery to the brain (disorder)
C0338418|Acute Necrotizing Encephalitides
C0338418|Acute Necrotizing Encephalitis
C0338418|Encephalitides, Acute Necrotizing
C0338418|Necrotizing Encephalitides, Acute
C0338418|Necrotizing Encephalitis, Acute
C0338418|ENCEPH ACUTE NECROTIZING
C0338418|viral encephalitis acute necrotizing
C0338418|Acute necrotizing encephalitis (diagnosis)
C0338418|Acute necrotising encephalitis
C0338418|Acute necrotizing viral encephalitis
C0338418|Acute necrotising viral encephalitis
C0338418|Acute necrotizing encephalitis (disorder)
C0338418|Encephalitis, Acute Necrotizing
C3897170|White Matter Injury
C1456496|Brain damage
C1456496|Traumatic AND/OR non-traumatic brain injury
C1456496|Traumatic AND/OR non-traumatic brain injury (disorder)
C0149843|Punch drunk
C0149843|Punch drunk syndrome
C0149843|Punch drunk syndrome (diagnosis)
C0149843|head injury with dementia punch drunk syndrome
C0149843|Boxer's dementia
C0149843|Dementia pugilistica
C0149843|Punchdrunk encephalopathy
C0149843|Punch drunk syndrome (disorder)
C0160293|Brain injury NEC-no coma
C0160293|Intcran inj of oth and unspec nature, w/o ment of open intcran wound, with no loc
C0160293|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with no loss of consciousness
C0160294|Brain inj NEC-brief coma
C0160294|Intcran inj of oth and unspec nature, w/o ment of open intcran wound, with brief loc
C0160294|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160298|Brain inj NEC-coma NOS
C0160298|Intcran inj of oth and unspec nature, w/o ment of open intcran wound, with loc of unspec dura
C0160298|Intracranial injury of other and unspecified nature without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0006109|Chronic brain syndrome
C0006109|Brain Damage, Chronic
C0006109|Chronic Brain Damage
C0006109|ENCEPH CHRONIC
C0006109|CHRONIC ENCEPH
C0006109|Brain syndrome chronic
C0006109|Syndrome brain chronic
C0006109|Encephalopathy, Chronic
C0006109|Brain Damage, Chronic [Disease/Finding]
C0006109|Chronic Encephalopathy
C0006109|Encephalopathy chronic
C0006109|Chronic brain syndrome (disorder)
C0006109|Chronic brain syndrome, NOS
C0006109|Chronic encephalopathy, NOS
C0160292|Intracranial injury of other and unspecified nature
C0021878|Intracranial injury of other and unspecified nature without mention of open intracranial wound
C1321905|Dysfunction, Minimal Brain
C1321905|minimal brain dysfunction
C1321905|Minimal brain dysfunction (disorder)
C1321905|MBD - Minimal brain dysfunction
C1321905|Minimal Brain Disorders
C1321905|Brain Dysfunction, Minimal
C0695222|Cerebellar or brain stem contusion with open intracranial wound, with concussion, unspecified
C0695222|Opn cerebel cont-concuss
C0695224|Cerebellar or brain stem laceration with open intracranial wound, with concussion, unspecified
C0695224|Opn cerebell lac-concuss
C0433815|Cortex (cerebral) contu w/o ment of open intcran wound, state of consciousness unspec
C0433815|Cerebral cortx contusion
C0433815|Cortex (cerebral) contusion without mention of open intracranial wound, unspecified state of consciousness
C0433815|Cortex contusion without mention of open intracranial wound, with unspecified state of consciousness (disorder)
C0433815|Cortex contusion without mention of open intracranial wound, with unspecified state of consciousness
C0433815|Cerebral cortex contusion without mention of open intracranial wound, state of consciousness unspecified
C0433815|Cortex contusion without mention of open intracranial wound, state of consciousness unspecified
C0433821|Cortex (cerebral) contu w/o ment of open intcran wound, with loc of unspec duration
C0433821|Cortex contus-coma NOS
C0433821|Cortex contusion without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433821|Cortex contusion without mention of open intracranial wound, with loss of consciousness of unspecified duration (disorder)
C0433821|Cortex (cerebral) contusion without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433821|Cerebral cortex contusion without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433846|Cortex (cerebral) laceration without mention of open intracranial wound
C0433846|Cortex laceration without mention of open intracranial wound (disorder)
C0433846|Cortex laceration without mention of open intracranial wound
C0433846|Cerebral cortex laceration without mention of open intracranial wound
C0433847|Cortex (cerebral) lacer w/o ment of open intcran wound, with state of consciousness unspec
C0433847|Cerebral cortex lacerat
C0433847|Cortex (cerebral) laceration without mention of open intracranial wound, unspecified state of consciousness
C0433847|Cortex laceration without mention of open intracranial wound, unspecified state of consciousness (disorder)
C0433847|Cortex laceration without mention of open intracranial wound, unspecified state of consciousness
C0433847|Cerebral cortex laceration without mention of open intracranial wound, with state of consciousness unspecified
C0433847|Cortex laceration without mention of open intracranial wound, with state of consciousness unspecified
C0433848|Cortex (cerebral) lacer w/o ment of open intcran wound, with no loc
C0433848|Cortex lacerat w/o coma
C0433848|Cortex laceration without mention of open intracranial wound, with no loss of consciousness
C0433848|Cortex laceration without mention of open intracranial wound, with no loss of consciousness (disorder)
C0433848|Cortex (cerebral) laceration without mention of open intracranial wound, with no loss of consciousness
C0433848|Cerebral cortex laceration without mention of open intracranial wound, with no loss of consciousness
C0433853|Cortex (cerebral) lacer w/o ment of open intcran wound, with loc of unspec duration
C0433853|Cortex lacerat-coma NOS
C0433853|Cortex laceration without mention of open intracranial wound, with loss of consciousness of unspecified duration (disorder)
C0433853|Cortex laceration without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433853|Cortex (cerebral) laceration without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433853|Cerebral cortex laceration without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433854|Cortex (cerebral) lacer w/o ment of open intcran wound, with concussion, unspec
C0433854|Cortex lacerat-concuss
C0433854|Cortex laceration without mention of open intracranial wound, with concussion, unspecified (disorder)
C0433854|Cortex laceration without mention of open intracranial wound, with concussion, unspecified
C0433854|Cortex (cerebral) laceration without mention of open intracranial wound, with concussion, unspecified
C0433854|Cerebral cortex laceration without mention of open intracranial wound, with concussion, unspecified
C0859613|Cortex (cerebral) contu w/o ment of open intcran wound, with no loc
C0160131|Cortex (cerebral) contu w/o ment of open intcran wound, with brief loc
C0160131|Cortex contus-brief coma
C0160131|Cortex (cerebral) contusion without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160131|Cerebral cortex contusion without mention of open intracranial wound, with brief loss of consciousness
C0160131|Cortex contusion without mention of open intracranial wound, with brief loss of consciousness
C0272955|Cortex contusion without open intracranial wound AND with moderate loss of consciousness (1-24 hours) (disorder)
C0272955|Cortex contusion without open intracranial wound and with moderate loss of consciousness (1-24 hours)
C0272955|Cortex (cerebral) contu w/o ment of open intcran wound, with moderate loc
C0272955|Cortex contus-mod coma
C0272955|Cortex contusion without mention of intracranial wound, with 1-24 hours loss of consciousness (disorder)
C0272955|Cortex contusion without mention of intracranial wound, with 1-24 hours loss of consciousness
C0272955|contusion of cortex w/o open intracranial wound, with moderate loc (1-24 hours)
C0272955|cortex contusion without open intracranial wound, with moderate loss of consciousness (1-24 hours)
C0272955|cortex contusion without open intracranial wound, with moderate loss of consciousness (1-24 hours) (diagnosis)
C0272955|Cortex (cerebral) contusion without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0272955|Cerebral cortex contusion without mention of open intracranial wound, with 1-24 hours loss of consciousness
C0272955|Cortex contusion without mention of open intracranial wound, with 1-24 hours loss of consciousness
C0272955|Cerebral cortex contusion without mention of open intracranial wound, with moderate loss of consciousness
C0272955|Cortex contusion without mention of open intracranial wound, with moderate loss of consciousness
C0160133|Cortex (cerebral) contu w/o ment of open intcran wound, with prolonged loc and rtrn to pecl
C0160133|Cortx contus-prolng coma
C0160133|Cortex (cerebral) contusion without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160133|Cerebral cortex contusion without mention of open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0160133|Cortex contusion without mention of open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0160134|Cortex (cerebral) contu w/o ment of open intcran wound, with prolonged loc, w/o rtrn to pecl
C0160134|Cortex contus-deep coma
C0160134|Cortex (cerebral) contusion without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160134|Cerebral cortex contusion without mention of open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C0160134|Cortex contusion without mention of open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C0695217|Cortex (cerebral) contu w/o ment of open intcran wound, with concussion, unspec
C0695217|Cortex contus-concus NOS
C0695217|Cortex (cerebral) contusion without mention of open intracranial wound, with concussion, unspecified
C0695217|Cerebral cortex contusion without mention of open intracranial wound, with concussion, unspecified
C0695217|Cortex contusion without mention of open intracranial wound, with concussion, unspecified
C0160138|Cortex (cerebral) contu with open intcran wound, w/o ment of specific state of consciousness
C0160138|Cortex (cerebral) contusion with open intracranial wound, with state of consciousness unspecified
C0160138|Cortex contusion/opn wnd
C0160138|Cortex (cerebral) contusion with open intracranial wound, without mention of specific state of consciousness
C0160138|Cortex (cerebral) contusion with open intracranial wound, unspecified state of consciousness
C0160138|Cerebral cortex contusion with open intracranial wound, without mention of specific state of consciousness
C0160138|Cortex contusion with open intracranial wound, without mention of specific state of consciousness
C0160140|Cortex (cerebral) contu with open intcran wound, with brief loc
C0160140|Opn cort contus-brf coma
C0160140|Cortex (cerebral) contusion with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160140|Cerebral cortex contusion with open intracranial wound, with brief loss of consciousness
C0160140|Cortex contusion with open intracranial wound, with brief loss of consciousness
C0160141|Cortex (cerebral) contu with open intcran wound, with moderate loc
C0160141|Opn cort contus-mod coma
C0160141|Cortex (cerebral) contusion with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160141|Cerebral cortex contusion with open intracranial wound, with moderate loss of consciousness
C0160141|Cortex contusion with open intracranial wound, with moderate loss of consciousness
C0160142|Cortex (cerebral) contu with open intcran wound, with prolonged loc and rtrn to pecl
C0160142|Opn cort contu-prol coma
C0160142|Cortex (cerebral) contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160142|Cerebral cortex contusion with open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0160142|Cortex contusion with open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0160143|Cortex (cerebral) contu with open intcran wound, with prolonged loc, w/o rtrn to pecl
C0160143|Opn cort contu-deep coma
C0160143|Cortex (cerebral) contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160143|Cerebral cortex contusion with open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C0160143|Cortex contusion with open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C0859614|Cortex (cerebral) contu with open intcran wound, with loc of unspec duration
C0160149|Cortex (cerebral) lacer w/o ment of open intcran wound, with brief loc
C0160149|Cortex lacera-brief coma
C0160149|Cortex (cerebral) laceration without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160149|Cerebral cortex laceration without mention of open intracranial wound, with brief loss of consciousness
C0160149|Cortex laceration without mention of open intracranial wound, with brief loss of consciousness
C0160150|Cortex (cerebral) lacer w/o ment of open intcran wound, with moderate loc
C0160150|Cortex lacerat-mod coma
C0160150|Cortex (cerebral) laceration without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160150|Cerebral cortex laceration without mention of open intracranial wound, with moderate loss of consciousness
C0160150|Cortex laceration without mention of open intracranial wound, with moderate loss of consciousness
C0160151|Cortex (cerebral) lacer w/o ment of open intcran wound, with prolonged loc and rtrn to pecl
C0160151|Cortex lacerat-prol coma
C0160151|Cortex (cerebral) laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160151|Cerebral cortex laceration without mention of open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0160151|Cortex laceration without mention of open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0160152|Cortex (cerebral) lacer w/o ment of open intcran wound, with prolonged loc, w/o rtrn to pecl
C0160152|Cortex lacerat-deep coma
C0160152|Cortex (cerebral) laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160152|Cerebral cortex laceration without mention of open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C0160152|Cortex laceration without mention of open intracranial wound, with prolonged loss of consciousness, without return to pre-existing conscious level
C0160158|Cortex (cerebral) lacer with open intcran wound, with brief loc
C0160158|Opn cortx lac-brief coma
C0160158|Cortex (cerebral) laceration with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160158|Cerebral cortex laceration with open intracranial wound, with brief loss of consciousness
C0160158|Cortex laceration with open intracranial wound, with brief loss of consciousness
C0160159|Cortex (cerebral) lacer with open intcran wound, with moderate loc
C0160159|Opn cortx lacer-mod coma
C0160159|Cortex (cerebral) laceration with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160159|Cerebral cortex laceration with open intracranial wound, with moderate loss of consciousness
C0160159|Cortex laceration with open intracranial wound, with moderate loss of consciousness
C0160160|Cortex (cerebral) lacer with open intcran wound, with prolonged loc and rtrn to pecl
C0160160|Opn cortx lac-proln coma
C0160160|Cortex (cerebral) laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160160|Cerebral cortex laceration with open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0160160|Cortex laceration with open intracranial wound, with prolonged loss of consciousness and return to pre-existing conscious level
C0859615|Cortex (cerebral) lacer with open intcran wound, with loc of unspec duration
C0160165|Cerebellar or brain stem contu w/o ment of open intcran wound, with state of cons unspec
C0160165|Cerebel/brain stm contus
C0160165|Cerebellar or brain stem contusion without mention of open intracranial wound, unspecified state of consciousness
C0160166|Cerebellar or brain stem contu w/o ment of open intcran wound, with no loc
C0160166|Cerebell contus w/o coma
C0160166|Cerebellar or brain stem contusion without mention of open intracranial wound, with no loss of consciousness
C0160167|Cerebellar or brain stem contu w/o ment of open intcran wound, with brief loc
C0160167|Cerebell contus-brf coma
C0160167|Cerebellar or brain stem contusion without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160168|Cerebellar or brain stem contu w/o ment of open intcran wound, with moderate loc
C0160168|Cerebell contus-mod coma
C0160168|Cerebellar or brain stem contusion without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160170|Cerebellar or brain stem contu w/o ment of open intcran wound, with prolonged loc, w/o rtrn to pecl
C0160170|Cerebel contus-deep coma
C0160170|Cerebellar or brain stem contusion without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160171|Cerebellar or brain stem contu w/o ment of open intcran wound, with loc of unspec duration
C0160171|Cerebell contus-coma NOS
C0160171|Cerebellar or brain stem contusion without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0695221|Cerebellar or brain stem contu w/o ment of open intcran wound, with concussion, unspec
C0695221|Cerebell contus-concuss
C0695221|Cerebellar or brain stem contusion without mention of open intracranial wound, with concussion, unspecified
C0160174|Cerebellar or brain stem contu with open intcran wound, with state of consciousness unspec
C0160174|Cerebel contus w opn wnd
C0160174|Cerebellar or brain stem contusion with open intracranial wound, unspecified state of consciousness
C0160176|Cerebellar or brain stem contu with open intcran wound, with brief loc
C0160176|Opn cerebe cont-brf coma
C0160176|Cerebellar or brain stem contusion with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160177|Cerebellar or brain stem contusion with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160177|Cerebellar or brain stem contu with open intcran wound, with moderate loc
C0160177|Opn cerebe cont-mod coma
C0160178|Cerebellar or brain stem contu with open intcran wound, with prolonged loc and return to pecl
C0160178|Opn cerebe cont-prol com
C0160178|Cerebellar or brain stem contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160179|Cerebellar or brain stem contu with open intcran wound, with prolonged loc, w/o return to pecl
C0160179|Opn cerebe cont-deep com
C0160179|Cerebellar or brain stem contusion with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160180|Cerebellar or brain stem contu with open intcran wound, with loc of unspec duration
C0160180|Opn cerebe cont-coma NOS
C0160180|Cerebellar or brain stem contusion with open intracranial wound, with loss of consciousness of unspecified duration
C0160183|Cerebellar or brain stem lacer w/o ment of open intcran wound, with state of consciousness unspec
C0160183|Cerebel/brain stem lacer
C0160183|Cerebellar or brain stem laceration without mention of open intracranial wound, unspecified state of consciousness
C0160184|Cerebellar or brain stem lacer w/o ment of open intcran wound, with no loc
C0160184|Cerebel lacerat w/o coma
C0160184|Cerebellar or brain stem laceration without mention of open intracranial wound, with no loss of consciousness
C0160185|Cerebellar or brain stem lacer w/o ment of open intcran wound, with brief loc
C0160185|Cerebel lacer-brief coma
C0160185|Cerebellar or brain stem laceration without mention of open intracranial wound, with brief [less than 1 hour] loss of consciousness
C0160186|Cerebellar or brain stem lacer w/o ment of open intcran wound, with moderate loc
C0160186|Cerebel lacerat-mod coma
C0160186|Cerebellar or brain stem laceration without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160187|Cerebellar or brain stem lacer w/o ment of open intcran wound, with prolonged loc and rtrn to pecl
C0160187|Cerebel lacer-proln coma
C0160187|Cerebellar or brain stem laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160188|Cerebellar or brain stem lacer w/o ment of open intcran wound, with prolonged loc, w/o rtrn to pecl
C0160188|Cerebell lacer-deep coma
C0160188|Cerebellar or brain stem laceration without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160189|Cerebellar or brain stem lacer w/o ment of open intcran wound, with loc of unspec duration
C0160189|Cerebel lacerat-coma NOS
C0160189|Cerebellar or brain stem laceration without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0695223|Cerebellar or brain stem lacer w/o ment of open intcran wound, with concussion, unspec
C0695223|Cerebel lacer-concussion
C0695223|Cerebellar or brain stem laceration without mention of open intracranial wound, with concussion, unspecified
C0160192|Cerebellar or brain stem lacer with open intcran wound, with state of consciousness unspec
C0160192|Cerebel lacer w open wnd
C0160192|Cerebellar or brain stem laceration with open intracranial wound, unspecified state of consciousness
C0160194|Cerebellar or brain stem lacer with open intcran wound, with brief loc
C0160194|Opn cerebel lac-brf coma
C0160194|Cerebellar or brain stem laceration with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160195|Cerebellar or brain stem lacer with open intcran wound, with moderate loc
C0160195|Opn cerebel lac-mod coma
C0160195|Cerebellar or brain stem laceration with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160196|Cerebellar or brain stem lacer with open intcran wound, with prolonged loc and return to pecl
C0160196|Opn cerebe lac-prol coma
C0160196|Cerebellar or brain stem laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160197|Cerebellar or brain stem lacer with open intcran wound, with prolonged loc, w/o return to pecl
C0160197|Opn cerebe lac-deep coma
C0160197|Cerebellar or brain stem laceration with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160198|Cerebellar or brain stem lacer with open intcran wound, with loc of unspec duration
C0160198|Opn cerebel lac-coma NOS
C0160198|Cerebellar or brain stem laceration with open intracranial wound, with loss of consciousness of unspecified duration
C0160201|Oth and unspec cerebral lacer and contu, w/o ment of open intcran wound, with state of cons unspec
C0160201|Brain laceration NEC
C0160201|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, unspecified state of consciousness
C0160202|Oth and unspec cerebral lacer and contu, w/o ment of open intcran wound, with no loc
C0160202|Brain lacer NEC w/o coma
C0160202|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with no loss of consciousness
C0160203|Oth and unspec cerebral lacer and contu, w/o ment of open intcran wound, with brief loc
C0160203|Brain lac NEC-brief coma
C0160203|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with brief [less than one hour] loss of consciousness
C0160204|Oth and unspec cerebral lacer and contu, w/o ment of open intcran wound, with moderate loc
C0160204|Brain lacer NEC-mod coma
C0160204|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160205|Oth and unspec cereb lacer and contu, w/o ment of open intcran wound, prol loc and rtrn to pecl
C0160205|Brain lac NEC-proln coma
C0160205|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre- existing conscious level
C0160206|Oth and unspec cereb lacer and contu, w/o ment of open intcran wound, prol loc, w/o rtrn to pecl
C0160206|Brain lac NEC-deep coma
C0160206|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160207|Oth and unspec cereb lacer and contu, w/o ment of open intcran wound, with loc of unspec duration
C0160207|Brain lacer NEC-coma NOS
C0160207|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0695225|Oth and unspec cerebral lacer and contu, w/o ment of open intcran wound, with concus, unspec
C0695225|Brain lacer NEC-concuss
C0695225|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound, with concussion, unspecified
C0160210|Oth and unspec cerebral lacer and contu, with open intcran wound, with state of cons unspec
C0160210|Brain lac NEC w open wnd
C0160210|Other and unspecified cerebral laceration and contusion, with open intracranial wound, unspecified state of consciousness
C0160211|Oth and unspec cerebral lacer and contu, with open intcran wound, with no loc
C0160211|Opn brain lacer w/o coma
C0160211|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with no loss of consciousness
C0160212|Oth and unspec cerebral lacer and contu, with open intcran wound, with brief loc
C0160212|Opn brain lac-brief coma
C0160212|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with brief [less than one hour] loss of consciousness
C0160213|Oth and unspec cerebral lacer and contu, with open intcran wound, with moderate loc
C0160213|Opn brain lacer-mod coma
C0160213|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with moderate [1-24 hours] loss of consciousness
C0160214|Oth and unspec cereb lacer and contu, with open intcran wound, with prol loc and rtrn to pecl
C0160214|Opn brain lac-proln coma
C0160214|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness and return to pre-existing conscious level
C0160215|Oth and unspec cereb lacer and contu, with open intcran wound, with prol loc, w/o rtrn to pecl
C0160215|Open brain lac-deep coma
C0160215|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0160216|Oth and unspec cerebral lacer and contu, with open intcran wound, with loc of unspec duration
C0160216|Opn brain lacer-coma NOS
C0160216|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with loss of consciousness of unspecified duration
C0695226|Oth and unspec cerebral lacer and contu, with open intcran wound, with concussion, unspec
C0695226|Open brain lacer-concuss
C0695226|Other and unspecified cerebral laceration and contusion, with open intracranial wound, with concussion, unspecified
C0859744|Cerebral laceration and contusion, without mention of open intracranial wound
C0859745|Cerebral laceration & contusion with open intracranial wound
C0859782|Cerebellar or brain stem contu w/o ment of open intcran wound, with prol loss cons and rtrn to pecl
C0859782|Cerebellar or brain stem contu w/o ment of open intcran wound, with prol loc and return to pecl
C0160128|Cortex (cerebral) contusion without mention of open intracranial wound
C0160128|Cerebral cortex contusion without mention of open intracranial wound
C0160128|Cortex contusion without mention of open intracranial wound
C0160164|Cerebellar or brain stem contusion without mention of open intracranial wound
C0160173|Cerebellar or brain stem contusion with open intracranial wound
C0160182|Cerebellar or brain stem laceration without mention of open intracranial wound
C0160191|Cerebellar or brain stem laceration with open intracranial wound
C0160200|Other and unspecified cerebral laceration and contusion, without mention of open intracranial wound
C0160209|Other and unspecified cerebral laceration and contusion, with open intracranial wound
C0160137|Cortex (cerebral) contusion with open intracranial wound
C0160137|Cortex contusion with open intracranial wound
C0160137|Cortex contusion with open intracranial wound (diagnosis)
C0160137|contusion of cortex with open intracranial wound
C0160137|Contusion of cerebral cortex with open intracranial wound
C0160137|Cortex contusion with open intracranial wound (disorder)
C0160137|Cerebral cortex contusion with open intracranial wound
C0160127|Cerebral laceration and contusion
C0160127|cerebral laceration and contusion (diagnosis)
C0160127|Cerebral laceration and contusion NOS
C0160127|Cerebral laceration and contusion (disorder)
C0160127|Cerebral laceration and contusion NOS (disorder)
C0160127|Brain laceration and contusion NOS
C0274278|Late effect of intracranial injury without mention of skull fracture
C0274278|Sequelae of intracranial injury
C0274278|Lt eff intracranial inj
C0274278|late effect of intracranial injury without skull fracture (diagnosis)
C0274278|Late effect of intracranial injury without skull fracture
C0274278|Late effect of intracranial injury without skull fracture (disorder)
C0272961|Cortex (cerebral) contusion with open intracranial wound, with no loss of consciousness
C0272961|Cortex contusion with open intracranial wound and no loss of consciousness
C0272961|cerebral contusion with open intracranial wound with no loss of consciousness (diagnosis)
C0272961|cerebral contusion with open intracranial wound with no loss of consciousness
C0272961|Opn cortx contus-no coma
C0272961|Cortex contusion with open intracranial wound AND no loss of consciousness (disorder)
C0272961|Cortex contusion with open intracranial wound, with no loss of consciousness
C0272961|Cortex contusion with open intracranial wound, with no loss of consciousness (disorder)
C0272961|Cerebral cortex contusion with open intracranial wound, with no loss of consciousness
C0160175|Cerebellar or brain stem contusion with open intracranial wound, with no loss of consciousness
C0160175|Opn cerebe cont w/o coma
C0160193|Cerebellar or brain stem laceration with open intracranial wound, with no loss of consciousness
C0160193|Opn cerebel lac w/o coma
C0272967|cerebral contusion with open intracranial wound with concussion (diagnosis)
C0272967|cerebral contusion w/ open intracranial wound w/ concussion
C0272967|cerebral contusion with open intracranial wound with concussion
C0272967|Cortex (cerebral) contusion with open intracranial wound, with concussion, unspecified
C0272967|Opn cortx contus-concuss
C0272967|Cortex contusion with open intracranial wound, with concussion, unspecified (disorder)
C0272967|Cortex contusion with open intracranial wound, with concussion, unspecified
C0272967|Cortex contusion with open intracranial wound AND concussion (disorder)
C0272967|Cortex contusion with open intracranial wound AND concussion
C0272967|Cortex contusion with open intracranial wound and unspecified concussion
C0272967|Cerebral cortex contusion with open intracranial wound, with concussion, unspecified
C0272977|Cortex (cerebral) laceration with open intracranial wound
C0272977|laceration of cerebrum with open intracranial wound
C0272977|laceration of cerebrum with open intracranial wound (diagnosis)
C0272977|Cortex laceration with open intracranial wound (finding)
C0272977|Cortex laceration with open intracranial wound
C0272977|Cortex laceration with open intracranial wound (disorder)
C0272977|Cerebral cortex laceration with open intracranial wound
C0272978|Cortex (cerebral) laceration with open intracranial wound, with state of consciousness unspecified
C0272978|Cortex laceration with open intracranial wound and unspecified state of consciousness -RETIRED-
C0272978|Cortex lacer w opn wound
C0272978|Cortex (cerebral) laceration with open intracranial wound, unspecified state of consciousness
C0272978|Cortex laceration with open intracranial wound and unspecified state of consciousness
C0272978|Cortex laceration with open intracranial wound and unspecified state of consciousness (disorder)
C0272978|Cortex laceration with open intracranial wound, unspecified state of consciousness
C0272978|Cortex laceration with open intracranial wound, unspecified state of consciousness (disorder)
C0272978|Cerebral cortex laceration with open intracranial wound, with state of consciousness unspecified
C0272978|Cortex laceration with open intracranial wound, with state of consciousness unspecified
C0272979|Cortex (cerebral) laceration with open intracranial wound, with no loss of consciousness
C0272979|Cortex laceration with open intracranial wound and no loss of consciousness
C0272979|laceration of cerebrum with open intracranial wound with no loss of consciousness
C0272979|laceration of cerebrum with open intracranial wound with no loss of consciousness (diagnosis)
C0272979|Opn cortex lacer-no coma
C0272979|Cortex laceration with open intracranial wound AND no loss of consciousness (disorder)
C0272979|Cortex laceration with open intracranial wound, with no loss of consciousness
C0272979|Cortex laceration with open intracranial wound, with no loss of consciousness (disorder)
C0272979|Cerebral cortex laceration with open intracranial wound, with no loss of consciousness
C0272985|Cortex (cerebral) laceration with open intracranial wound, with concussion, unspecified
C0272985|laceration of cerebrum with open intracranial wound with concussion
C0272985|laceration of cerebrum with open intracranial wound with concussion (diagnosis)
C0272985|Opn cortx lacer-concuss
C0272985|Cortex laceration with open intracranial wound, with concussion, unspecified (disorder)
C0272985|Cortex laceration with open intracranial wound, with concussion, unspecified
C0272985|Cortex laceration with open intracranial wound AND concussion (disorder)
C0272985|Cortex laceration with open intracranial wound AND concussion
C0272985|Cortex laceration with open intracranial wound and unspecified concussion
C0272985|Cerebral cortex laceration with open intracranial wound, with concussion, unspecified
C1708044|Fetal Brain Injury
C0270088|Tentorial Tear
C0270088|Tentorial tear due to birth injury
C0270088|tentorial tear due to birth trauma
C0270088|tentorial tear due to birth trauma (diagnosis)
C0270088|Tears, Tentorial
C0270088|Tentorial Tears
C0270088|Tentorial laceration due to birth trauma
C0270088|Tentorial tear as birth trauma
C0270088|Tentorial tear as birth trauma (disorder)
C0270088|Tentorial tear due to birth trauma (disorder)
C0270088|birth; injury, tentorial tear
C0270088|injury; birth, tentorial tear
C2347482|Perinatal Brain Injury
C0478211|Other intracranial injuries
C0478211|Other intracranial injury
C0478211|[X]Other intracranial injuries (disorder)
C0478211|[X]Other intracranial injuries
C0238154|Epidural hemorrhage
C0238154|Epidural haemorrhage
C0238154|Extradural haematoma
C0238154|Extradural hemorrhage NOS
C0238154|Extradural Hemorrhage, Cranial
C0238154|Hematoma, Epidural, Intracranial
C0238154|Extradural Hematoma, Cranial
C0238154|Hematoma, Epidural, Cranial [Disease/Finding]
C0238154|Hemorrhage, Cranial Epidural
C0238154|Cranial Epidural Hematoma
C0238154|Hematoma, Epidural, Cranial
C0238154|Intracranial Epidural Hematoma
C0238154|Epidural Hemorrhage, Cranial
C0238154|Haemorrhage;epidural
C0238154|Haemorrhage;epidural;traumatic
C0238154|Epidural haematoma
C0238154|Epidural hematoma
C0238154|Epidural hemorrhage NOS
C0238154|Extradural hematoma
C0238154|Epidural hematoma (disorder)
C0238154|Epidural intracranial hemorrhage
C0238154|Epidural intracranial hematoma
C0238154|Epidural intracranial hemorrhage (disorder)
C0238154|Epidural intracranial haemorrhage
C0238154|Epidural hemorrhage (disorder)
C0238154|Epidural intracranial hematoma (disorder)
C0238154|Epidural intracranial haematoma
C0238154|Extradural haematoma (disorder)
C0238154|Extradural intracranial haematoma
C0238154|Extradural intracranial hematoma
C0238154|Hemorrhage, Extradural
C0238154|Extradural Hemorrhage
C0238154|Intracranial epidural haematoma
C0238154|Epidural bleeding
C0238154|Extradural haemorrhage
C0238154|EDH - Extradural haematoma
C0238154|EDH - Extradural hematoma
C0238154|epidural; hematoma
C0238154|extradural; hemorrhage
C0238154|hematoma; epidural
C0238154|hemorrhage; extradural
C0238154|Epidural hemorrhage, NOS
C0238154|Extradural hemorrhage, NOS
C0238154|Epidural hemorrhage [dup] (disorder)
C0238154|Cranial Epidural Hematomas
C0238154|Cranial Epidural Hemorrhages
C0238154|Cranial Epidural Hemorrhage
C0238154|Cranial Extradural Hematomas
C0238154|Cranial Extradural Hematoma
C0238154|Cranial Extradural Hemorrhages
C0238154|Cranial Extradural Hemorrhage
C0238154|Epidural Hematoma, Cranial
C0238154|Epidural Hematoma, Intracranial
C0238154|Epidural Hematomas, Cranial
C0238154|Epidural Hematomas, Intracranial
C0238154|Epidural Hemorrhages, Cranial
C0238154|Extradural Hematomas, Cranial
C0238154|Extradural Hemorrhages, Cranial
C0238154|Hematoma, Cranial Epidural
C0238154|Hematoma, Cranial Extradural
C0238154|Hematoma, Intracranial Epidural
C0238154|Hematomas, Cranial Epidural
C0238154|Hematomas, Cranial Extradural
C0238154|Hematomas, Intracranial Epidural
C0238154|Hemorrhage, Cranial Extradural
C0238154|Hemorrhages, Cranial Epidural
C0238154|Hemorrhages, Cranial Extradural
C0238154|Intracranial Epidural Hematomas
C0238154|Hemorrhage;epidural
C0238154|Hemorrhage;epidural;traumatic
C0238154|traumatic epidural hemorrhage
C0238154|traumatic epidural haemorrhage
C0452048|Intracranial injury with prolonged coma
C0452048|Intracranial injury with prolonged coma (diagnosis)
C0452048|intracranial injury unspecified nature with prolonged coma
C0452048|Intracranial injury with prolonged coma (disorder)
C0452048|injury; intracranial, with prolonged coma
C0452048|intracranial; injury, with prolonged coma
C0347535|Intracranial injury
C0347535|Intracranial injury, unspecified
C0347535|intracranial injury of unspecified nature
C0347535|intracranial injury of unspecified nature (diagnosis)
C0347535|unspecified intracranial injury (diagnosis)
C0347535|unspecified intracranial injury
C0347535|Injury;intracranial
C0347535|Intracranial injury (disorder)
C0347535|Intracranial injury NOS
C0347535|Intracranial injury NOS (disorder)
C0347535|[X]Intracranial injury, unspecified
C0347535|[X]Intracranial injury, unspecified (disorder)
C0347535|injury; intracranial
C0347535|intracranial; injury
C0347535|Intracranial injury [Ambiguous]
C0472391|Traumatic cerebral edema
C0472391|Traumatic cerebral oedema
C0472391|Traumatic cerebral edema NOS
C0472391|cerebral edema traumatic
C0472391|traumatic cerebral edema (diagnosis)
C0472391|Traumatic cerebral oedema (disorder)
C0472391|Traumatic cerebral edema (disorder)
C0472391|edema; brain, traumatic
C0475073|Traumatic subarachnoid haemorrhage
C0475073|Traumatic subarachnoid hemorrhage
C0475073|Hemorrhage, Post-Traumatic Subarachnoid
C0475073|Hemorrhages, Post-Traumatic Subarachnoid
C0475073|Post Traumatic Subarachnoid Hemorrhage
C0475073|Post-Traumatic Subarachnoid Hemorrhages
C0475073|Subarachnoid Hemorrhage, Post-Traumatic
C0475073|Subarachnoid Hemorrhages, Post-Traumatic
C0475073|Hemorrhage, Traumatic Subarachnoid
C0475073|Subarachnoid Hemorrhage, Traumatic
C0475073|Subarachnoid Hemorrhages, Traumatic
C0475073|Traumatic Subarachnoid Hemorrhages
C0475073|Post-Traumatic Subarachnoid Hemorrhage
C0475073|Subarachnoid Hemorrhage, Traumatic [Disease/Finding]
C0475073|Traumatic subarachnoid hemorrhage NOS
C0475073|Traumatic subarachnoid hemorrhage (disorder)
C0475073|Subarachnoid hemorrhage following injury
C0475073|Traumatic subarachnoid intracranial hemorrhage (disorder)
C0475073|Subarachnoid haemorrhage following injury
C0475073|Traumatic subarachnoid haemorrhage (disorder)
C0475073|Traumatic subarachnoid intracranial haemorrhage
C0475073|Traumatic subarachnoid intracranial hemorrhage
C0475073|hemorrhage; subarachnoid, traumatic
C0475073|subarachnoid; hemorrhage, traumatic
C1367166|Traumatic subdural haemorrhage
C1367166|Traumatic subdural hemorrhage
C1367166|head injury with subdural hemorrhage
C1367166|head injury with subdural hemorrhage (diagnosis)
C1367166|Haemorrhage;subdural;traumatic
C1367166|Traumatic subdural hemorrhage NOS
C1367166|Traumatic subdural intracranial hemorrhage
C1367166|Traumatic subdural intracranial haemorrhage
C1367166|Traumatic subdural intracranial hemorrhage (disorder)
C1367166|Traumatic subdural hemorrhage (disorder)
C1367166|Subdural haemorrhage following injury
C1367166|Subdural hemorrhage following injury
C1367166|hemorrhage; subdural, traumatic
C1367166|subdural; hemorrhage, traumatic
C1367166|Hemorrhage;subdural;traumatic
C2832047|Diffuse traumatic brain injury
C2832047|Diffuse traumatic brain injury NOS
C2832047|brain injury traumatic diffuse
C2832047|diffuse traumatic brain injury (diagnosis)
C2832052|Focal traumatic brain injury
C2832052|focal traumatic brain injury (diagnosis)
C2832052|brain injury traumatic focal
C2977736|Other specified intracranial injuries
C0272936|intracranial injury unspecified nature with open intracranial wound (diagnosis)
C0272936|intracranial injury unspecified nature with open intracranial wound
C0272936|intracranial injury of unspecified nature with open intracranial wound
C0272936|Brain injury with open intracranial wound (disorder)
C0272936|Brain injury with open intracranial wound
C0272936|Brain injury with open intracranial wound, NOS
C2118964|unspecified intracranial injury with no loss of consciousness (diagnosis)
C2118964|unspecified intracranial injury with no loss of consciousness
C2118964|unspecified intracranial injury with no LOC
C2118965|unspecified intracranial injury with brief (< 1 hr) loss of consciousness (diagnosis)
C2118965|unspecified intracranial injury brief (under 1 hr) unconsciousness
C2118965|unspecified intracranial injury with brief (< 1 hr) loss of consciousness
C2118965|unspecified intracranial injury with brief (< 1 hr) LOC
C2118965|unspecified intracranial injury with brief (under 1 hr) unconsciousness
C2118966|unspecified intracranial injury with moderate (1-24 hrs) loss of consciousness (diagnosis)
C2118966|unspecified intracranial injury moderate (1-24 hrs) unconsciousness
C2118966|unspecified intracranial injury with moderate (1-24 hrs) loss of consciousness
C2118966|unspecified intracranial injury with moderate (1-24 hrs) LOC
C2118966|unspecified intracranial injury with moderate (1-24 hrs) unconsciousness
C2118967|unspecified intracranial injury with prolonged (> 24 hrs) loss of consciousness with return to prior level of consciousness (diagnosis)
C2118967|unspecified intracranial injury loss of consciousness >24 hr then return to prior level
C2118967|unspecified intracranial injury with prolonged (> 24 hrs) loss of consciousness with return to prior level of consciousness
C2118967|unspecified intracranial injury with LOC over 24 hr, then return to prior level
C2118968|unspecified intracranial injury with prolonged (> 24 hrs) loss of consciousness without return to prior level of consciousness
C2118968|unspecified intracranial injury loss of consciousness > 24 hr without return to prior level
C2118968|unspecified intracranial injury with prolonged (> 24 hrs) loss of consciousness without return to prior level of consciousness (diagnosis)
C2118968|unspecified intracranial injury with LOC over 24 hours without return to prior level
C2118969|unspecified intracranial injury with unconsciousness of unspecified duration (diagnosis)
C2118969|unspecified intracranial injury with unconsciousness of unspecified duration
C2118970|unspecified intracranial injury with concussion (diagnosis)
C2118970|unspecified intracranial injury with concussion
C2832671|Unspecified intracranial injury without loss of consciousness
C2832675|Unspecified intracranial injury with loss of consciousness of 30 minutes or less
C2832679|Unspecified intracranial injury with loss of consciousness of 31 minutes to 59 minutes
C2832683|Unspecified intracranial injury with loss of consciousness of 1 hour to 5 hours 59 minutes
C2832687|Unspecified intracranial injury with loss of consciousness of 6 hours to 24 hours
C2832691|Unspecified intracranial injury with loss of consciousness greater than 24 hours with return to pre-existing conscious level
C2832695|Unspecified intracranial injury with loss of consciousness greater than 24 hours without return to pre-existing conscious level with patient surviving
C2832699|Unspecified intracranial injury with loss of consciousness of any duration with death due to brain injury prior to regaining consciousness
C2832703|Unspecified intracranial injury with loss of consciousness of any duration with death due to other cause prior to regaining consciousness
C2832707|Unspecified intracranial injury with loss of consciousness of unspecified duration
C0435306|open fracture of skull with intracranial injury (diagnosis)
C0435306|open skull fracture with intracranial injury
C0435306|open fracture of skull with intracranial injury
C0435306|Open fracture of skull NOS with intracranial injury
C0435306|Open fracture of skull NOS with intracranial injury (disorder)
C0435306|Open skull fracture with intracranial injury (disorder)
C0085094|Closed Head Injury
C0085094|Head Injuries, Closed
C0085094|Head Injury, Closed
C0085094|Closed head injuries
C0085094|HEAD INJ NONPENETRATING
C0085094|INJ CLOSED HEAD
C0085094|CLOSED HEAD INJ
C0085094|HEAD INJ CLOSED
C0085094|Closed Head Trauma
C0085094|Closed Head Traumas
C0085094|Head Traumas, Closed
C0085094|Trauma, Closed Head
C0085094|Traumas, Closed Head
C0085094|Nonpenetrating Head Injuries
C0085094|Nonpenetrating Head Injury
C0085094|Head Injuries, Nonpenetrating
C0085094|Head Trauma, Closed
C0085094|Head Injuries, Closed [Disease/Finding]
C0085094|Injuries, Closed Head
C0085094|Head Injury, Nonpenetrating
C0085094|Closed injury of head
C0085094|Closed injury of head (disorder)
C0085094|Injury;closed head
C3506613|injury of internal carotid artery, intracranial portion (diagnosis)
C3506613|injury of internal carotid artery, intracranial portion
C3506613|injury internal carotid artery intracranial portion
C3506611|unspecified intracranial injury with LOC with death due to brain injury prior to regaining consciousness (diagnosis)
C3506611|unspecified intracranial injury with LOC with death due to brain injury prior to regaining consciousness
C3506611|unspec intracranial injury loc w/ death d/t brain injury prior to regain consc
C3506612|unspec intracranial injury loc w/ death d/t other cause prior to regain consc (diagnosis)
C3506612|unspec intracranial injury loc w/ death d/t other cause prior to regain consc
C0161401|Injury of visual cortex
C0161401|injury of visual cortex (diagnosis)
C0161401|injury to the visual cortex
C0161401|Injury to visual cortex
C0161401|Injury of visual cortex NOS
C0161401|Traumatic injury of visual cortex
C0161401|Traumatic injury of visual cortex (disorder)
C0161401|Visual cortex injury
C0161401|Visual cortex injury (disorder)
C0161401|cortex; injury, visual
C0161401|injury; cortex, visual
C0161401|injury; visual cortex
C0161401|visual cortex; injury
C0270802|Spastic paralysis due to intracranial birth injury
C0270802|Spastic paralysis due to intracranial birth injury (disorder)
C0475075|Closed traumatic subarachnoid haemorrhage
C0475075|Closed traumatic subarachnoid hemorrhage
C0475075|Closed traumatic subarachnoid hemorrhage (disorder)
C0473821|Subdural haemorrhage due to birth injury
C0473821|Subdural hemorrhage due to birth injury
C0473821|subdural hemorrhage due to birth trauma
C0473821|subdural hemorrhage due to birth trauma (diagnosis)
C0473821|Subdural intracranial hemorrhage due to birth trauma (disorder)
C0473821|Subdural intracranial haemorrhage due to birth trauma
C0473821|Subdural intracranial hemorrhage due to birth trauma
C0473821|Subdural hemorrhage due to birth trauma (disorder)
C0473821|Subdural haemorrhage unspecified, due to birth trauma
C0473821|Subdural hemorrhage unspecified, due to birth trauma
C0473821|Subdural hemorrhage unspecified, due to birth trauma (disorder)
C0473821|Subdural haemorrhage due to birth trauma
C0475054|Open traumatic extradural haemorrhage
C0475054|Open traumatic extradural hemorrhage
C0475054|Open traumatic extradural hemorrhage (disorder)
C0475061|Closed traumatic subdural intracranial haemorrhage
C0475061|Closed traumatic subdural intracranial hemorrhage
C0475061|Closed traumatic subdural intracranial hemorrhage (disorder)
C0475061|Closed traumatic subdural hemorrhage (disorder)
C0475061|Subdural hemorrhage following injury without open intracranial wound
C0475061|Subdural haemorrhage following injury without open intracranial wound
C0475061|Subdural hemorrhage following injury without open intracranial wound (disorder)
C0475061|head injury - subdural hemorrhage without open intracranial wound
C0475061|subdural hemorrhage following head injury without open intracranial wound (diagnosis)
C0475061|subdural hemorrhage following head injury without open intracranial wound
C0475061|Closed traumatic subdural haemorrhage
C0475061|Closed traumatic subdural hemorrhage
C0475059|Hematoma, Traumatic Subdural
C0475059|Hematomas, Traumatic Subdural
C0475059|Subdural Hematomas, Traumatic
C0475059|Traumatic Subdural Hematoma
C0475059|Traumatic Subdural Hematomas
C0475059|Haematoma;subdural;traumatic
C0475059|Subdural Hematoma, Traumatic
C0475059|Traumatic subdural haematoma
C0475059|Traumatic subdural haematoma (disorder)
C0475059|Traumatic subdural hematoma (disorder)
C0475059|Traumatic subdural hematoma (diagnosis)
C0475059|subdural hematoma - traumatic
C0475059|Subdural hematoma (traumatic)
C0475059|Subdural haematoma (traumatic)
C0475059|Hematoma;subdural;traumatic
C0273487|olfactory nerve injury
C0273487|traumatic olfactory nerve injury
C0273487|olfactory nerve injury (diagnosis)
C0273487|traumatic olfactory nerve injury (diagnosis)
C0273487|Injury of olfactory [1st ] nerve
C0273487|Injuries, Olfactory Nerve
C0273487|Nerve Trauma, Olfactory
C0273487|Trauma, Olfactory Nerve
C0273487|Traumatic Olfactory Neuropathies
C0273487|First Nerve Palsy, Traumatic
C0273487|Palsy, Traumatic First-Nerve
C0273487|Olfactory Nerve Injuries
C0273487|First-Nerve Traumas
C0273487|Palsies, Traumatic First-Nerve
C0273487|Traumatic First-Nerve Palsies
C0273487|Traumas, First-Nerve
C0273487|Nerve Injury, Olfactory
C0273487|Nerve Traumas, Olfactory
C0273487|Neuropathy, Traumatic Olfactory
C0273487|Traumatic First Nerve Palsy
C0273487|First Nerve Trauma
C0273487|Olfactory Neuropathies, Traumatic
C0273487|Traumatic Olfactory Neuropathy
C0273487|Injury, Olfactory Nerve
C0273487|Nerve Injuries, Olfactory
C0273487|Trauma, First-Nerve
C0273487|Traumas, Olfactory Nerve
C0273487|First-Nerve Palsies, Traumatic
C0273487|Olfactory Nerve Traumas
C0273487|Neuropathies, Traumatic Olfactory
C0273487|Cranial Nerve I Injury
C0273487|First Cranial Nerve Injury
C0273487|Injury, First Cranial Nerve
C0273487|Olfactory Neuropathy, Traumatic
C0273487|First-Nerve Trauma
C0273487|Olfactory Nerve Injuries [Disease/Finding]
C0273487|Traumatic First-Nerve Palsy
C0273487|Olfactory Nerve Trauma
C0273487|First Cranial Nerve Injuries
C0273487|First-Nerve Palsy, Traumatic
C0273487|Injury, Cranial Nerve I
C0273487|Olfactory (1st) nerve injury
C0273487|Olfactory nerve injury (disorder)
C0273487|Injury of first cranial nerve
C0273487|Injury of olfactory nerve
C0273487|Injury to olfactory nerve
C0273487|Injury of olfactory nerve (disorder)
C0273487|injury; olfactory nerve
C0273487|n.olfactorius; injury
C0273487|Injury to 1st cranial nerve
C0475592|Subarachnoid haemorrhage due to birth injury
C0475592|Subarachnoid hemorrhage due to birth injury
C0475592|Intracranial subarachnoid haemorrhage due to birth injury
C0475592|Subarachnoid hemorrhage due to birth injury (disorder)
C0475592|Intracranial subarachnoid hemorrhage due to birth injury
C0475592|Intracranial subarachnoid hemorrhage due to birth injury (disorder)
C0475592|birth trauma subarachnoid hemorrhage
C0475592|subarachnoid hemorrhage due to birth trauma
C0475592|subarachnoid hemorrhage due to birth trauma (diagnosis)
C0475592|birth; injury, subarachnoid hemorrhage
C0433912|Injury of vertebral artery
C0433912|vertebral artery injury (diagnosis)
C0433912|vertebral artery injury
C0433912|Injury of vertebral artery (disorder)
C0433912|a.vertebralis; injury
C0433912|injury; vertebral artery
C0474996|Traumatic spinal subarachnoid hemorrhage
C0474996|hemorrhage subarachnoid traumatic spinal
C0474996|Traumatic spinal subarachnoid hemorrhage (diagnosis)
C0474996|Traumatic spinal subarachnoid haemorrhage
C0474996|Traumatic spinal subarachnoid hemorrhage (disorder)
C0433070|Crushing injury of head
C0433070|Crushing injury of head, part unspecified
C0433070|Crushing injury of skull and intracranial contents
C0433070|crush injury of head (diagnosis)
C0433070|crush injury head
C0433070|crush injury of head
C0433070|[X]Crushing injury of head, part unspecified
C0433070|[X]Crushing injury of head, part unspecified (disorder)
C0433070|Crushing injury of skull and intracranial contents (disorder)
C0433070|crushing injury; head
C0433070|head; crushing injury
C0272937|Brain injury with open intracranial wound and unspecified state of consciousness -RETIRED-
C0272937|Brain injury with open intracranial wound and unspecified state of consciousness
C0272937|Intracranial injury NOS with open intracranial wound, unspecified state of consciousness (disorder)
C0272937|Brain injury with open intracranial wound and unspecified state of consciousness (disorder)
C0272937|Intracranial injury NOS with open intracranial wound, unspecified state of consciousness
C0433774|Intracranial injury NOS with open intracranial wound, with more than 24 hours loss of consciousness and return to pre-existing conscious level
C0433774|Intracranial injury NOS with open intracranial wound, with more than 24 hours loss of consciousness and return to pre-existing conscious level (disorder)
C0433783|Intracranial injury NOS without mention of open intracranial wound, with more than 24 hours loss of consciousness and return to pre-existing conscious level
C0433783|Intracranial injury NOS without mention of open intracranial wound, with more than 24 hours loss of consciousness and return to pre-existing conscious level (disorder)
C0433769|Intracranial injury NOS with open intracranial wound (disorder)
C0433769|Intracranial injury NOS with open intracranial wound
C0433776|Intracranial injury NOS with open intracranial wound, with loss of consciousness of unspecified duration (disorder)
C0433776|Intracranial injury NOS with open intracranial wound, with loss of consciousness of unspecified duration
C0433784|Intracranial injury NOS without mention of open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious state
C0433784|Intracranial injury NOS without mention of open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious state (disorder)
C0433786|Intracranial injury NOS without mention of open intracranial wound, with concussion, unspecified
C0433786|Intracranial injury NOS without mention of open intracranial wound, with concussion, unspecified (disorder)
C0433780|Intracranial injury NOS without mention of open intracranial wound, with no loss of consciousness (disorder)
C0433780|Intracranial injury NOS without mention of open intracranial wound, with no loss of consciousness
C0433785|Intracranial injury NOS without mention of open intracranial wound, with loss of consciousness of unspecified duration (disorder)
C0433785|Intracranial injury NOS without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0433775|Intracranial injury NOS with open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious level
C0433775|Intracranial injury NOS with open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious level (disorder)
C0433782|Intracranial injury NOS without mention of open intracranial wound, with 1-24 hours loss of consciousness (disorder)
C0433782|Intracranial injury NOS without mention of open intracranial wound, with 1-24 hours loss of consciousness
C0433773|Intracranial injury NOS with open intracranial wound, with 1-24 hours loss of consciousness
C0433773|Intracranial injury NOS with open intracranial wound, with 1-24 hours loss of consciousness (disorder)
C0433779|Intracranial injury NOS without mention of open intracranial wound, unspecified state of consciousness (disorder)
C0433779|Intracranial injury NOS without mention of open intracranial wound, unspecified state of consciousness
C0272938|Brain injury with open intracranial wound and no loss of consciousness
C0272938|head injury with open intracranial wound with no loss of consciousness (diagnosis)
C0272938|head injury with open intracranial wound with no loss of consciousness
C0272938|Intracranial injury NOS with open intracranial wound, with no loss of consciousness (disorder)
C0272938|Intracranial injury NOS with open intracranial wound, with no loss of consciousness
C0272938|Brain injury with open intracranial wound AND no loss of consciousness (disorder)
C0433778|Intracranial injury NOS without mention of open intracranial wound (disorder)
C0433778|Intracranial injury NOS without mention of open intracranial wound
C0433781|Intracranial injury NOS without mention of open intracranial wound, with less than 1 hour loss of consciousness
C0433781|Intracranial injury NOS without mention of open intracranial wound, with less than 1 hour loss of consciousness (disorder)
C0433777|Intracranial injury NOS with open intracranial wound, with concussion, unspecified (disorder)
C0433777|Intracranial injury NOS with open intracranial wound, with concussion, unspecified
C0433772|Intracranial injury NOS with open intracranial wound, with less than 1 hours loss of consciousness (disorder)
C0433772|Intracranial injury NOS with open intracranial wound, with less than 1 hours loss of consciousness
C0272925|intracranial injury without skull fracture
C0272925|head injury unspecified intracranial injury without skull fracture
C0272925|intracranial injury without skull fracture (diagnosis)
C0272925|Head injury, without skull fracture
C0272925|Intracranial injury, without skull fracture (disorder)
C0272925|Intracranial injury, without skull fracture
C0272925|Head injury, NOS, without skull fracture
C0272925|Intracranial injury, NOS, without skull fracture
C0558400|H'ge - cerebral trauma
C0558400|Cerebral trauma
C0558400|cerebral trauma (diagnosis)
C0558400|Cerebral trauma (disorder)
C0411045|Cerebral injury due to birth trauma
C0411045|Cerebral injury due to birth trauma (disorder)
C0433855|brain injury traumatic burst lobe
C0433855|Burst lobe of brain
C0433855|Burst lobe of brain (diagnosis)
C0433855|Burst lobe of brain (disorder)
C0442857|Hypothalamic injury
C0442857|hypothalamic injury (diagnosis)
C0442857|Hypothalamic injury (disorder)
C0456045|brain laceration tentorial
C0456045|tentorial brain laceration
C0456045|tentorial brain laceration (diagnosis)
C0456045|Tentorial laceration
C0456045|Tentorial laceration (disorder)
C0435236|closed fracture of skull vault with intracranial injury
C0435236|closed fracture of skull vault with intracranial injury (diagnosis)
C0435236|Closed fracture of vault of skull with intracranial injury (disorder)
C0435236|Closed fracture of vault of skull with intracranial injury
C0435236|Fracture of vault of skull, closed with intracranial injury
C0435236|Closed fracture vault of skull with intracranial injury
C0435236|Closed fracture vault of skull with intracranial injury (disorder)
C0435223|open fracture of skull vault with intracranial injury
C0435223|open fracture of skull vault with intracranial injury (diagnosis)
C0435223|Open fracture of vault of skull with intracranial injury
C0435223|Open fracture of vault of skull with intracranial injury (disorder)
C0435223|Fracture of vault of skull, open with intracranial injury
C0435223|Open fracture vault of skull with intracranial injury
C0435223|Open fracture vault of skull with intracranial injury (disorder)
C0273058|head injury with intracranial hemorrhage
C0273058|head injury with intracranial hemorrhage (diagnosis)
C0273058|Hemorrhage, Traumatic Intracranial
C0273058|Hemorrhages, Traumatic Intracranial
C0273058|Intracranial Hemorrhage, Traumatic
C0273058|Intracranial Hemorrhages, Traumatic
C0273058|Traumatic Intracranial Hemorrhages
C0273058|Intracranial Hemorrhage, Traumatic [Disease/Finding]
C0273058|Traumatic Intracranial Hemorrhage
C0273058|Hemorrhage, Intracranial, Traumatic
C0273058|Intracranial hemorrhage following injury
C0273058|Traumatic intracranial haemorrhage (disorder)
C0273058|Intracranial hemorrhage following injury (disorder)
C0273058|Traumatic intracranial hemorrhage (disorder)
C0273058|Traumatic intracranial haemorrhage
C0273058|Intracranial haemorrhage following injury
C0273058|Traumatic intracranial bleeding
C0273058|Traumatic intracranial haemorrhage NOS
C0273058|Traumatic intracranial hemorrhage NOS
C0273058|hemorrhage; intracranial, traumatic
C0273058|hemorrhage; traumatic, intracranial
C0273058|intracranial; hemorrhage, traumatic
C0273058|traumatic; hemorrhage, intracranial
C0273058|Intracranial hemorrhage following injury, NOS
C1264285|Intracranial injury with loss of consciousness (disorder)
C1264285|Intracranial injury with loss of consciousness
C0435249|open fracture of base of skull with intracranial injury (diagnosis)
C0435249|open basilar skull fracture with intracranial injury
C0435249|open fracture of base of skull with intracranial injury
C0435249|Open fracture base of skull with intracranial injury (disorder)
C0435249|Open fracture base of skull with intracranial injury
C0435249|Fracture of base of skull, open with intracranial injury
C0435249|Open fracture of base of skull with intracranial injury (disorder)
C0435262|closed fracture of base of skull with intracranial injury (diagnosis)
C0435262|closed basilar skull fracture with intracranial injury
C0435262|closed fracture of base of skull with intracranial injury
C0435262|Closed fracture base of skull with intracranial injury (disorder)
C0435262|Closed fracture base of skull with intracranial injury
C0435262|Fracture of base of skull, closed with intracranial injury
C0435262|Closed fracture of base of skull with intracranial injury (disorder)
C0273098|Closed traumatic extradural hemorrhage
C0273098|Closed traumatic extradural haemorrhage
C0273098|Closed traumatic extradural hemorrhage (disorder)
C0273098|Extradural hemorrhage following injury without open intracranial wound (diagnosis)
C0273098|head injury - with extradural hemorrhage, without open intracranial wound
C0273098|Extradural hemorrhage following injury without open intracranial wound
C0273098|Extradural haemorrhage following injury without open intracranial wound
C0273098|Extradural hemorrhage following injury without open intracranial wound (disorder)
C0272499|multiple open fractures of skull or face with subarachnoid, subdural, or extradural hemorrhage (diagnosis)
C0272499|multi skull/face fractures open w/ subarachnoid, subdural, extradural hemorrhage
C0272499|multiple open fractures of skull or face with subarachnoid, subdural, or extradural hemorrhage
C0272499|Multiple open fractures of skull AND/OR face with subarachnoid, subdural AND/OR extradural haemorrhage
C0272499|Multiple open fractures of skull AND/OR face with subarachnoid, subdural AND/OR extradural hemorrhage (disorder)
C0272499|Multiple open fractures of skull AND/OR face with subarachnoid, subdural AND/OR extradural hemorrhage
C0272499|Multiple open fractures of skull and face with subarachnoid, subdural and extradural hemorrhage
C0161399|injury of optic chiasm
C0161399|injury of optic chiasm (diagnosis)
C0161399|injury to the optic chiasm
C0161399|Injury to optic chiasm
C0161399|Injury of optic chiasm (disorder)
C0161399|Optic chiasm injury
C0751814|INJ VASCULAR BRAIN
C0751814|VASCULAR INJ BRAIN
C0751814|BRAIN INJ VASCULAR
C0751814|Brain Vascular Injury
C0751814|Injury, Brain Vascular
C0751814|Injury, Vascular Brain
C0751814|Vascular Brain Injuries
C0751814|Vascular Brain Injury
C0751814|Brain Vascular Trauma
C0751814|Trauma, Brain Vascular
C0751814|Vascular Traumas, Brain
C0751814|Cerebrovascular Trauma
C0751814|Trauma, Cerebrovascular
C0751814|Brain Injury, Vascular
C0751814|Cerebrovascular Trauma [Disease/Finding]
C0751814|Injury, Vascular, Brain
C0751814|Vascular Injury, Brain
C0751814|Vascular Trauma, Brain
C0751814|cerebral vessels; injury
C0751814|injury; cerebral vessels
C0273106|open intracranial wound and extradural hemorrhage with concussion (diagnosis)
C0273106|open intracranial wound and extradural hemorrhage with concussion
C0273106|head injury with open intracranial wound and extradural hemorrhage with concussion
C0273106|Extradural hem-concuss
C0273106|Extradural hemorrhage following injury with open intracranial wound, with concussion, unspecified
C0273106|Extradural haemorrhage following injury with open intracranial wound, with concussion, unspecified
C0273106|Extradural hemorrhage following injury with open intracranial wound, with concussion, unspecified (disorder)
C0273106|Extradural hemorrhage following injury, with open intracranial wound, with concussion, unspecified
C0273106|Extradural haemorrhage following injury with open intracranial wound AND concussion
C0273106|Extradural hemorrhage following injury with open intracranial wound AND concussion (disorder)
C0273106|Extradural hemorrhage following injury with open intracranial wound AND concussion
C0273106|Extradural hemorrhage following injury with open intracranial wound and unspecified concussion
C0475077|head injury with subarachnoid hemorrhage with moderate (1-24 hrs) loss of consciousness
C0475077|head injury with subarachnoid hemorrhage with moderate (1-24 hrs) loss of consciousness (diagnosis)
C0475077|head injury with subarachnoid hemorrhage moderate (1-24 hr) loss of consciousness
C0475077|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with 1-24 hours loss of consciousness (disorder)
C0475077|Subarachnoid hemorrhage following injury without mention of open intracranial wound, with 1-24 hours loss of consciousness
C0475077|Subarachnoid haemorrhage following injury without mention of open intracranial wound, with 1-24 hours loss of consciousness
C0273070|head injury with open intracranial wound and intracranial hemorrhage
C0273070|open intracranial wound and hemorrhage (diagnosis)
C0273070|open intracranial wound and hemorrhage
C0273070|Intracranial hemorrhage following injury with open intracranial wound
C0273070|Intracranial haemorrhage following injury with open intracranial wound
C0273070|Intracranial hemorrhage following injury with open intracranial wound (disorder)
C0273087|Middle meningeal hemorrhage following injury
C0273087|Middle meningeal hemorrhage following injury (disorder)
C0273087|Middle meningeal haemorrhage following injury
C0273087|Middle meningeal hemorrhage following injury [dup] (disorder)
C0273104|Extradural hemorrhage following injury without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0273104|Extradural hem following inj, w/o ment of open intcran wound, with loc of unspec duration
C0273104|Extradural hem following inj, w/o ment of open intcran wound, with prol loc, w/o rtrn to pecl
C0273104|Extradural hem-deep coma
C0273104|Extradural hem-coma NOS
C0273104|Extradural hemorrhage following injury without mention of open intracranial wound, with prolonged [more than 24 hours] loss of consciousness without return to pre-existing conscious level
C0273104|Extradural hemorrhage following injury without mention of open intracranial wound, with loss of consciousness of unspecified duration (disorder)
C0273104|Extradural haemorrhage following injury without mention of open intracranial wound, with loss of consciousness of unspecified duration
C0273104|extradural hemorrhage following injury without open intracranial wound, with loss of consciousness (diagnosis)
C0273104|extradural hemorrhage following injury without open intracranial wound, with loss of consciousness
C0273104|head inj - w/ extradural hemorrhage, w/o open intracranial wound w/ loc
C0273104|Extradural haemorrhage following injury without open intracranial wound AND with loss of consciousness
C0273104|Extradural hemorrhage following injury without open intracranial wound AND with loss of consciousness (disorder)
C0273104|Extradural hemorrhage following injury without open intracranial wound AND with loss of consciousness
C0273104|Extradural hemorrhage following injury without open intracranial wound and with loss of consciousness of unspecified duration
C0475083|Subarachnoid haemorrhage following injury with open intracranial wound, with 1-24 hours loss of consciousness
C0475083|Subarachnoid hemorrhage following injury with open intracranial wound, with 1-24 hours loss of consciousness
C0475083|Subarachnoid hemorrhage following injury with open intracranial wound, with 1-24 hours loss of consciousness (disorder)
C0475082|Subarachnoid hemorrhage following injury with open intracranial wound, with less than 1 hour loss of consciousness
C0475082|Subarachnoid hemorrhage following injury with open intracranial wound, with less than 1 hour loss of consciousness (disorder)
C0475082|Subarachnoid haemorrhage following injury with open intracranial wound, with less than 1 hour loss of consciousness
C0475085|Subarachnoid hemorrhage following injury with open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious level
C0475085|Subarachnoid haemorrhage following injury with open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious level
C0475085|Subarachnoid hemorrhage following injury with open intracranial wound, with more than 24 hours loss of consciousness without return to pre-existing conscious level (disorder)
C0160228|head injury with open intracranial wound and subarachnoid hemorrhage (diagnosis)
C0160228|head injury with open intracranial wound and subarachnoid hemorrhage
C0160228|open intracranial wound and subarachnoid hemorrhage
C0160228|Subarachnoid hemorrhage following injury with open intracranial wound
C0160228|Subarachnoid haemorrhage following injury with open intracranial wound
C0160228|Subarachnoid hemorrhage following injury with open intracranial wound (disorder)
C0160233|Subarachnoid hemorrhage following injury with open intracranial wound and prolonged loss of consciousness (more than 24 hours) and return to pre-existing conscious level
C0160233|open intracranial wound and subarachnoid hemorrhage loss of consciousness greater than 24 hours then return to previous level
C0160233|open intracranial wound and subarachnoid hemorrhage with prolonged (> 24 hrs) loss of consciousness with return to prior level of consciousness (diagnosis)
C0160233|open intracranial wound and subarachnoid hemorrhage with prolonged (> 24 hrs) loss of consciousness with return to prior level of consciousness
C0160233|head injury with open intracranial wound and subarachnoid hemorrhage with LOC over 24 hr, then return to prior level
C0160233|Subarac hem following inj, with open intcran wound, with prolonged loc and return to pecl
C0160233|Op subarach hem-prol com
C0160233|Subarachnoid hemorrhage following injury with open intracranial wound, with prolonged [more than 24 hours) loss of consciousness and return to pre-existing conscious level
C0160233|Subarachnoid haemorrhage following injury with open intracranial wound, with more than 24 hours loss of consciousness and return to pre-existing conscious level
C0160233|Subarachnoid hemorrhage following injury with open intracranial wound, with more than 24 hours loss of consciousness and return to pre-existing conscious level
C0160233|Subarachnoid hemorrhage following injury with open intracranial wound, with more than 24 hours loss of consciousness and return to pre-existing conscious level (disorder)
C0160233|Subarachnoid haemorrhage following injury with open intracranial wound AND prolonged loss of consciousness (more than 24 hours) AND return to pre-existing conscious level
C0160233|Subarachnoid hemorrhage following injury with open intracranial wound AND prolonged loss of consciousness (more than 24 hours) AND return to pre-existing conscious level (disorder)
C0541931|Encephalitis toxic chronic
C0007789|Cerebral Palsy
C0007789|Cerebral palsy NOS
C0007789|Cerebral palsy, unspecified
C0007789|CP (Cerebral Palsy)
C0007789|Cerebral Palsy [Disease/Finding]
C0007789|cerebral palsy (diagnosis)
C0007789|Palsy;cerebral
C0007789|CP
C0007789|Cerebral palsy (CP)
C0007789|Cerebral palsy (disorder)
C0007789|Congenital cerebral palsy
C0007789|Infantile cerebral palsy
C0007789|Cerebral paralysis
C0007789|Palsy cerebral
C0007789|CP - Cerebral palsy
C0007789|cerebral; paralysis
C0007789|paralysis; cerebral
C0007789|Cerebral palsy, NOS
C0007789|Cerebral palsy [Ambiguous]
C0553767|CONGEN CEREBRAL PALSY
C0553767|Congenital cerebral palsy NOS (disorder)
C0553767|Congenital cerebral palsy
C0553767|Congenital cerebral palsy NOS
C0553767|cerebral palsy congenital
C0553767|Congenital cerebral palsy (diagnosis)
C0553767|Congenital cerebral palsy (disorder)
C0553767|Cerebral Palsy, Congenital
C0270719|Chatter-box syndrome
C0270719|Chronic brain-hydrocephalus syndrome
C0270719|Cocktail party syndrome
C0270719|Chronic brain-hydrocephalus syndrome (disorder)
C0270674|Chronic non-psychotic brain syndrome
C0270674|Chronic non-psychotic brain syndrome (disorder)
C0236656|alcohol-induced persistent dementia (diagnosis)
C0236656|alcohol-induced persistent dementia
C0236656|alcohol dependence with dementia (diagnosis)
C0236656|alcohol dependence with dementia
C0236656|Alcohol induced persisting dementia
C0236656|Alcohol persist dementia
C0236656|Dementia;alcoholic
C0236656|Alcoholic dementia NOS
C0236656|[X]Alcoholic dementia NOS
C0236656|[X]Chronic alcoholic brain syndrome
C0236656|Alcoholic dementia NOS (disorder)
C0236656|chronic organic mental disorder alcoholic brain syndrome
C0236656|Chronic alcoholic brain syndrome
C0236656|Chronic alcoholic brain syndrome (diagnosis)
C0236656|Dementia associated with alcoholism
C0236656|Alcohol-induced persisting dementia
C0236656|Alcoholic dementia
C0236656|Chronic alcoholic brain syndrome (disorder)
C0236656|Dementia associated with alcoholism (disorder)
C0236656|brain; syndrome, alcoholic (chronic)
C0236656|dementia; alcoholic
C0236656|dementia; alcohol
C0236656|alcohol; dementia
C0236656|syndrome; brain, alcoholic (chronic)
C0236656|Alcoholism associated with dementia NOS
C0019151|Encephalopathies, Hepatic
C0019151|Encephalopathies, Portosystemic
C0019151|Hepatic Encephalopathies
C0019151|Hepatic Encephalopathy
C0019151|Portosystemic Encephalopathies
C0019151|ENCEPH HEPATOCEREBRAL
C0019151|ENCEPH PORTAL SYSTEMIC
C0019151|HEPATIC ENCEPH
C0019151|PORTOSYSTEMIC ENCEPH
C0019151|ENCEPH PORTOSYSTEMIC
C0019151|PORTAL SYSTEMIC ENCEPH
C0019151|HEPATOCEREBRAL ENCEPH
C0019151|ENCEPH HEPATIC
C0019151|hepatic encephalopathy (diagnosis)
C0019151|Hepatocerebral encephalopathy -RETIRED-
C0019151|Encephalopathies, Hepatocerebral
C0019151|Hepatocerebral Encephalopathies
C0019151|Encephalopathies, Portal-Systemic
C0019151|Portal Systemic Encephalopathy
C0019151|Portal-Systemic Encephalopathies
C0019151|hepatic encephalopathy NOS
C0019151|Portosystemic Encephalopathy
C0019151|Encephalopathy, Hepatocerebral
C0019151|Hepatocerebral Encephalopathy
C0019151|Hepatic Encephalopathy [Disease/Finding]
C0019151|Portal-Systemic Encephalopathy
C0019151|Encephalopathy, Hepatic
C0019151|Encephalopathy, Portal-Systemic
C0019151|Encephalopathy, Portosystemic
C0019151|hepatic coma/encephalopathy
C0019151|Encephalopathy, Portal Systemic
C0019151|Gaustad's syndrome
C0019151|Portal systemic encephalopathy (disorder)
C0019151|Transient hepatargy syndrome
C0019151|Encephalopathy - hepatic
C0019151|Hepatocerebral encephalopathy (disorder)
C0019151|Encephalopathy hepatic
C0019151|HE - Hepatic encephalopathy
C0019151|Hepatic encephalopathy (disorder)
C0019151|encephalopathy; hepatic
C0019151|encephalopathy; portosystemic
C0019151|hepatic; encephalopathy
C0019151|portosystemic; encephalopathy
C2729507|hepatic encephalopathy with coma (diagnosis)
C2729507|hepatic encephalopathy with coma
C0019147|Comas, Hepatic
C0019147|Hepatic Comas
C0019147|Coma, Hepatic
C0019147|Hepatic coma
C0019147|Coma hepatic
C0019147|Hepatic coma NOS
C0019147|Coma;hepatic
C0019147|Hepatic coma (disorder)
C0019147|Hepatocerebral intoxication
C0019147|coma; hepatic
C0019147|hepatic; coma
C3266165|Hepatic encephalopathy in fulminant hepatic failure
C3266165|Hepatic encephalopathy in fulminant hepatic failure (disorder)
C0751198|Hepatic Stupors
C0751198|Stupor, Hepatic
C0751198|Stupors, Hepatic
C0751198|Hepatic Stupor
C1836797|COXPD1
C1836797|COMBINED OXIDATIVE PHOSPHORYLATION DEFICIENCY 1
C1836797|Hepatoencephalopathy, Early Fatal Progressive
C4024937|Chronic hepatic encephalopathy
