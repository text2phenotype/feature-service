C0079500|Hepatitis C-Like Viruses
C0220847|Hepatitis C virus
C0019196|Hepatitis C
C0220847|Hepatitis C virus
C3839041|Reactivation of hepatitis C viral hepatitis
C0369335|Hepatitis C virus RNA
C0400914|Acute hepatitis C
C0400920|Hepatitis C carrier (finding)
C1112419|Hepatitis C positive
C1698259|HCV coinfection
C0700073|hepatitis nonA nonB virus
C0700073|enterically-transmitted non-A, non-B hepatitis virus ET-NANBHV
C0700073|non-A non-B hepatitis virus
C0700073|non-A, non-B hepatitis virus ET-NANBHV
C0700073|non-A, non-B hepatitis-associated virus
C0700073|Non-A, non-B hepatitis virus
C0700073|Non-A, non-B hepatitis virus (organism)
C0376573|GB virus B
C0376573|Hepatitis GB virus B
C0376573|GBV-B
C0079500|Hepatitis C Like Viruses
C0079500|Hepatitis C-Like Virus
C0079500|Hepatitis C-Like Viruses
C0079500|Genus Hepacivirus
C0079500|Hepacavirus
C0079500|Hepacivirus
C0079500|Hepaciviruses
C0079500|Hepatitis C virus group
C0079500|Hepatitis C viruses
C0079500|Genus: Hepatitis C virus group
C0079500|Hepacavirus (organism)
C0079500|Genus Hepacivirus (organism)
C0079500|Hepacivirus (organism)
C3601684|unclassified Hepacivirus
C0220847|Hepatitis C virus
C0220847|Hepatitis C viruses
C0220847|Hepatitis C
C0220847|Hepatitis C virus (HCV)
C0220847|HCV
C0220847|hepatitis C virus HCV
C0220847|human hepatitis C virus
C0220847|human hepatitis C virus HCV
C0220847|human hepatitis virus C HCV
C0220847|post-transfusion hepatitis non A non B virus
C0220847|HCV - Hepatitis C virus
C0220847|Hepatitis C virus (organism)
C0220847|Virus-Hepatitis C
C3532919|Hepatitis C virus genotype 1 (organism)
C3532919|Hepatitis C virus genotype 1
C3532920|Hepatitis C virus genotype 2
C3532920|Hepatitis C virus genotype 2 (organism)
C3532921|Hepatitis C virus genotype 3 (organism)
C3532921|Hepatitis C virus genotype 3
C3532922|Hepatitis C virus genotype 4 (organism)
C3532922|Hepatitis C virus genotype 4
C3532923|Hepatitis C virus genotype 5 (organism)
C3532923|Hepatitis C virus genotype 5
C3532924|Hepatitis C virus genotype 6
C3532924|Hepatitis C virus genotype 6 (organism)
C3494961|Hepatitis C virus subtype 3b (organism)
C3494961|Hepatitis C virus subtype 3b
C3494962|Hepatitis C virus subtype 3a
C3494962|Hepatitis C virus subtype 3a (organism)
C3494958|Hepatitis C virus subtype 6a (organism)
C3494958|Hepatitis C virus subtype 6a
C3494966|Hepatitis C virus subtype 1a (organism)
C3494966|Hepatitis C virus subtype 1a
C3494964|Hepatitis C virus subtype 2a
C3494964|Hepatitis C virus subtype 2a (organism)
C3494959|Hepatitis C virus subtype 5a (organism)
C3494959|Hepatitis C virus subtype 5a
C3494963|Hepatitis C virus subtype 2b (organism)
C3494963|Hepatitis C virus subtype 2b
C3494965|Hepatitis C virus subtype 1b (organism)
C3494965|Hepatitis C virus subtype 1b
C3662864|Hepatitis C virus subtype 4
C3662864|Hepatitis C virus subtype 4 (organism)
C1989112|Hepatitis C virus c22p Ab &#x7C; bld-ser-plas
C0369335|Hepatitis C virus RNA
C0369335|Hepatitis C virus ribonucleic acid (substance)
C0369335|Hepatitis C virus ribonucleic acid
C0369335|Hepatitis C virus RNA (substance)
C1989101|Hepatitis C virus 100-3 Ab &#x7C; bld-ser-plas
C1989113|Hepatitis C virus c33c Ab &#x7C; bld-ser-plas
C3700145|Hepatitis C virus NS3 gene &#x7C; Isolate
C1989123|Hepatitis C virus sod Ab &#x7C; bld-ser-plas
C0166049|Anti HCV Antibodies
C0166049|Hepatitis C Antibodies
C0166049|ANTIHCV ANTIBODIES
C0166049|ANTIHEPATITIS C VIRUS ANTIBODIES
C0166049|Anti-HCV Antibodies
C0166049|Hepatitis C Antibodies [Chemical/Ingredient]
C0166049|Anti-Hepatitis C Virus Antibodies
C0166049|Hepatitis C Virus Antibodies
C0166049|HCV Antibodies
C0166049|Hepatitis C virus Ab
C0166049|Anti Hepatitis C Virus Antibodies
C0166049|Hepatitis C virus Antibody
C0166049|Anti-HCV Antibody
C0166049|Hepatitis C Antibody
C0166049|HCV Antibody
C0166049|Anti-Hepatitis C Antibody
C0166049|Anti HCV
C0166049|Antibody to hepatitis C
C0166049|Antibody to hepatitis C virus (substance)
C0166049|Antibody to hepatitis C virus
C2738068|Hepatitis C virus E2 Ab &#x7C; Bld-Ser-Plas
C1989099|Hepatitis C virus &#x7C; XXX
C2587456|Hepatitis C virus &#x7C; Body fluid
C1989097|Hepatitis C virus &#x7C; bld-ser-plas
C2738069|Hepatitis C virus NS3 Ab &#x7C; Bld-Ser-Plas
C2357726|Hepatitis C Virus C100p+5-1-1 Ab &#x7C; Bld-Ser-Plas
C1989102|Hepatitis C virus 22-3 Ab &#x7C; bld-ser-plas
C2357722|Hepatitis C virus 100+5-1-1 Ab &#x7C; Bld-Ser-Plas
C1989117|Hepatitis C virus NS5 Ab &#x7C; bld-ser-plas
C1989103|Hepatitis C virus 5-1-1 Ab &#x7C; bld-ser-plas
C2738067|Hepatitis C virus c2 Ab &#x7C; Bld-Ser-Plas
C3700146|Hepatitis C virus NS5 gene &#x7C; Isolate
C1989098|Hepatitis C virus &#x7C; Tissue and Smears
C2738066|Hepatitis C virus c1 Ab &#x7C; Bld-Ser-Plas
C2738070|Hepatitis C virus NS4 Ab &#x7C; Bld-Ser-Plas
C4068643|Hepatitis C virus core Antigen
C4068643|Hepatitis C virus core Ag
C0524910|Chronic viral hepatitis C
C0524910|Hepatitis C, Chronic
C0524910|chronic hepatitis, C virus
C0524910|chronic viral hepatitis C infection
C0524910|chronic hepatitis C infection (diagnosis)
C0524910|chronic hepatitis C infection
C0524910|Chronic Hepatitis C
C0524910|Hepatitis C, Chronic [Disease/Finding]
C0524910|Chronic viral hepatitis C (disorder)
C0524910|Chronic hepatitis C (disorder)
C0524910|Chronic type C viral hepatitis
C0524910|hepatitis; virus, chronic, type C
C0019196|Hepatitis C
C0019196|PT NANBH
C0019196|Viral hepatitis, non-A, non-B -RETIRED-
C0019196|viral hepatitis C infection
C0019196|hepatitis C infection (diagnosis)
C0019196|hepatitis C infection
C0019196|Hepatitis non-A non-B
C0019196|Unspecified viral hepatitis C
C0019196|Viral hepatitis C NOS
C0019196|Hepatitis C [Disease/Finding]
C0019196|PT-NANBH
C0019196|Parenterally-Transmitted Non-A, Non-B Hepatitis
C0019196|Hepatitis, Viral, Non-A, Non-B, Parenterally-Transmitted
C0019196|Parenterally Transmitted Non A, Non B Hepatitis
C0019196|Viral hepatitis, non-A, non-B
C0019196|Hepatitis C (disorder)
C0019196|Viral hepatitis, non-A, non-B (disorder)
C0019196|Viral hepatitis C (disorder)
C0019196|Viral hepatitis type C (disorder)
C0019196|Viral hepatitis type C
C0019196|Non-A non-B hepatitis
C0019196|Hep non-A non-B
C0019196|Viral hepatitis C
C0019196|Hepatitis (non-A non-B)
C0019196|Type C viral hepatitis
C0019196|Hepatitis non-A non-B (disorder)
C0019196|hepatitis nonA nonB
C0019196|hepatitis non A non B
C0019196|hepatitis; virus, non-A, non-B
C0019196|hepatitis; virus, type C
C0019196|non-A non-B-hepatitis
C0019196|virus; hepatitis, non-A, non-B
C0019196|Non-A, non-B hepatitis
C0019196|NANBH
C0019196|Unspecified viral hepatitis C NOS
C2711110|Hepatitis B and hepatitis C (disorder)
C2711110|Hepatitis B and hepatitis C
C2711110|Hepatitis B and hepatitis C (diagnosis)
C2711110|hepatitis viral b and c
C1456263|Hpt C w/o hepat coma NOS
C1456263|Unspecified viral hepatitis C without hepatic coma
C1456265|Hpt C w hepatic coma NOS
C1456265|Unspecified viral hepatitis C with hepatic coma
C2063424|chronic hepatitis C infection with hepatic coma (diagnosis)
C2063424|hepatitis, C virus with hepatic coma
C2063424|chronic viral hepatitis C infection with hepatic coma
C2063424|chronic hepatitis, C virus with hepatic coma
C2063424|hepatitis C infection with hepatic coma (diagnosis)
C2063424|hepatitis C infection with hepatic coma
C2063424|chronic hepatitis C infection with hepatic coma
C0400914|Acute hepatitis C
C0400914|acute viral hepatitis C infection
C0400914|acute hepatitis C infection (diagnosis)
C0400914|acute hepatitis C infection
C0400914|acute type C viral hepatitis
C0400914|Acute hepatitis C NOS
C0400914|Hepatitis C, acute
C0400914|Acute hepatitis C (disorder)
C0520788|posttransfusion hepatitis
C0520788|Hepatitis post transfusion
C0520788|Post transfusion hepatitis
C0520788|Posttransfusion viral hepatitis (disorder)
C0520788|Posttransfusion viral hepatitis
C0520788|Transfusion hepatitis
C0520788|hepatitis; post-transfusion
C0520788|post-transfusion; hepatitis
C0520788|Posttransfusion hepatitis, NOS
C0520788|Posttransfusion viral hepatitis, NOS
C0520788|Transfusion hepatitis, NOS
C0400900|Viral hepatitis C without mention of hepatic coma (disorder)
C0400900|Viral hepatitis C without mention of hepatic coma
C0375009|Chrnc hpt C w hepat Coma
C0375009|Chronic hepatitis C with hepatic coma
C0375009|Chronic viral hepatitis C with hepatic coma (disorder)
C0375009|Chronic viral hepatitis C with hepatic coma
C3837244|hepatitis, c virus - without hepatic coma
C3837244|hepatitis, C virus without hepatic coma
C3837244|hepatitis, C virus without hepatic coma (diagnosis)
C3839041|Reactivation of hepatitis C viral hepatitis (disorder)
C3839041|Reactivation of hepatitis C viral hepatitis
C0400915|Viral hepatitis C with coma
C0400915|Viral hepatitis C with coma (disorder)
C0241911|Chronic non-A non-B hepatitis
C0241911|Chronic non-A non-B hepatitis (disorder)
C0458009|Congenital hepatitis C infection
C0458009|Congenital hepatitis C infection (disorder)
C2357728|Hepatitis C virus RNA &#x7C; Body Fluid
C1989118|Hepatitis C virus RNA &#x7C; bld-ser-plas
C1989120|Hepatitis C virus RNA &#x7C; Cerebral spinal fluid
C1989119|Hepatitis C virus RNA &#x7C; Bone marrow
C1989121|Hepatitis C virus RNA &#x7C; Tissue and Smears
C1989122|Hepatitis C virus RNA &#x7C; XXX
C1545335|HIV 1+Hepatitis C virus RNA
C1545335|human immunodeficiency virus 1+Hepatitis C virus ribonucleic acid
C2911593|Acute hepatitis C without hepatic coma
C1456261|Hpt C acute w hepat Coma
C1456261|Acute hepatitis C with hepatic coma
C2215293|acute hepatitis C infection with hepatic coma
C2215293|acute hepatitis C infection with hepatic coma (diagnosis)
C2215293|acute type C viral hepatitis with hepatic coma
C2118423|acute hepatitis C infection with fulminant hepatic failure
C2118423|acute hepatitis C infection with fulminant hepatic failure (diagnosis)
C2118423|acute type C viral hepatitis with fulminant hepatic failure
C3838646|acute hepatitis, C virus without hepatic coma
C3838646|acute hepatitis, C virus without hepatic coma (diagnosis)
C3838646|hepatitis, c virus - acute without hepatic coma
C0400920|Hepatitis C carrier (finding)
C0400920|Hepatitis C carrier
C2025298|carrying viral hepatitis type C
C2025298|carrier of type C viral hepatitis
C2025298|carrier of type C viral hepatitis (history)
C1112419|Hepatitis C positive
C1698259|HCV coinfection
