C0005910|Body Weight
C0944911|Body weight:Mass:Point in time:^Patient:Quantitative
C0178684|human birth weight
C0028754|Obesity
C0028754|Obesity, unspecified
C0028754|obesity (diagnosis)
C0028754|Obesity NOS
C0028754|Obesity [Disease/Finding]
C0028754|Obesity (disorder)
C0028754|Med: Obesity
C0028754|Obese
C0028754|Obesity, NOS
C0028754|Obesity [Ambiguous]
C0028754|Obese (finding)
C1262477|Losses, Weight
C1262477|Reduction, Weight
C1262477|Reductions, Weight
C1262477|Weight Loss
C1262477|Weight Losses
C1262477|Weight Reductions
C1262477|Loss, Weight
C1262477|Weight decreased
C1262477|Progressive weight loss
C1262477|Weight loss, progressive
C1262477|Decreased weight
C1262477|Decreased body weight
C1262477|weight loss on exam (physical finding)
C1262477|weight loss on exam
C1262477|weight loss (on exam)
C1262477|Abnormal loss of weight
C1262477|Weight Loss [Disease/Finding]
C1262477|Weight Reduction
C1262477|Decreased;weight
C1262477|Loss (of);weight
C1262477|Weight decreasing
C1262477|Loss of weight
C1262477|Weight decreasing (finding)
C1262477|Weight loss finding
C1262477|Weight loss (finding)
C1262477|Weight loss finding (finding)
C1262477|Weight Decrease
C1262477|Lost weight
C1262477|Losing wt
C1262477|Wt loss
C1262477|Losing weight
C1262477|Weight decreased (finding)
C1262477|loss; weight
C1262477|weight; loss
C1262477|Weight decreased (observable entity)
C0596091|animal birth weight
C0043094|Gains, Weight
C0043094|Weight Gain
C0043094|Weight Gains
C0043094|Gain, Weight
C0043094|Weight increased
C0043094|Increased body weight
C0043094|weight gain (physical finding)
C0043094|Weight Gain [Disease/Finding]
C0043094|Increased;weight
C0043094|Increased weight
C0043094|Weight increasing
C0043094|Weight increasing (finding)
C0043094|Weight gain (finding)
C0043094|Weight gain finding
C0043094|Weight gain finding (finding)
C0043094|Body Weight Gain
C0043094|BWGAIN
C0043094|Weight Increase
C0043094|Ponderal increased
C0043094|Wt gain
C0043094|Weight increased (finding)
C0043094|Weight increased (observable entity)
C0005612|Birth Weight
C0005612|Birth Weights
C0005612|Weight, Birth
C0005612|Weights, Birth
C0005612|birth weight (physical finding)
C0005612|Birth Weight [Disease/Finding]
C0005612|Finding of birth weight
C0005612|Birth weight of baby NOS (finding)
C0005612|Observation of birth weight
C0005612|Birth weight of baby NOS
C0005612|Finding of birth weight (finding)
C0005612|Birth weight (observable entity)
C0005612|Birth weight of baby NOS (observable entity)
C0005612|Weight - baby
C0005612|BW - Birth weight
C0005612|Birth weight finding (finding)
C0005612|Birth weight finding
C0005612|Birth weight of baby
C0005612|Birth weight, NOS
C0005911|Body Weight Changes
C0005911|Body Weight Change
C0005911|Change, Body Weight
C0005911|Changes, Body Weight
C0005911|Weight Change, Body
C0005911|Weight Changes, Body
C0005911|Weight change
C0005911|Body Weight Changes [Disease/Finding]
C0005911|Weight change (observable entity)
C0005911|weight changes
C0039870|Thinness
C0039870|LEANNESS
C0039870|Thinness [Disease/Finding]
C0039870|Thin build
C0039870|Thin build (finding)
C0039870|Skinny build
C0039870|Thinness, NOS
C0751992|Body Weights, Fetal
C0751992|Fetal Body Weight
C0751992|Fetal Body Weights
C0751992|Fetal Weight
C0751992|Fetal Weights
C0751992|Weight, Fetal
C0751992|Weights, Fetal
C0751992|Fetal Weight [Disease/Finding]
C0751992|Body Weight, Fetal
C0497406|OVERWEIGHT
C0497406|overweight (diagnosis)
C0497406|overweight (physical finding)
C0497406|Overweight [Disease/Finding]
C0497406|Patient overweight
C0497406|Overweight (finding)
C0497406|overweight (BMI<30)
C0497406|Overweight (BMI 25-30)
C0005910|Body Weight
C0005910|Body Weights
C0005910|Weight, Body
C0005910|Weights, Body
C0005910|Weight
C0005910|weight (physical finding)
C0005910|Body Weight [Disease/Finding]
C0005910|Body weight - observation
C0005910|Body weight (observable entity)
C0005910|BW
C0005910|Body weight, NOS
C0005910|Body weight [dup] (observable entity)
C0005910|Weight (Body)
C0421272|ideal weight ___
C0421272|IBW (ideal body weight) ___
C0421272|ideal weight
C0421272|ideal body weight
C0421272|ideal body weight (physical finding)
C0421272|Body Weight, Ideal
C0421272|Weight, Ideal Body
C0421272|Ideal Body Masses
C0421272|Normal Body Weights
C0421272|Body Masses, Ideal
C0421272|Masses, Ideal Body
C0421272|Body Weights, Ideal
C0421272|Weight, Normal Body
C0421272|Mass, Ideal Body
C0421272|Weights, Ideal Body
C0421272|Body Weight, Normal
C0421272|Body Weights, Normal
C0421272|Body Mass, Ideal
C0421272|Ideal Body Weights
C0421272|Weights, Normal Body
C0421272|Body weight ideal
C0421272|Ideal body weight (finding)
C0421272|IDEALWT
C0421272|Ideal Body Mass
C0421272|Normal Body Weight
C0421272|IBW - Ideal body weight
C0421272|Ideal body weight (observable entity)
C2709005|Dry body weight
C2709005|Dry weight
C2709005|Dry body weight (observable entity)
C0041667|Underweight
C0041667|Low body weight
C0041667|Low weight
C0041667|underweight (diagnosis)
C0041667|the patient's weight was too low
C0041667|weight of patient too low (physical finding)
C0041667|weight of patient too low
C0041667|Excessive body weight loss (finding)
C0041667|Excessive body weight loss
C0041667|Patient underweight
C0041667|Underweight (finding)
C0041667|Excessive body weight loss (finding) [Ambiguous]
C2195744|bitemporal wasting
C2195744|bitemporal wasting (physical finding)
C2195744|bitemporal wasting was noted
C0517416|Weight percentile for age
C0517416|weight ___ percentile for age
C0517416|weight percentile for age (physical finding)
C2197572|weight proportional to height (physical finding)
C2197572|weight proportional to height
C2197572|the weight was proportional to the height
C2188871|usual weight (physical finding)
C2188871|usual weight
C0517417|Weight percentile for height
C0517417|weight ___ percentile for height
C0517417|weight percentile for height (physical finding)
C2012267|goal weight (___ lbs)
C2012267|goal weight in pounds
C2012267|goal weight in pounds (physical finding)
C2012267|goal weight
C2227317|body weight adjusted for prescription (physical finding)
C2227317|body weight adjusted for prescription
C2227317|adjusted body weight (for Rx)
C1439839|dry weight (physical finding)
C1439839|dry weight
C2266789|weight recorded
C2266789|weight recorded (physical finding)
C2266789|weight was recorded
C2203027|weight in wheelchair (___ lbs)
C2203027|weight in wheelchair
C2203027|weight in wheelchair (physical finding)
C0424680|skin fold thickness
C0424680|Skin-fold thickness (finding)
C0424680|thickness of skin fold
C0424680|thickness of skin fold (physical finding)
C0424680|Skin-fold thickness
C0424680|Skin-fold thickness (observable entity)
C0006625|Cachexia
C0006625|[D]Cachexia (context-dependent category)
C0006625|[D]Cachexia NOS (context-dependent category)
C0006625|cachectic (physical finding)
C0006625|cachectic
C0006625|Cachexia [Disease/Finding]
C0006625|[D]Cachexia
C0006625|Cachexia (disorder)
C0006625|[D]Cachexia NOS (situation)
C0006625|[D]Cachexia (situation)
C0006625|[D]Cachexia NOS
C0006625|Wasting
C0006625|General body deterioration
C0006625|Cachexia (finding)
C0006625|Cachexia, NOS
C0006625|Cachexia (disorder) [Ambiguous]
C2230143|obesity (10+% over ideal weight)
C2230143|obesity (more than 10% over ideal weight) (physical finding)
C2230143|obesity (more than 10% over ideal weight)
C2230143|patient was observed to be obese
C2203039|weight within normal limits (+/- 10% ideal weight) (physical finding)
C2203039|weight within normal limits (+/- 10% ideal weight)
C2203028|weight less than 75% ideal body weight
C2203028|weight less than 75% ideal body weight (physical finding)
C0424631|Decreased subcutaneous fat
C0424631|Sparse subcutaneous fat
C0424631|Little subcutaneous fat
C0424631|Loss of subcutaneous fat
C0424631|loss of subcutaneous fat (physical finding)
C0424631|Subcutaneous fat loss
C0424631|Loss of subcutaneous fat (finding)
C2983672|Terminal Body Weight
C2983672|TERMBW
C1303013|Baseline weight (observable entity)
C1303013|Baseline weight
C0424662|Reference weight
C0424662|Reference weight (observable entity)
C3645728|weight obtained from prior medical record (___ lbs) (physical finding)
C3645728|weight obtained from prior medical record (___ lbs)
C1975565|Weight &#x7C; calculus (stone)
C1830806|Wt Wat Qn
C1830806|Weight:Mass:Pt:Water:Qn
C1830806|Weight of Water
C1830806|Weight:Mass:Point in time:Water:Quantitative
C3834630|weight with clothes (physical finding)
C3834630|weight with clothes
C3834629|weight without clothes (physical finding)
C3834629|weight without clothes
C3834631|weight at initial encounter ___
C3834631|weight at initial encounter ___ (physical finding)
C2751656|Slender habitus
C2751656|slender habitus (physical finding)
C4032003|antepartum weight (___lbs)
C4032003|antepartum weight
C4032003|antepartum weight (physical finding)
C4027960|weight post-surgery (___ lbs)
C4027960|post-surgery weight (physical finding)
C4027960|post-surgery weight
C4027367|weight pre-surgery (___ lbs)
C4027367|weight pre-surgery (___ lbs) (physical finding)
C4042910|Body Weight Maintenance
C4042910|Weight Maintenances, Body
C4042910|Maintenance, Body Weight
C4042910|Maintenances, Body Weight
C4042910|Body Weight Maintenances
C4042910|Weight Maintenance, Body
C1827199|Body weight without shoes
C1827199|Body weight without shoes (observable entity)
C1828456|Body weight with shoes (observable entity)
C1828456|Body weight with shoes
C0944911|Body weight:Mass:Point in time:^Patient:Quantitative
C0944911|Body weight:Mass:Pt:^Patient:Qn
C0944911|Weight
C0944911|Body weight
