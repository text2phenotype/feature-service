C0024117|Chronic Obstructive Airway Disease
C0034067|Emphysema
C0034067|Pulmonary Emphysema
C0034067|Emphysema, unspecified
C0034067|EMPHYSEMAS PULM
C0034067|EMPHYSEMA PULM
C0034067|PULM EMPHYSEMAS
C0034067|PULM EMPHYSEMA
C0034067|emphysema (diagnosis)
C0034067|Emphysema (lung)(pulmonary) NOS
C0034067|Emphysemas, Pulmonary
C0034067|Pulmonary Emphysemas
C0034067|Pulmonary Emphysema [Disease/Finding]
C0034067|Emphysema, Pulmonary
C0034067|Emphysema (disorder)
C0034067|Emphysema pulmonary
C0034067|Emphysema of lung
C0034067|Pulmonary emphysema (disorder)
C0034067|Emphysema of lung, NOS
C0034067|Pulmonary emphysema, NOS
C0034067|Emphysema (Pulmonary)
C0008677|Unspecified chronic bronchitis
C0008677|chronic bronchitis
C0008677|chronic bronchitis (diagnosis)
C0008677|Chronic bronchitis NOS
C0008677|Bronchitis, Chronic
C0008677|Bronchitis, Chronic [Disease/Finding]
C0008677|Bronchitis;chronic
C0008677|Chronic bronchitis (disorder)
C0008677|Chronic bronchitis NOS (disorder)
C0008677|-- Chronic Bronchitis
C0008677|Chronic bronchitis, unspecified
C0008677|Bronchitis chronic
C0008677|Bronchitis chronic NOS
C0008677|bronchitis; chronic
C0008677|chronic; bronchitis
C0008677|Chronic bronchitis, NOS
C0004096|Asthma
C0004096|Asthmas
C0004096|Asthma, unspecified
C0004096|Bronchial asthma
C0004096|asthma (diagnosis)
C0004096|Br. asthma
C0004096|Asthma NOS
C0004096|Unspecified asthma
C0004096|Asthma [Disease/Finding]
C0004096|Asthma, Bronchial
C0004096|Asthma (disorder)
C0004096|Asthma unspecified (disorder)
C0004096|Asthma NOS (disorder)
C0004096|Asthma unspecified
C0004096|-- Asthma
C0004096|Asthmatic
C0004096|Asthma bronchial
C0004096|Bronchitic asthma
C0004096|Cardio/pulm: Asthma
C0004096|Airway hyperreactivity
C0004096|Asthma, NOS
C0004096|Bronchial asthma, NOS
C0004096|Asthma (disorder) [Ambiguous]
C0006266|Bronchial Spasm
C0006266|Bronchial Spasms
C0006266|Bronchospasm
C0006266|Bronchospasms
C0006266|Spasm, Bronchial
C0006266|Spasms, Bronchial
C0006266|Bronchospasm NOS
C0006266|Broncho spasms
C0006266|bronchospasm (diagnosis)
C0006266|Bronchial Spasm [Disease/Finding]
C0006266|Bronchospasm (disorder)
C0006266|Spasm bronchial
C0006266|Bronchospasm (finding)
C0006266|bronchus; constriction
C0006266|bronchus; spasm
C0006266|constriction; bronchus
C0006266|spasm; bronchial
C0024117|COPD
C0024117|Pulmonary Disease, Chronic Obstructive
C0024117|CHRONIC OBSTRUCTIVE PULMONARY DISEASE
C0024117|Chronic Obstructive Airway Disease
C0024117|Chronic obstructive pulmonary disease, unspecified
C0024117|Chronic Obstructive Lung Disease
C0024117|Chronic Obstructive Airways Disease
C0024117|CHRONIC OBSTRUCTIVE LUNG DIS
C0024117|PULM DIS CHRONIC OBSTRUCTIVE
C0024117|CHRONIC OBSTRUCTIVE PULM DIS
C0024117|CHRONIC OBSTRUCTIVE AIRWAY DIS
C0024117|small airways disease
C0024117|COLD (chronic obstructive lung disease)
C0024117|chronic obstructive pulmonary disease (diagnosis)
C0024117|Chronic Obstructive Pulmonary Disease (COPD)
C0024117|COLD
C0024117|Chronic obstructive airway disease NOS
C0024117|Chronic obstructive lung disease NOS
C0024117|Pulmonary Disease, Chronic Obstructive [Disease/Finding]
C0024117|COAD
C0024117|Chronic airways disease
C0024117|Chronic obstructive airways disease NOS (disorder)
C0024117|Chronic obstructive lung disease (disorder)
C0024117|Chronic obstructive airways disease NOS
C0024117|Chronic obstructive pulmonary disease NOS
C0024117|-- COPD
C0024117|Obstructive Pulmonary Disease (COPD), Chronic
C0024117|COPD, Chronic Obstructive Pulmonary Disease
C0024117|Pulmonary Disease (COPD), Chronic Obstructive
C0024117|Chronic Obstructive Pulmonary Disease, (COPD)
C0024117|Disease (COPD), Chronic Obstructive
C0024117|Chronic obstructive pulmonary disease finding
C0024117|Chronic obstructive pulmonary disease finding (finding)
C0024117|Chronic obstruct airways disease
C0024117|Chronic obstructive bronchopneumopathy
C0024117|Hyperactive airway disease
C0024117|Obstructive airways disease (chronic)
C0024117|Chronic airflow limitation
C0024117|Chronic airway obstruction
C0024117|COAD - Chronic obstructive airways disease
C0024117|COLD - Chronic obstructive lung disease
C0024117|COPD - Chronic obstructive pulmonary disease
C0024117|Chronic airway disease
C0024117|Chronic irreversible airway obstruction
C0024117|CAFL - Chronic airflow limitation
C0024117|CAL - Chronic airflow limitation
C0024117|disease (or disorder); respiratory tract, chronic, obstructive
C0024117|disease (or disorder); respiratory tract, obstructive, chronic
C0024117|lung; disease, obstructive (chronic)
C0024117|lung; obstruction, disease, chronic
C0024117|obstruction; airway, chronic
C0024117|obstruction; lung, disease, chronic
C0024117|airway; obstruction, chronic
C0024117|respiratory tract; disorder, chronic, obstructive
C0024117|respiratory tract; disorder, obstructive, chronic
C0024117|Chronic obstructive lung disease, NOS
C0024117|Chronic obstructive lung disease [Ambiguous]
C0024117|Chronic airway obstruction; not otherwise specified
C0024117|COPD NOS
C0024117|Chronic obstr airways disease
C0024117|Chronic obstr lung disease
C0024117|Chronic obstr pulmon disease
C0006267|Bronchiectases
C0006267|Bronchiectasis
C0006267|bronchiectasis (diagnosis)
C0006267|Bronchiectasis NOS
C0006267|Bronchiectasis [Disease/Finding]
C0006267|Bronchiectasis NOS (disorder)
C0006267|Bronchiectasis (disorder)
C0006267|Chronic dilatation of bronchus and bronchiole
C0006267|Bronchi dilated
C0006267|Cardio/pulm: Bronchiectasis
C0006267|Bronchiectasis, NOS
C0375334|chronic obstructive asthma with status asthmaticus
C0375334|chronic obstructive asthma with status asthmaticus (diagnosis)
C0375334|Ch ob asthma w stat asth
C0348818|Chronic obstructive pulmonary disease with acute lower respiratory infection
C0348818|Chronic obstructive pulmon disease w acute lower resp infct
C0348818|chronic obstructive pulmonary disease with acute lower respiratory infection (diagnosis)
C0348818|Chronic obstructive pulmonary disease with acute lower respiratory infection (disorder)
C3508933|chronic obstructive pulmonary disease with exacerbation (diagnosis)
C3508933|chronic obstructive pulmonary disease with exacerbation
C1527303|Airflow Obstructions, Chronic
C1527303|Chronic Airflow Obstructions
C1527303|Chronic Airflow Obstruction
C1527303|CAO - Chronic airflow obstruction
C1527303|Airflow Obstruction, Chronic
C3714496|Allergic bronchiolitis
C3714496|Reactive airway disease
C3714496|Small airway disease
C3714496|Recurrent airway obstruction
C3714496|Recurrent airway obstruction (disorder)
C3714496|Chronic airway disease
C3714496|Heaves
C3714496|COPD
C3714496|Chronic obstructive pulmonary disease of horses
C3714496|Broken wind
C3714496|Chronic alveolar emphysema of horses
C3714496|Heaves (disorder)
C0348693|Other specified chronic obstructive pulmonary disease
C0348693|Other specified chronic obstructive airways disease
C0348693|[X]Other specified chronic obstructive pulmonary disease (disorder)
C0348693|Other specified chronic obstructive airways disease (disorder)
C0348693|[X]Other specified chronic obstructive pulmonary disease
C0155874|Obstructive chronic bronchitis
C0155874|Chronic obstructive bronchitis
C0155874|chronic bronchitis with emphysema
C0155874|Emphysematous bronchitis
C0155874|Chronic obstructive bronchitis (disorder)
C0155874|Obstructive chronic bronchitis NOS (disorder)
C0155874|Emphysematous bronchitis (disorder)
C0155874|Obstructive chronic bronchitis NOS
C0155874|Bronchitis with airway obstruction
C0155874|COB - Chronic obstructive bronchitis
C0155874|bronchitis; chronic, obstructive
C0155874|bronchitis; emphysematous
C0155874|chronic; bronchitis, obstructive
C0155874|emphysematous; bronchitis
C0155874|Chronic obstructive bronchitis (disorder) [Ambiguous]
C0155874|Chronic bronchitis & emphysema
C0155874|Emphysema with chronic bronchitis
C0155874|Chronic bronchitis, obstructive
C0155874|Bronchitis with emphysema
C0155874|Bronchitis, emphysematous
C0730607|Severe chronic obstructive pulmonary disease
C0730607|Severe chronic obstructive pulmonary disease (disorder)
C0730607|Severe chronic obstructive pulmonary disease (diagnosis)
C0730607|chronic obstructive pulmonary disease severe
C0730604|Mild chronic obstructive pulmonary disease
C0730604|Mild chronic obstructive pulmonary disease (disorder)
C0730604|chronic obstructive pulmonary disease mild
C0730604|Mild chronic obstructive pulmonary disease (diagnosis)
C0730605|Moderate chronic obstructive pulmonary disease (disorder)
C0730605|Moderate chronic obstructive pulmonary disease
C0730605|chronic obstructive pulmonary disease moderate
C0730605|Moderate chronic obstructive pulmonary disease (diagnosis)
C3662842|Chronic obstructive airway disease with asthma (disorder)
C3662842|Chronic obstructive airway disease with asthma
C1847014|PULMONARY DISEASE, CHRONIC OBSTRUCTIVE, SEVERE EARLY-ONSET
C0494659|Other chronic obstructive pulmonary disease
C0494660|Predominantly allergic asthma
C0494660|allergic (predominantly) asthma
C0494660|asthma; predominantly allergic
C0494660|predominantly allergic; asthma
C0029607|Other emphysema
C0029607|Emphysema NEC
C0029607|Other emphysema (morphologic abnormality)
C0029607|Other emphysema NOS
C0029607|[X]Other emphysema
C0029607|[X]Other emphysema (morphologic abnormality)
C0029607|Other emphysema NOS (morphologic abnormality)
C0849659|Chronic airways limitation
C0348817|Chronic obstructive pulmonary disease with acute exacerbation, unspecified
C0348817|Chronic obstructive pulmonary disease with acute exacerbation, unspecified (disorder)
C0348819|Mixed asthma
C0348819|asthma mixed
C0348819|mixed asthma (diagnosis)
C0348819|Mixed asthma (disorder)
C0348819|asthma; mixed
C0348819|mixed; asthma
C0221227|Centrilobular emphysema
C0221227|centriacinar emphysema (diagnosis)
C0221227|centriacinar emphysema
C0221227|Emphysema, Centrilobular
C0221227|Emphysemas, Centriacinar
C0221227|Centriacinar Emphysemas
C0221227|Emphysema, Centriacinar
C0221227|Centrilobular Emphysemas
C0221227|Emphysemas, Centrilobular
C0221227|Centriacinar emphysema (disorder)
C0221227|centrilobular; emphysema
C0221227|emphysema; centrilobular
C0221227|Lung or pulmonary emphysema, centriacinar
C0221227|Lung or pulmonary emphysema, centrilobular
C0264393|Panlobular emphysema
C0264393|panacinar emphysema
C0264393|panacinar emphysema (diagnosis)
C0264393|Panlobular Emphysemas
C0264393|Panacinar Emphysemas
C0264393|Emphysemas, Panlobular
C0264393|Emphysema, Panacinar
C0264393|Emphysemas, Panacinar
C0264393|Emphysema, Panlobular
C0264393|Alveolar emphysema of lung
C0264393|Vesicular emphysema
C0264393|Panacinar emphysema (disorder)
C0264393|emphysema; panacinar
C0264393|emphysema; panlobular
C0264393|emphysema; vesicular
C0264393|panacinar; emphysema
C0264393|panlobular; emphysema
C0264393|vesicular; emphysema
C0264393|Emphysema, vesicular
C0264393|Lung or pulmonary emphysema, panacinar
C0264393|Lung or pulmonary emphysema, panlobular
C0264393|Lung or pulmonary emphysema, vesicular
C0155880|Nonallergic asthma
C0155880|Intrinsic asthma
C0155880|intrinsic asthma (diagnosis)
C0155880|intrinsic nonallergic asthma
C0155880|Intrinsic asthma (disorder)
C0155880|Intrinsic asthma NOS
C0155880|Intrinsic asthma NOS (disorder)
C0155880|Non-allergic asthma
C0155880|Non-allergic asthma (diagnosis)
C0155880|asthma non-allergic
C0155880|Asthma due to internal immunological process
C0155880|Non-allergic asthma (disorder)
C0155880|asthma; intrinsic, nonallergic
C0155880|asthma; intrinsic
C0155880|asthma; nonallergic
C0155880|intrinsic; asthma, nonallergic
C0155880|intrinsic; asthma
C0155880|nonallergic; asthma
C0155880|Intrinsic asthma (disorder) [Ambiguous]
C1277261|end stage chronic obstructive pulmonary disease
C1277261|end stage chronic obstructive pulmonary disease (diagnosis)
C1277261|chronic obstructive pulmonary disease end stage
C1277261|End stage chronic obstructive airways disease (disorder)
C1277261|End stage chronic obstructive airways disease
C1854729|MUCUS INSPISSATION OF RESPIRATORY TRACT
C1969833|COPD, SEVERE EARLY-ONSET
C3714497|Reactive airway disease
C3714497|reactive airway disease (diagnosis)
C3714497|Reactive airway disease (disorder)
C3714497|Hyperactive Airway Disease
C3714497|Reactive airways disease
C3714497|Reactive Airway Disease (AQ)
C3714497|Disease;hyperactive airways
C3714497|hyperactive airways disease
C3838076|chronic obstructive pulmonary disease susceptibility
C3838076|COPD susceptibility
C3838076|COPD susceptibility (diagnosis)
C3838076|PULMONARY DISEASE, CHRONIC OBSTRUCTIVE, SUSCEPTIBILITY TO
C4040148|Chronic obstructive lung disease co-occurrent with acute bronchitis (disorder)
C4040148|Chronic obstructive lung disease co-occurrent with acute bronchitis
C0340044|Chronic obstructive pulmonary disease with (acute) exacerbation
C0340044|Chronic obstructive pulmonary disease w (acute) exacerbation
C0340044|Acute exacerbation of chronic obstructive airways disease (disorder)
C0340044|Acute exacerbation of chronic obstructive airways disease
C0340044|Acute exacerbation of COPD
C0340044|Acute exacerbation of chronic obstructive pulmonary disease
C0006272|Bronchiolitis Obliterans
C0006272|Obliterative bronchiolitis
C0006272|BO
C0006272|bronchiolitis obliterans (diagnosis)
C0006272|obliterative bronchiolitis (diagnosis)
C0006272|Bronchiolitis Obliterans [Disease/Finding]
C0006272|Obliterative bonchiolitis
C0006272|OB - Obliterative bronchiolitis
C0006272|Obliterative bronchiolitis (disorder)
C0006272|bronchiolitis; obliterative
C0006272|obliterative; bronchiolitis
C0006272|Obliterative bronchiolitis, NOS
C1385064|disease (or disorder); lung, obstructive (chronic)
C0001883|Airway Obstruction
C0001883|Airway Obstructions
C0001883|Obstruction, Airway
C0001883|Obstructions, Airway
C0001883|airway obstructed
C0001883|obstructed airway
C0001883|airway obstructed (physical finding)
C0001883|Airway Obstruction [Disease/Finding]
C0001883|Respiratory obstruction
C0001883|Airways obstruction
C0001883|Airway obstruction NOS
C0001883|Embarrassed airway
C0001883|Respiratory obstruction (disorder)
C0001883|obstruction; airway
C0001883|obstruction; respiratory
C0001883|airway; obstruction
C0001883|respiratory; obstruction
C0001883|Airway obstruction, NOS
C0155883|Chronic obstructive asthma
C0155883|chronic obstructive asthma (diagnosis)
C0155883|Chronic obstructive asthma (with obstructive pulmonary disease)
