C0086287|Females
C0086287|Female
C0086287|Woman
C0086287|W
C0086582|Males
C0086582|Male
C0086582|Man
C0086582|M
C1550327|Administrative Gender
C0079399|Gender
C1522384|sex
C1706180|Male Gender, Self Report
C1710069|Sex or Gender
C3839079|Masculine gender
C3839293|Feminine gender
C0043210|Women
C0043210|Human Females
C0043210|Woman
C0043210|Woman (person)
C0043210|Females (Human)
C0043210|Human, Female
C0015671|Father
C0015671|Fathers
C0015671|Father (person)
C0015671|Father, NOS
C0025266|Men
C0025266|Male population group
C0025266|Man
C0025266|Man (person)
C0025266|Human, Male
C0682275|House husband (context-dependent category)
C0682275|House husband (person)
C0682275|House husband
C0682275|House husband (situation)
C0682275|House husband (occupation)
C0242658|Homosexuality, Male
C0242658|Male Homosexuality
C0242658|Male homosexual state
C0242658|Male homosexual
C0242658|Male homosexual (finding)
C0043174|Widower
C0043174|Widower (person)
C0043174|Widowerhood
C0043174|Widower (finding)
C0043174|Widowers
C0521319|Boyfriend
C0521319|Boyfriend (person)
C0337527|brother
C0337527|Brother (person)
C0337527|Brothers
C0337527|Brother, NOS
C0037683|Son
C0037683|Son (person)
C0037683|Sons
C0037683|Son, NOS
C0086582|Male
C0086582|Human Males
C0086582|M
C0086582|Male Gender
C0086582|Male Gender [Disease/Finding]
C0086582|Male (finding)
C0086582|Males
C0086582|Male individual
C0086582|Male structure (body structure)
C0086582|Male structure
C0086582|Male individual, NOS
C0086582|Male, NOS
C0086582|Males (Human)
C0086582|Human, Male
C0432475|XX Male
C0432475|male with 46,XX karyotype
C0432475|male with 46,XX karyotype (diagnosis)
C0432475|XX males
C0432475|Male with 46, XX karyotype
C0432475|XX males (disorder)
C0432475|karyotype; 46,XX, male
C0458452|Male urethra
C0458452|Male urethral structure
C0458452|Male urethral structure (body structure)
C1291683|Male reproductive finding (finding)
C1291683|Male reproductive finding
C3687554|Intact male
C3687554|Intact male (finding)
C1319065|Castrated Male
C1319065|Neutered Male
C1319065|Neutered male (finding)
C1319065|Castrated male (finding)
C1319065|Neutered
C1284842|Entire male (body structure)
C1284842|Entire male
C0227926|Male genitourinary system
C0227926|Male genitourinary system structure (body structure)
C0227926|Male genitourinary system structure
C0227926|Male genitourinary tract
C0227926|Male genitourinary system, NOS
C0227926|Male genitourinary tract, NOS
C0242664|Husband
C0242664|Husband (person)
C0242664|Husbands
C0870831|Male Criminals
C1706429|Male
C1706429|Male, Self-Reported
C1706429|Male, Self-Report
C1706429|Male Sex, Self Report
C1706428|Male
C1706428|Male Phenotype
C1706180|Male
C1706180|Male Gender, Self Reported
C1706180|Male Gender, Self Report
C1706180|Male Gender
C0729953|Male genital vein
C0729953|Male genital vein (body structure)
C0419384|Male baby
C0419384|Baby male
C0419384|Baby male (finding)
C0574034|Spermatic cord and male perineal structures
C0574034|Spermatic cord and/or male perineal structures (body structure)
C0574034|Spermatic cord and/or male perineal structures
C0574034|Spermatic cord and male perineal structures (body structure)
C0447084|Artery of male pelvic region
C0447084|Artery of male pelvic region (body structure)
C1276151|Lymphatics of male pelvis
C1276151|Structure of lymphatic vessel of male pelvis (body structure)
C1276151|Structure of lymphatic vessel of male pelvis
C1276151|Lymphatics of male pelvis (body structure)
C0015780|Female
C0015780|F
C0015780|Female Gender, Self Reported
C0015780|Female Gender, Self Report
C0015780|Female Gender
C0015780|Female Gender [Disease/Finding]
C0015780|Female (finding)
C0015780|Females
C0015780|Female individual
C0015780|Female structure (body structure)
C0015780|Female structure
C0015780|Female individual, NOS
C0015780|Female, NOS
C1561593|Undifferentiated
C1561593|Administrative Gender - Undifferentiated
C0036866|Characteristic, Sex
C0036866|Characteristics, Sex
C0036866|Difference, Sex
C0036866|Differences, Sex
C0036866|Dimorphism, Sex
C0036866|Dimorphisms, Sex
C0036866|Sex Characteristic
C0036866|Sex Characteristics
C0036866|Sex Difference
C0036866|Sex Dimorphisms
C0036866|sexual dimorphism (noncellular)
C0036866|gender difference
C0036866|Sex differences
C0036866|Sex Dimorphism
C0036866|Gender Differences
C0079399|Gender
C0079399|Gender [Disease/Finding]
C0079399|Gender (finding)
C0079399|Gender (observable entity)
C1522384|Sex
C1522384|Sex of individual
C1522384|Gender
C1522384|Sex structure (body structure)
C1522384|Sex structure
C1522384|Sex of individual, NOS
C1522384|Sex, NOS
C1257955|Genotypic Sex
C1257955|Sex, Genotypic
C1257956|Phenotypic Sex
C1257956|Sex, Phenotypic
C0278457|Indeterminate sex, unspecified
C0278457|Indeterminate sex
C0278457|indeterminate sex (diagnosis)
C0278457|Indeterminate sex NOS
C0278457|Indeterminate sex NOS (disorder)
C0278457|Indeterminate sex (finding)
C0278457|Indeterminate sex (body structure)
C0278457|sex; indeterminate
