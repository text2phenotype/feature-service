C0040615|Antipsychotic Agents
C4048284|Benzodiazepine
C0005064|Benzodiazepines
C0023870|Lithium
C3540800|Lithium antipsychotics
C0287163|Seroquel
C0072953|raclopride
C0072953|Benzamide, 3,5-dichloro-N-((1-ethyl-2-pyrrolidinyl)-methyl)-2-hydroxy-6-methoxy-
C0072953|Raclopride [Chemical/Ingredient]
C0073393|risperidone
C0073393|4H-Pyrido(1,2-a)pyrimidin-4-one, 3-(2-(4-(6-fluoro-1,2-benzisoxazol-3-yl)-1-piperidinyl)ethyl)-6 ,7,8,9-tetrahydro-2-methyl-
C0073393|risperidone (medication)
C0073393|Risperidone [Chemical/Ingredient]
C0073393|Risperidone (product)
C0073393|Risperidone (substance)
C0008286|Chlorpromazine
C0008286|10H-Phenothiazine-10-propanamine, 2-chloro-N,N-dimethyl-
C0008286|2-Chloro-10-(3-(dimethylamino)propyl)phenothiazine
C0008286|chlorpromazines (medication)
C0008286|chlorpromazines
C0008286|Chlorpromazine [Chemical/Ingredient]
C0008286|CPZ - Chlorpromazine
C0008286|Chlorpromazine (product)
C0008286|Chlorpromazine (substance)
C0016368|Fluphenazine
C0016368|1-Piperazineethanol, 4-(3-(2-(trifluoromethyl)-10H-phenothiazin-10-yl)propyl)-
C0016368|1-Piperazineethanol, 4-(3-(2-(trifluoromethyl)-10H-phenothiazin-10-yl)propyl)-(9CI)
C0016368|Fluphenazine [Chemical/Ingredient]
C0016368|Flufenazin
C0016368|Fluphenazine (product)
C0016368|Fluphenazine (substance)
C0018546|Haloperidol
C0018546|1-Butanone, 4-(4-(4-chlorophenyl)-4-hydroxy-1-piperidinyl)-1-(4-fluorophenyl)-
C0018546|4-[4-(4-Chlorophenyl)-4-hydroxy-1-piperidinyl]-1-(4-fluorophenyl)-1-butanone
C0018546|haloperidol (medication)
C0018546|Haloperidol [Chemical/Ingredient]
C0018546|Haloperidol [antipsychotic]
C0018546|Haloperidol [tics, chorea] [see D47..]
C0018546|Haloperidol [tics, chorea] [see D47..] (product)
C0018546|Haloperidol [antipsychotic] (product)
C0018546|Haloperidol (product)
C0018546|Haloperidol (substance)
C0018546|Haloperidol [antipsychotic] (substance)
C0018546|Haloperidol [tics, chorea] [see D47..] (substance)
C0031935|Pimozide
C0031935|2H-Benzimidazol-2-one, 1-(1-(4,4-bis(4-fluorophenyl)butyl)-4-piperidinyl)-1,3-dihydro-
C0031935|Opiran
C0031935|pimozide (medication)
C0031935|Pimozide [Chemical/Ingredient]
C0031935|Pimozide (product)
C0031935|Pimozide (substance)
C0033229|Prochlorperazine
C0033229|10H-Phenothiazine, 2-chloro-10-(3-(4-methyl-1-piperazinyl)propyl)-
C0033229|2-Chloro-10-(3-(1-methyl-4-piperazinyl)propyl)-phenothiazine
C0033229|prochlorperazine (medication)
C0033229|Prochlorperazine [Chemical/Ingredient]
C0033229|Prochlorperazine [nausea]
C0033229|Prochlorperazine [nausea] (product)
C0033229|Prochlorperazine [antipsych] [see dhe..]
C0033229|Prochlorperazine [antipsych] [see dhe..] (product)
C0033229|Prochlorperazine (product)
C0033229|Prochlorperazine (substance)
C0033229|PCPZ
C0033229|Prochlorperazine [antipsych] [see dhe..] (substance)
C0033229|Prochlorperazine [nausea] (substance)
C0039943|Thioridazine
C0039943|10H-Phenothiazine, 10-(2-(1-methyl-2-piperidinyl)ethyl)-2-(methylthio)-
C0039943|thioridazine (discontinued)
C0039943|thioridazine (discontinued) (medication)
C0039943|Thioridazine [Chemical/Ingredient]
C0039943|Thioridazine (product)
C0039943|Thioridazine (substance)
C0009079|Clozapine
C0009079|5H-Dibenzo(b,e)(1,4)diazepine, 8-chloro-11-(4-methyl-1-piperazinyl)-
C0009079|clozapine (medication)
C0009079|Clozapine [Chemical/Ingredient]
C0009079|8-Chloro-11-(4-methyl-1-piperazinyl)-5H-dibenzo(b,e)(1,4)diazepine
C0009079|Clozapine (product)
C0009079|Clozapine (substance)
C0016367|Flupenthixol
C0016367|1-Piperazineethanol, 4-(3-(2-(trifluoromethyl)-9H-thioxanthen-9-ylidene)propyl)-
C0016367|Flupentixol
C0016367|alpha-Flupenthixol
C0016367|Flupenthixol [Chemical/Ingredient]
C0016367|cis-Flupenthixol
C0016367|antipsychotics flupentixol
C0016367|Flupentixol (medication)
C0016367|Flupentixol [antipsychotic]
C0016367|Flupenthixol [antipsychotic] (product)
C0016367|Flupenthixol [antidepressant]
C0016367|Flupenthixol [antidepressant] (product)
C0016367|Flupenthixol [antipsychotic]
C0016367|Flupentixol [antidepressant]
C0016367|Flupentixol (product)
C0016367|Flupentixol (substance)
C0016367|Flupenthixol [antidepressant] (substance)
C0016367|Flupenthixol [antipsychotic] (substance)
C0026388|Molindone
C0026388|4H-Indol-4-one, 3-ethyl-1,5,6,7-tetrahydro-2-methyl-5-(4-morpholinylmethyl)-
C0026388|Molindone [Chemical/Ingredient]
C0026388|Molindone (product)
C0026388|Molindone (substance)
C0027999|Nialamide
C0027999|4-Pyridinecarboxylic acid, 2-(3-oxo-3-((phenylmethyl)amino)propyl)hydrazide
C0027999|1-(2-(Benzylcarbamoyl)ethyl)-2-isonicotinoylhydrazine
C0027999|Nialamide [Chemical/Ingredient]
C0027999|Nialamide (substance)
C0030815|Penfluridol
C0030815|4-Piperidinol, 1-(4,4-bis(4-fluorophenyl)butyl)-4-(4-chloro-3-(trifluoromethyl)phenyl)-
C0030815|Penfluridol [Chemical/Ingredient]
C0030815|Penfluridol (substance)
C0035179|Reserpine
C0035179|Yohimban-16-carboxylic acid, 11,17-dimethoxy-18-((3,4,5-trimethoxybenzoyl)oxy)-, methyl ester, (3beta,16beta,17alpha,18beta,20alpha)-
C0035179|(3beta,16beta,17alpha,18beta,20alpha)-11,17-Dimethoxy-18-[(3,4,5-trimethoxybenzoyl)oxy]yohimban-16-carboxylic Acid Methyl Ester
C0035179|reserpine (medication)
C0035179|Reserpine [Chemical/Ingredient]
C0035179|Reserpine - chemical
C0035179|Reserpine - chemical (substance)
C0035179|Reserpine (product)
C0035179|Reserpine (substance)
C0037956|Spiperone
C0037956|1,3,8-Triazaspiro(4.5)decan-4-one, 8-(4-(4-fluorophenyl)-4-oxobutyl)-1-phenyl-
C0037956|Spiroperidol
C0037956|Spiperone [Chemical/Ingredient]
C0037956|Spiroperone
C0037956|Spiperone - chemical (substance)
C0037956|Spiperone - chemical
C0037956|Spiperone (substance)
C0038803|Sulpiride
C0038803|Benzamide, 5-(aminosulfonyl)-N-((1-ethyl-2-pyrrolidinyl)methyl)-2-methoxy-
C0038803|Sulpiride [Chemical/Ingredient]
C0038803|Sulperide
C0038803|N-((1-Ethyl-2-Pyrrolidinyl)Methyl)-5-Sulfamoyl-O-Anisamide
C0038803|antidepressants sulpiride
C0038803|sulpiride (medication)
C0038803|Sulpiride (product)
C0038803|Sulpiride (substance)
C0039955|Thiothixene
C0039955|9H-Thioxanthene-2-sulfonamide, N,N-dimethyl-9-(3-(4-methyl-1-piperazinyl)propylidene)-
C0039955|Thioxanthene-2-sulfonamide, N,N-dimethyl-9-(3-(4-methyl-1-piperazinyl)propylidene)-
C0039955|N,N-Dimethyl-9-(3-(4-methylpiperazin-1-yl)propylidene)-9H-thioxanthene-2-sulphonamide
C0039955|Navaron
C0039955|Orbinamon
C0039955|thiothixene (medication)
C0039955|Thiothixene [Chemical/Ingredient]
C0039955|Tiotixene
C0039955|Thiothixene (product)
C0039955|Thiothixene (substance)
C0040979|Trifluoperazine
C0040979|10H-Phenothiazine, 10-(3-(4-methyl-1-piperazinyl)propyl)-2-(trifluoromethyl)-
C0040979|10-(3-(4-Methyl-1-piperazinyl)propyl)-2-(trifluoromethyl)-10H-phenothiazine
C0040979|TFP
C0040979|Trifluoperazine [Chemical/Ingredient]
C0040979|Trifluoroperazine
C0040979|Trifluperazine
C0040979|Trifluoperazine [antipsychotic]
C0040979|Trifluoperazine [antipsychotic] (product)
C0040979|Trifluoperazine [nausea] [see dh4..] (product)
C0040979|Trifluoperazine [nausea] [see dh4..]
C0040979|10-[3-(4-Methyl-1-piperazinyl)propyl]-2-(trifluoromethyl)-10H-phenothiazine
C0040979|Trifluoperazine (product)
C0040979|Trifluoperazine (substance)
C0040979|Trifluoperazine [antipsychotic] (substance)
C0040979|Trifluoperazine [nausea] [see dh4..] (substance)
C0871650|Antischizophrenic Drugs
C0701357|ICI204636
C0701357|204636, ICI
C0701357|204,636, ICI
C0701357|ICI 204,636
C0701357|ICI-204636
C0701357|ICI 204636
C0171023|2-methyl-4-(4-methyl-1-piperazinyl)-10H-thieno(2,3-b)(1,5)benzodiazepine
C0171023|olanzapine
C0171023|olanzapine (medication)
C0171023|olanzapine [Chemical/Ingredient]
C0171023|olanzapine (Zyprexa)
C0171023|Olanzapine (product)
C0171023|Olanzapine (substance)
C0380393|5-(2-(4-(3-benzisothiazolyl)piperazinyl)ethyl)-6-chloro-1,3-dihydro-2H-indol-2-one
C0380393|ziprasidone
C0380393|2H-Indol-2-one, 5-(2-(4-(1,2-benzisothiazol-3-yl)-1-piperazinyl)ethyl)-6-chloro-1,3-dihydro-
C0380393|ziprasidone [Chemical/Ingredient]
C0380393|ziprazidone
C0380393|Ziprasidone (product)
C0380393|Ziprasidone (substance)
C0597883|alentemol
C0597884|antischizophrenic
C0000959|Acepromazine
C0000959|Ethanone, 1-(10-(3-(dimethylamino)propyl)-10H-phenothiazin-2-yl)-
C0000959|Acepromazine [Chemical/Ingredient]
C0000959|Acetopromazine
C0000959|Acetazine
C0000959|Acetylpromazine
C0000959|10-(3-Dimethylaminopropyl)phenothiazine-3-ethylone
C0000959|Acepromazine (substance)
C0004477|Azaperone
C0004477|1-Butanone, 1-(4-fluorophenyl)-4-(4-(2-pyridinyl)-1-piperazinyl)-
C0004477|Azaperone [Chemical/Ingredient]
C0004477|Azaperone (substance)
C0005013|Benperidol
C0005013|2H-Benzimidazol-2-one, 1-(1-(4-(4-fluorophenyl)-4-oxobutyl)-4-piperidinyl)-1,3-dihydro-
C0005013|benperidol (medication)
C0005013|Benperidol - chemical
C0005013|Benperidol (substance)
C0005013|Benperidol - chemical (substance)
C0005013|Benperidol [Chemical/Ingredient]
C0005013|Benperidol (product)
C0006467|Butaclamol
C0006467|Butaclamol [Chemical/Ingredient]
C0008290|Chlorprothixene
C0008290|1-Propanamine, 3-(2-chloro-9H-thioxanthen-9-ylidene)-N,N-dimethyl-, (Z)-
C0008290|chlorprothixene (medication)
C0008290|Chlorprotixen
C0008290|Chlorprothixene [Chemical/Ingredient]
C0008290|Chlorprothixene (product)
C0008290|Chlorprothixene (substance)
C0009026|Clopenthixol
C0009026|1-Piperazineethanol, 4-(3-(2-chloro-9H-thioxanthen-9-ylidene)propyl)-
C0009026|Clopenthixol (product)
C0009026|Clopenthixol [Chemical/Ingredient]
C0009026|Clopenthixol, Trans
C0009026|Clopenthixol (substance)
C0013136|Droperidol
C0013136|2H-Benzimidazol-2-one, 1-(1-(4-(4-fluorophenyl)-4-oxobutyl)-1,2,3,6-tetrahydro-4-pyridinyl)-1,3-dihydro-
C0013136|droperidol (medication)
C0013136|Droperidol [Chemical/Ingredient]
C0013136|Droperidol [central nervous system use] (product)
C0013136|Droperidol [central nervous system use]
C0013136|Droperidol [anesthesia] (product)
C0013136|Droperidol [anaesthesia]
C0013136|Droperidol [anesthesia]
C0013136|Droperidol (product)
C0013136|Droperidol (substance)
C0013136|Droperidol [anesthesia] (substance)
C0013136|Droperidol [central nervous system use] (substance)
C0014958|Etazolate
C0014958|1H-Pyrazolo(3,4-b)pyridine-5-carboxylic acid, 1-ethyl-4-((1-methylethylidene)hydrazino)-, ethyl ester
C0014958|Etazolate [Chemical/Ingredient]
C0016383|Fluspirilene
C0016383|1,3,8-Triazaspiro(4.5)decan-4-one, 8-(4,4-bis(4-fluorophenyl)butyl)-1-phenyl-
C0016383|Spirodiflamine
C0016383|Fluspirilene [Chemical/Ingredient]
C0016383|Fluspirilene (product)
C0016383|Fluspirilene (substance)
C0024056|Loxapine
C0024056|Dibenz(b,f)(1,4)oxazepine, 2-chloro-11-(4-methyl-1-piperazinyl)-
C0024056|loxapine (medication)
C0024056|Oxilapine
C0024056|2-Chloro-11-(4-methyl-1-piperazinyl)-dibenz(b,f)(1,4)oxazepine
C0024056|Cloxazepine
C0024056|Loxapine [Chemical/Ingredient]
C0024056|Loxapine (product)
C0024056|Loxapine (substance)
C0025497|Mesoridazine
C0025497|10H-Phenothiazine, 10-(2-(1-methyl-2-piperidinyl)ethyl)-2-(methylsulfinyl)-
C0025497|mesoridazine (medication)
C0025497|Mesoridazine [Chemical/Ingredient]
C0025497|Mesoridazine (product)
C0025497|Mesoridazine (substance)
C0025654|Methiothepin
C0025654|Piperazine, 1-(10,11-dihydro-8-(methylthio)dibenzo(b,f)thiepin-10-yl)-4-methyl-
C0025654|Metitepine
C0025654|Methiothepine
C0025654|Methiothepin [Chemical/Ingredient]
C0025678|Methotrimeprazine
C0025678|10H-Phenothiazine-10-propanamine, 2-methoxy-N,N,beta-trimethyl-, (R)-
C0025678|Methotrimeprazine product
C0025678|methotrimeprazine (discontinued) (medication)
C0025678|methotrimeprazine (discontinued)
C0025678|Levomepromazine
C0025678|Methotrimeprazine [Chemical/Ingredient]
C0025678|Levomeprazin
C0025678|Levopromazine
C0025678|(-)-10-(3-(Dimethylamino)-2-methylpropyl)-2-methoxyphenothiazine
C0025678|Levomepromazine product
C0025678|Methotrimeprazine product (substance)
C0025678|Levomeprazine
C0025678|Methotrimeprazine (product)
C0025678|Methotrimeprazine (substance)
C0025678|Levomepromazine product (substance)
C0030969|Perazine
C0030969|10H-Phenothiazine, 10-(3-(4-methyl-1-piperazinyl)propyl)-
C0030969|Perazine [Chemical/Ingredient]
C0030969|Pernazine
C0030969|Perazine (substance)
C0031184|Perphenazine
C0031184|1-Piperazineethanol, 4-(3-(2-chloro-10H-phenothiazin-10-yl)propyl)-
C0031184|4-[3-(2-Chloro-10H-phenothiazin-10-yl)propyl]-1-piperazineethanol
C0031184|perphenazine (medication)
C0031184|Chlorpiprazine
C0031184|Perphenazine [Chemical/Ingredient]
C0031184|Perfenazine
C0031184|Perphenazine [central nervous system use]
C0031184|Perphenazine [anesthesia]
C0031184|Perphenazine [central nervous system use] (product)
C0031184|Perphenazine [anesthesia] (product)
C0031184|Perphenazine [anaesthesia]
C0031184|Perphenazine (product)
C0031184|Perphenazine (substance)
C0031184|Perphenazine [anesthesia] (substance)
C0031184|Perphenazine [central nervous system use] (substance)
C0033399|Promazine
C0033399|10H-Phenothiazine-10-propanamine, N,N-dimethyl-
C0033399|Promazine [Chemical/Ingredient]
C0033399|Promazine (product)
C0033399|Promazine (substance)
C0040988|Trifluperidol
C0040988|1-Butanone, 1-(4-fluorophenyl)-4-(4-hydroxy-4-(3-(trifluoromethyl)phenyl)-1-piperidinyl)-
C0040988|Trifluridol
C0040988|Trifluperidol [Chemical/Ingredient]
C0040988|Trifluperidol (product)
C0040988|Trifluperidol (substance)
C0040989|Triflupromazine
C0040989|10H-Phenothiazine-10-propanamine, N,N-dimethyl-2-(trifluoromethyl)-
C0040989|triflupromazine (discontinued) (medication)
C0040989|triflupromazine (discontinued)
C0040989|Trifluopromazine
C0040989|Triflupromazine [Chemical/Ingredient]
C0040989|Fluopromazine
C0040989|Triflupromazine (product)
C0040989|Triflupromazine (substance)
C0085260|Ritanserin
C0085260|5H-Thiazolo(3,2-a)pyrimidin-5-one, 6-(2-(4-(bis(4-fluorophenyl)methylene)-1-piperidinyl)ethyl)-7-methyl-
C0085260|Ritanserin [Chemical/Ingredient]
C0085260|6-(2-(4-(Bis(4-fluorophenyl)methylene)-1-piperidinyl)ethyl)-7-methyl-5H-thiazolo(3,2-a)pyrimidin-5-one
C0085260|6-(2-(4-(Bis(P-Fluorophenyl)Methylene)-Piperidino)Ethyl)-7-Methyl-5h-Thiazolo-(3,2-A)Pyrimidin-5-One
C0061851|Ondansetron
C0061851|4H-Carbazol-4-one, 1,2,3,9-tetrahydro-9-methyl-3-((2-methyl-1H-imidazol-1-yl)methyl)-
C0061851|ondansetron (medication)
C0061851|Ondansetron [Chemical/Ingredient]
C0061851|Ondansetron, (+,-)-Isomer
C0061851|Ondansetron (product)
C0061851|Ondansetron (substance)
C0073047|Remoxipride
C0073047|Benzamide, 3-bromo-N-((1-ethyl-2-pyrrolidinyl)methyl)-2,6-dimethoxy-, (S)-
C0073047|Remoxipride [Chemical/Ingredient]
C0073047|(S)-3-Bromo-N-((1-ethyl-2-pyrrolidinyl)methyl)-2,6-dimethoxybenzamide
C0073047|Remoxipride (product)
C0073047|Remoxipride (substance)
C0023870|Lithium
C0023870|Lithium product
C0023870|lithium (medication)
C0023870|Lithium [Chemical/Ingredient]
C0023870|Lithium Metallicum
C0023870|Li
C0023870|Li element
C0023870|Li+ element
C0023870|Li - Lithium
C0023870|Lithium (product)
C0023870|Lithium (substance)
C0023870|Lithium, NOS
C0023870|Lithium product (product)
C0023870|Lithium product (substance)
C3179399|Hydrochloride, Tiapamil
C3179399|Tiapamil Hydrochloride
C3179399|Tiapamil Hydrochloride [Chemical/Ingredient]
C3179399|1,3-Dithiane-2-propanamine, 2-(3,4-dimethoxyphenyl)-N-(2-(3,4-dimethoxyphenyl)ethyl)-N-methyl-, 1,1,3,3-tetraoxide, hydrochloride
C3179399|N-(3,4-dimethoxyphenethyl)-2-(3,4-dimethoxyphenyl)-N-methyl-m-dithian-2-propylamin-1,1,3,3-tetroxide hydrochloride
C0040615|Agents, Antipsychotic
C0040615|Agents, Major Tranquilizing
C0040615|Agents, Major Tranquillizing
C0040615|Antipsychotic Agents
C0040615|Major Tranquilizing Agents
C0040615|Major Tranquillizing Agents
C0040615|antipsychotic agent
C0040615|Agents, Neuroleptic
C0040615|Drugs, Antipsychotic
C0040615|Drugs, Neuroleptic
C0040615|Tranquilizers, Major
C0040615|neuroleptic
C0040615|ANTIPSYCHOTICS
C0040615|Neuroleptic Agent
C0040615|Antischizophrenic Agent
C0040615|Major Tranquilizer
C0040615|neurological agents neuroleptics
C0040615|antipsychotics (medication)
C0040615|neuroleptics
C0040615|neuroleptics (medication)
C0040615|Antipsychotic Agent [TC]
C0040615|Antipsychotic
C0040615|[CN700] ANTIPSYCHOTICS
C0040615|Antipsychotic drug
C0040615|Antipsychotic drug (product)
C0040615|Antipsychotic drugs
C0040615|Neuroleptic Agents
C0040615|Major Tranquilizers
C0040615|Neuroleptic Drugs
C0040615|Tranquillizing Agents, Major
C0040615|Tranquilizing Agents, Major
C0040615|Neuroleptic drug
C0040615|Anti-psychotic agent (product)
C0040615|Anti-psychotic agent (substance)
C0040615|Anti-psychotic agent
C0040615|Anti-psychotic agent, NOS
C0040615|Neuroleptic drug, NOS
C0039623|Tetrabenazine
C0039623|2H-Benzo(a)quinolizin-2-one, 1,3,4,6,7,11b-hexahydro-9,10-dimethoxy-3-(2-methylpropyl)-
C0039623|Tetrabenazine Orphan Brand
C0039623|2-Oxo-3-isobutyl-9,10-dimethoxy-1,3,4,6,7,11-beta-hexahydro-
C0039623|Orphan Brand of Tetrabenazine
C0039623|Tetrabenazine [Chemical/Ingredient]
C0039623|neurological agents tetrabenazine
C0039623|tetrabenazine (medication)
C0039623|Tetrabenazine product
C0039623|Tetrabenazine (substance)
C0039623|Tetrabenazine product (product)
C0039623|Tetrabenazine product (substance)
C0304370|phenothiazine derivatives
C0304370|phenothiazine derivatives (medication)
C0304370|Phenothiazine derivative (substance)
C0304370|Phenothiazine derivative antipsychotic
C0304370|Phenothiazine derivative
C0304370|Phenothiazine derivative antipsychotic (product)
C0304370|Phenothiazine derivative antipsychotic agent (substance)
C0304370|Phenothiazine derivative antipsychotic agent
C0304370|Phenothiazine AND/OR derivative
C0304370|Phenothiazine AND/OR derivative (product)
C0304370|Phenothiazine derivative (product)
C0304370|Phenothiazine AND/OR derivative (substance)
C0304370|Phenothiazines
C0301410|Hydroxyphenamate
C0301410|2-hydroxy-2-phenylbutyl carbamate
C0301410|Hydroxyphenamate (substance)
C0301410|Oxyfenamate
C0165561|2-methyl-5-(4-methyl-1-piperazinyl)-11H-(1,2,4)triazolo(1,5-C)(1,3)benzodiazepine
C0165561|11H-(1,2,4)Triazolo(1,5-c)(1,3)benzodiazepine, 2-methyl-5-(4-methyl-1-piperazinyl)-
C0165561|batelapine
C2698335|Batelapine Maleate
C0054138|4-(4-(4-bromophenyl)-4-hydroxypiperidino)-4'-fluorobutyrophenone
C0054138|bromoperidol
C0054138|bromperidol
C0054138|bromperidol (medication)
C1321935|butaperazine maleate (medication)
C1321935|butaperazine maleate
C0133602|(2-(4-(6-fluoro-1,2-benzisoxazol-3-yl)-1-piperidinyl)ethyl)-2,9-dimethyl-4H-pyrido(1,2-a)pyrimidin-4-one
C0133602|ocaperidone
C0133602|4H-Pyrido(1,2-a)pyrimidin-4-one, 3-(2-(4-(6-fluoro-1,2-benzisoxazol-3-yl)-1-piperidinyl)ethyl)-2,9-dimethyl-
C2698647|Olanzapine Pamoate
C0137024|Benzamide, 3,5-dimethyl-N-(4-pyridinylmethyl)-
C0137024|N-(4-picolyl)-3,5-dimethylbenzamide
C0137024|picobenzide
C2699086|Rilapine
C0076043|2-trifluormethyl-6-fluoro-9-(3-(4-(2-hydroxypiperazin-1-yl))propyl)thioxanthene
C0076043|teflutixol
C2699912|Tenilapine
C0076666|tienocarbin
C0076666|tienocarbine
C0076685|10-fluoro-1,2,3,4,4a,5-hexahydro-3-methyl-7-(2-thienyl)pyrazino(1,2-a)(1,4)benzodiazepine
C0076685|timelotem
C2699946|Timirdine
C2699963|Tolpiprazole
C2700075|Triclodazol
C2699390|Cloxypendyl
C2698342|Belaperidone
C2698342|(+)-3-(2-((1S,5R,6S)-6-(p-Fluorophenyl)-3-azabicyclo(3.2.0)hept-3-yl)ethyl)-2,4(1H,3H)-quinazolinedione
C2699631|3,5-Dichlor-N-(2-(diethylamino)ethyl)-2-methoxybenzamid
C2699631|Diclometide
C2719618|Asenapine Maleate
C2719618|1H-Dibenz(2,3:6,7)oxepino(4,5-c)pyrrole, 5-chloro-2,3,3a,12b-tetrahydro-2-methyl-,(3aR,12bR)-rel-, (2Z)-2-butenedioate (1:1)
C2719618|5-chloro-2,3,3a,12b-tetrahydro-2-methyl-1H-dibenz(2,3-6,7)oxepino(4,5-c)pyrrole
C2699376|4-(2-Chloroxanthen-9-ylidene)-1-methylpiperidine
C2699376|Clopipazan
C0668910|carvotroline
C0668910|1H-Pyrido(4,3-b)indole, 8-fluoro-2,3,4,5-tetrahydro-2-(2-(4-pyridinyl)ethyl)-
C0770896|Thioproperazine Mesylate
C0770896|Thioproperazine Methanesulfonate
C0936105|Amitriptyline + perphenazine (product)
C0936105|Amitriptyline + perphenazine
C0936105|AMITRIPTYLINE/PERPHENAZINE
C0936105|amitriptyline-perphenazine
C0936105|amitriptyline, perphenazine drug combination
C0936105|amitriptyline - perphenazine
C0936105|amitriptyline-perphenazine combination
C0936105|Amitriptyline / Perphenazine
C0936105|perphenazine-amitriptyline combination
C0066682|fluphenazine enanthate
C0066682|Fluohenazine enanthate
C0066682|fluphenazine enanthate (discontinued) (medication)
C0066682|fluphenazine enanthate (discontinued)
C0066682|fluphenazine enanthate [Chemical/Ingredient]
C0066682|Fluphenazine enanthate (product)
C0066682|Fluphenazine enanthate (substance)
C0066682|Fluophenazine enanthate
C0066682|Fluophenazine enanthate (substance)
C0078168|veralipride
C0078168|N-(1-allyl-2-pyrrolidinyl)methyl-2,3-dimethoxy-5-sulfamoylbenzamide
C0078168|Veralipride (substance)
C0009071|clothiapine
C0009071|clotiapine
C0009071|Dibenzo(b,f)(1,4)thiazepine, 2-chloro-11-(4-methyl-1-piperazinyl)-
C0009071|clothiapine (medication)
C0009071|Clotiapine (substance)
C2000088|Asenapine
C2000088|Asenapine (product)
C2000088|Asenapine (substance)
C2000088|antipsychotics asenapine
C2000088|asenapine (medication)
C0951571|carpipramine dihydrochloride
C0050458|acetophenazine
C0050458|acetophenazine [Chemical/Ingredient]
C0050458|Acetophenazine (substance)
C2825691|Lorpiprazole
C0033459|Pericyazine
C0033459|Periciazine
C0033459|pericyazine (medication)
C0033459|propericiazine
C0033459|Pericyazine (product)
C0033459|Pericyazine (substance)
C2825692|Clopipazan Mesylate
C0060479|6,8-difluoro-2,3,4,9-tetrahydro-N,N-dimethyl-1H-carbazole-3-amine
C0060479|flucindole
C2825693|Fenimide
C0772014|prothipendyl hydrochloride
C2825694|Clothixamide Maleate
C2825695|Cyclophenazine Hydrochloride
C0068168|3-(3-hydroxyphenyl)-N-n-propylpiperidine
C0068168|3-PPP
C0068168|n-N-propyl-3(N-hydroxyphenyl)piperidine
C0068168|Phenol, 3-(1-propyl-3-piperidinyl)-
C0068168|Preclamol
C0068168|(-)-(S)-m-(1-Propyl-3-piperidyl)phenol
C0068168|n-N-propyl-3-(3-hydroxyphenyl)piperidine
C2827084|Benzindopyrine
C0247194|Ethanone, 1-(4-(3-(4-(6-fluoro-1,2-benzisoxazol-3-yl)-1-piperidinyl)propoxy)-3-methoxyphenyl)-
C0247194|iloperidone
C0247194|Iloperidone (substance)
C0247194|Iloperidone (product)
C0247194|4'-(3-(4-(6-Fluoro-1,2-benzisoxazol-3-yl)piperidino)propoxy)-3'-methoxyacetophenone
C0247194|antipsychotics iloperidone
C0247194|Iloperidone (medication)
C0072200|propionylpromazine
C0072200|propiopromazine
C0072200|1-Propanone, 1-(10-(3-(Dimethylamino)Propyl)-10H-Phenothiazin-2-yl)-
C0072200|1-Propanone, 1-(10-(3-(Dimethylamino)Propyl)Phenothiazin-2-yl)-
C0072200|1-(10-(3-(Dimethylamino)Propyl)-10H-Phenothiazin-2-yl)Propan-1-One
C0954036|Propiopromazine Hydrochloride
C0954036|1-(10-(3-(Dimethylamino)Propyl)-10H-Phenothiazin-2-yl)-1-Propanone
C0954036|1-Propanone, 1-(10-(3-(Dimethylamino)Propyl)-10H-Phenothiazin-2-yl)-, Monohydrochloride
C0954036|Propionylpromazine Hydrochloride
C0954036|Propiopromazine hydrochloride (substance)
C0139007|prothipendyl
C0139007|Prothipendyl (substance)
C0075591|sulforidazine
C2026712|ceruletide diethylamine (discontinued) (medication)
C2026712|neuroleptics ceruletide diethylamine (discontinued)
C2026712|ceruletide diethylamine (discontinued)
C2092061|traditional antipsychotics (medication)
C2092061|traditional antipsychotics
C2092062|novel antipsychotics
C2092062|novel antipsychotics (medication)
C1875654|PHENOTHIAZINE/RELATED ANTIPSYCHOTICS
C1875654|[CN701] PHENOTHIAZINE/RELATED ANTIPSYCHOTICS
C1874317|ANTIPSYCHOTICS,OTHER
C1874317|[CN709] ANTIPSYCHOTICS,OTHER
C2719626|paliperidone palmitate
C2719626|Hexadecanoic Acid, 3-(2-(4-(6-fluoro-1,2-benzisoxazol-3-yl)-1-piperidinyl)ethyl)-6,7,8,9-tetrahydro-2-methyl-4-oxo-4H-pyrido(1,2-a)pyrimidin-9-yl Ester
C2719626|Paliperidone palmitate (substance)
C2719626|Palmitate, Paliperidone
C2719626|Paliperidone Palmitate [Chemical/Ingredient]
C2719626|antipsychotics paliperidone palmitate
C2719626|paliperidone palmitate (medication)
C0031968|10H-Phenothiazine-2-sulfonamide,10-(3-(4-(2-hydroxyethyl)-1-piperidinyl)propyl)-N,N-dimethyl-
C0031968|pipothiazine
C0031968|pipotiazin
C0031968|Pipotiazine
C0031968|10-[3-[4-(2-Hydroxyethyl)Piperidino]Propyl]-N,N-Dimethylphenothiazine-2-Sulfonamide
C0031968|Pipothiazine (product)
C0031968|Pipotiazine (substance)
C0031968|Pipothiazine (substance)
C2983804|Cinuperone
C2983866|Lusaperidone
C0066451|2-methyl-11-(4-methyl-1-piperazinyl)-dibenzo (b,f)(1,4)thiazepine
C0066451|metiapine
C0069710|10-(3-(4-(2-(1,3-dioxan-2-yl)ethyl)-1- piperazinyl)propyl)-2-trifluoromethylphenothiazine
C0069710|oxaflumazine
C0533453|3-(3-(4--(5-methoxy-4-pyrimidinyl)-1-piperazinyl)propyl)-N-methyl-1H-indole-5-methanesulfonamide fumarate
C0533453|3-(3-(4-(5-Methoxy-4-pyrimidinyl)-1-piperazinyl)propyl)-N-methylindole-5-methanesulfonamide
C0533453|Avitriptan
C0006481|butaperazine
C0006481|butyrylperazine
C0006481|1-Butanone, 1-(10-(3-(4-methyl-1-piperazinyl)propyl)-10H-phenothiazin-2-yl)-
C0006481|Butaperizine
C0006481|Butaperazine (substance)
C2825448|Clothixamide
C2825448|Clotixamide
C0770895|pipothiazin palmitate
C0770895|pipothiazine palmitate
C0770895|Hexadecanoic acid, 2-(1-(3-(2-((dimethylamino)sulfonyl)-10H-phenothiazin-10-yl)propyl)-4-piperidinyl)ethyl ester
C0770895|pipotiazine palmitate
C0770895|pipotiazine palmitate (medication)
C0770895|10-(3-(4-(2-Hydroxyethyl)Piperidino)Propyl)-N,N-Dimethylphenothiazine-2-Sulfonamide Palmitate (Ester)
C0770895|Pipothiazine palmitate (product)
C0770895|Pipotiazine palmitate (substance)
C0770895|Pipothiazine palmitate (substance)
C0149491|clopenthixol acetate ester
C0149491|Zuclopenthixol acetate
C0149491|(Z)-4-[3-(2-chlorothioxanthen-9-ylidene)propyl]-1-piperazineethanol Acetate
C0149491|Zuclopenthixol acetate (product)
C0149491|Zuclopenthixol acetate (substance)
C0149492|Zuclopenthixol decanoate
C0149492|Decanoic acid, 2-(4-(3-(2-chloro-9H-thioxanthen-9-ylidene)propyl)-1-piperazinyl)ethyl ester, (Z)-
C0149492|Zuclopenthixol decanoate (product)
C0149492|Zuclopenthixol decanoate (substance)
C0149492|zuclopenthixole decanoate
C0350505|Zuclopenthixol dihydrochloride
C0350505|Zuclopenthixol dihydrochloride (substance)
C0350505|cis-Clopenthixol Hydrochloride
C0350505|(Z)-4-(3-(2-Chloro-9H-thioxanthen-9-ylidene)propyl)-1-piperazineethanol Dihydrochloride
C0350505|Zuclopenthixol Hydrochloride
C0350505|Zuclopenthixol dihydrochloride (product)
C0075662|6-(7-chloro-1,8-naphthyridin-2-yl)-2,3,6,7-tetrahydro-7-oxo-5H-(1,4)dithiino(2,3-c)pyrrol-5-yl-4-methylpiperazine-1-carboxylate
C0075662|suriclone
C0075662|(R,S)-6-(7-Chlor-1,8-naphthyridin-2-yl)-3,5,6,7-tetrahydro-5-oxo-2H-(1,4)dithixino(2,3-c)pyrrol-7-yl-4-methyl-1-piperazinylcarboxylat
C0075662|4-Methyl-1-piperazinecarboxylic acid ester with (+-)-6-(7-chloro-1,8-naphthyridin-2-yl)-2,3,6,7-tetrahydro-7-hydroxy-5H-p-dithiino(2,3-c)pyrrol-5-one
C0075662|(8-(7-chloro(1,8)naphthyridin-2-yl)-7-oxo-2,5-dithia-8-azabicyclo(4.3.0)non-10-en-9-yl) 4-methylpiperazine-1-carboxylate
C0006525|Butyrophenones
C0006525|butyrophenone
C0006525|butyrophenone (medication)
C0006525|Butyrophenones [Chemical/Ingredient]
C0006525|1-phenylbutan-1-one
C0006525|Butyrophenone product
C0006525|Butyrophenone (substance)
C0886927|Tiapride Hydrochloride
C0886927|Monohydrochloride, Tiapride
C0886927|Hydrochloride, Tiapride
C0886927|Tiapride Hydrochloride [Chemical/Ingredient]
C0886927|Tiapride Monohydrochloride
C0886927|N,N-Diethyl-2-((2-methoxy-5-(methylsulfonyl)benzoyl)amino)ethanaminium chloride
C2983907|Pentiapine Maleate
C0039961|Thioxanthenes
C0039961|Thioxanthenes [Chemical/Ingredient]
C0039961|Thioxanthene (product)
C0039961|Thioxanthene
C0039961|Thioxanthene (substance)
C0064748|4'-fluoro-4-(4-(p-fluorobenozyl)piperidino)butyrophenone
C0064748|lenperone
C0064748|Lenperone (substance)
C0175156|azacyclonol
C0175156|Diphenyl carbinol
C0175156|Azacyclonol (substance)
C0380392|Ziprasidone Hydrochloride
C0380392|5-(2-(4-(1,2-Benzisothiazol-3-yl)-1-piperazinyl)ethyl)-6-chloro-1,3-dihydro-2H-Indol-2-one Monohydrochloride
C0380392|ziprasidone hydrochloride (medication)
C0380392|antipsychotics ziprasidone hydrochloride
C0380392|Ziprasidone hydrochloride (substance)
C0608826|aceprometazine
C0608826|1-(10-(2-(dimethylamino)propyl)-10H-phenothiazin- 2-yl)ethanone
C0654391|4-(4-bromophenyl)-1-(4-(4-fluorophenyl)-4-oxobutyl)-4-piperidinyl decanoate
C0654391|bromperidol decanoate
C0654391|bromperidol decanoate (medication)
C1981574|Antipsychotics &#x7C; urine
C1994723|Pimozide &#x7C; bld-ser-plas
C0060157|2-ethylamino-3-phenylnorcamphane
C0060157|bicyclo(2.2.1)heptan-2-amine, N-ethyl-3-phenyl-
C0060157|fencamfamine
C0060157|N-ethyl-3-phenylbicyclo(2.2.1)heptan-2-amine
C0060157|Fencamfamin
C0060157|2-Norbornanamine, N-Ethyl-3-Phenyl-
C0060157|3-Phenyl-N-Ethyl-2-Norbornanamine
C0060157|2-Phenyl-3-Ethylaminobicyclo(2.2.1)Heptane
C0060157|2-Ethylamino-3-Phenylnorbornane
C0060157|Fencamfamin (substance)
C1974051|Sulpiride &#x7C; bld-ser-plas
C1981573|Antipsychotics &#x7C; bld-ser-plas
C1980662|Acetophenazine &#x7C; bld-ser-plas
C0043513|Zolazepam
C0043513|Pyrazolo(3,4-e)(1,4)diazepin-7(1H)-one, 4-(2-fluorophenyl)-6,8-dihydro-1,3,8-trimethyl-
C0043513|Zolazepam [Chemical/Ingredient]
C0043513|Zolasepam
C1981247|Amilsulpride &#x7C; bld-ser-plas
C0123091|quetiapine
C0123091|quetiapine (medication)
C0123091|2-(2-(4-dibenzo(b,f)(1,4)thiazepine-11-yl-1-piperazinyl)ethoxy)ethanol
C0123091|Quetiapine (product)
C0123091|Quetiapine (substance)
C0031436|Phenothiazines
C0031436|phenothiazines (medication)
C0031436|Phenothiazines [Chemical/Ingredient]
C1533126|Cyclopropanecarboxamide, 2-(aminomethyl)-N,N-diethyl-1-phenyl-, cis-(+-)-
C1533126|MILNACIPRAN
C1533126|Milnacipran (product)
C1533126|Milnacipran (substance)
C1533126|midalcipran
C1533126|milnacipran [Chemical/Ingredient]
C1533126|antidepressants snri milnacipran
C1533126|milnacipran (medication)
C2925168|Iloperidone &#x7C; Bld-Ser-Plas
C1994732|Pipamperone &#x7C; bld-ser-plas
C1983134|Bromperidol &#x7C; bld-ser-plas
C2925288|Methotrimeprazine metabolite &#x7C; Urine
C2738464|Norolanzapine &#x7C; Bld-Ser-Plas
C0770404|Carphenazine Maleate
C0770404|carphenazine maleate (discontinued) (medication)
C0770404|carphenazine maleate (discontinued)
C0770404|Carphenazine maleate (substance)
C3847696|Fluspirilene &#x7C; Bld-Ser-Plas
C3871108|Antipsychotics &#x7C; Blood or Urine
C0299792|aripiprazole
C0299792|2(1H)-Quinolinone, 7-(4-(4-(2,3-Dichlorophenyl)-1-piperazinyl)butoxy)-3,4-dihydro-
C0299792|aripiprazole (medication)
C0299792|7-(4-(4-(2,3-dichlorophenyl)-1-piperazinyl)butyloxy)-3,4-dihydro-2(1H)-quinolinone
C0299792|Aripiprazole [Chemical/Ingredient]
C0299792|Aripiprazol
C0299792|Aripiprazole (product)
C0299792|Aripiprazole (substance)
C4038379|7-Hydroxyquetiapine &#x7C; Urine
C0724680|Quetiapine Fumarate
C0724680|Ethanol, 2-(2-(4-dibenzo(b,f)(1,4)thiazepin-11-yl-1-piperazinyl)ethoxy)-,(E)-2-butenedioate(2:1)(salt)
C0724680|Fumarate, Quetiapine
C0724680|Ethanol, 2-(2-(4-dibenzo(b,f)(1,4)thiazepin-11-yl-1-piperazinyl)ethoxy)-, (E)-2-butenedioate (2:1) (salt)
C0724680|Quetiapine Fumarate [Chemical/Ingredient]
C0724680|Quetiapine fumarate (substance)
C2697950|Lurasidone Hydrochloride
C2697950|Lurasidone hydrochloride (substance)
C2697950|HCl, Lurasidone
C2697950|Hydrochloride, Lurasidone
C2697950|Lurasidone HCl
C2697950|Lurasidone Hydrochloride [Chemical/Ingredient]
C4072501|Benperidol &#x7C; Bld-Ser-Plas
C0103045|Amisulpride
C0103045|Amisulpride - chemical
C0103045|Amisulpride (substance)
C0103045|Amisulpride - chemical (substance)
C0103045|Amisulpride (product)
C4072058|Penfluridol &#x7C; Bld-Ser-Plas
C2003424|Lurasidone
C2003424|N-(2-(4-(1,2-benzisothiazol-3-yl)-1-piperazinylmethyl)-1-cyclohexylmethyl)-2,3-bicyclo(2.2.1)heptanedicarboximide
C2003424|Lurasidone (substance)
C2003424|lurasidone (medication)
C2003424|antipsychotics lurasidone
C4056439|aripiprazole lauroxil
C4056439|antipsychotics aripiprazole lauroxil
C4056439|aripiprazole lauroxil (medication)
C0358425|Anxiolytics and neuroleptic perioperative drugs (product)
C0358425|Anxiolytics and neuroleptic perioperative drugs
C0358425|Anxiolytics and neuroleptic perioperative drugs (substance)
C0030077|oxypertine
C0030077|1H-Indole, 5,6-dimethoxy-2-methyl-3-(2-(4-phenyl-1-piperazinyl)ethyl)-
C0030077|5,6-Dimethoxy-2-Methyl-3-(2-(4-Phenyl-1-Piperazinyl)Ethyl)Indole
C0030077|Win 18,501-2
C0030077|Oxypertine (product)
C0030077|Oxypertine (substance)
C0355185|Antipsychotic depot injections (product)
C0355185|Antipsychotic depot injections
C0355185|Antipsychotic depot injections (substance)
C0304387|Butyrophenone derivative antipsychotic agent (product)
C0304387|Butyrophenone derivative antipsychotic agent (substance)
C0304387|Butyrophenone derivative antipsychotic agent
C0304387|Butyrophenone derivative antipsychotic agent, NOS
C0304389|Dibenzoxazepine derivative antipsychotic agent (product)
C0304389|Dibenzoxazepine derivative antipsychotic agent (substance)
C0304389|Dibenzoxazepine derivative antipsychotic agent
C0304389|Dibenzoxazepine derivative antipsychotic agent, NOS
C0304392|Dihydroindolone derivative antipsychotic agent (product)
C0304392|Dihydroindolone derivative antipsychotic agent (substance)
C0304392|Dihydroindolone derivative antipsychotic agent
C0304392|Dihydroindolone derivative antipsychotic agent, NOS
C0304393|Diphenylbutylpiperidine derivative antipsychotic agent (product)
C0304393|Diphenylbutylpiperidine derivative antipsychotic agent (substance)
C0304393|Diphenylbutylpiperidine derivative antipsychotic agent
C0304393|Diphenylbutylpiperidine derivative antipsychotic agent, NOS
C1268911|Phenylbutylpiperadine derivative antipsychotic agent (product)
C1268911|Phenylbutylpiperadine derivative antipsychotic agent (substance)
C1268911|Phenylbutylpiperadine derivative antipsychotic agent
C1276996|Atypical antipsychotic
C1276996|Atypical antipsychotic (product)
C1276996|Atypical antipsychotic (substance)
C0304383|Thioxanthene derivative antipsychotic agent (product)
C0304383|Thioxanthene derivative antipsychotic agent (substance)
C0304383|Thioxanthene derivative antipsychotic agent
C0304383|Thioxanthene derivative antipsychotic agent, NOS
C1268910|Benzisoxazole derivative antipsychotic agent (product)
C1268910|Benzisoxazole derivative antipsychotic agent (substance)
C1268910|Benzisoxazole derivative antipsychotic agent
C1320173|Dihydrocarbostyril derivative antipsychotic (product)
C1320173|Dihydrocarbostyril derivative antipsychotic agent (substance)
C1320173|Dihydrocarbostyril derivative antipsychotic agent
C1320173|Dihydrocarbostyril derivative antipsychotic
C0100267|8-hydroxyloxapine
C0100267|Dibenz(b,f)(1,4)oxazepin-8-ol, 2-chloro-11-(4-methyl-1-piperazinyl)-
C0100267|8-hydroxyloxapine (substance)
C0304394|Dimozide
C0304394|Dimozide (substance)
C0753678|paliperidone
C0753678|Paliperidone (substance)
C0753678|Paliperidone (product)
C0753678|paliperidone (medication)
C0753678|9-Hydroxyrisperidone
C0753678|4H-Pyrido(1,2-a)pyrimidin-4-one, 3-(2-(4-(6-fluoro-1,2-benzisoxazol-3-yl)-1-piperidinyl)ethyl)-6,7,8,9-tetrahydro-9-hydroxy-2-methyl-
C0753678|9 Hydroxy risperidone
C0753678|9 OH risperidone
C0753678|9 Hydroxyrisperidone
C0753678|9-Hydroxy-risperidone
C0753678|3-(2-(4-(6-fluoro-3-(1,2-benzisoxazolyl))-1-piperidinyl)ethyl)-6,7,8,9-tetrahydro-9-hydroxy-2-methyl-4H-pyrido(1,2-a)pyrimidin-4-one
C0753678|9-OH-risperidone
C0753678|9-Hydroxyrisperidone (substance)
C0060473|4'-fluoro-4-(4-(o-methoxyphenyl)-1-piperazinyl)- butyrophenone
C0060473|fluanisone
C0060473|haloanisone
C0060473|haloanizone
C0071098|1'-(3-(4-fluorobenzoyl)propyl)-(1,4'-bipiperidine) -4'-carboxamide
C0071098|pipamperone
C0071098|Pipamperone (product)
C0071098|Pipamperone (substance)
C0066477|4'-fluor-4-(4-methylpiperidino)-butyrophenone
C0066477|melperon
C0066477|melperone
C0066477|methylperon
C0066477|metylperon
C0066477|Melperone (substance)
C0066477|Melperone (product)
C0075226|stepholidine
C0075630|N-(ethyl-1-pyrrolidinyl- 2-methyl)methoxy-2-ethylsulfonyl-5-benzamide
C0075630|sultopride
C0075630|N-((1-ethyl-2-pyrrolidinyl)methyl)-5-(ethylsulfonyl)-O-anisamide
C0074587|2,6-methano-3-benzazocin-8-ol, 1,2,3,4,5,6-hexahydro-6,11-dimethyl-3-(2-propenyl)-
C0074587|SK&F 10047
C0074587|SKF 10047
C0074587|SKF-10047
C0058518|10-(2-methyl 3-(1-hydroxyethoxyethyl-4-piperazinyl)propyl)phenothiazine
C0058518|dixyrazine
C0076278|5,8,13,13a-tetrahydro-2,3,9,10-tetramethoxy-6H-dibenzo(a,g)quinolizine
C0076278|tetrahydropalmatine
C0076278|tetrahydropalmitine
C0071053|6-fluoro-9-(3-(4-(2-hydroxyethyl)piperidino) propylidene)-2-trifluoromethyl-thioxanthene
C0071053|piflutixol
C0063970|1-Piperazineethanol, 4-(3-fluoro-10,11-dihydro-8-(1-methylethyl)dibenzo(b,f)thiepin-10-yl)-
C0063970|3-fluor-8-isopropyl-10-(4-(2-hydroxyethyl)piperazino)-10,11-dihydrodibenzo(b,f)thiepin
C0063970|isofloxythepin
C0078849|2-chloro-11-(2-dimethylaminoethoxy)dibenzo(b,f)thiepine
C0078849|zotepine
C0078849|2-((8-Chlorodibenzo(b,f)thiepin-10-yl)oxy)-N,N-dimethylethanamine
C0078849|Zotepine (product)
C0078849|Zotepine (substance)
C0076688|4'-fluoro-4-(4-(2-thioxo-1-benzimidazolinyl)piperidino)butyrophenone
C0076688|4-(4-(2,3-dihydro-2-thioxo-1H-benzimidazol-1-yl)-1-piperidinyl)-1-(4-fluorophenyl)-1- butanone
C0076688|timiperone
C0078761|1-(3-chlorophenyl)-3-(2-(3,3-dimethyl-1-azetidinyl)ethyl)imidazolidin-2-one
C0078761|2-Imidazolidinone, 1-(3-chlorophenyl)-3-(2-(3,3-dimethyl-1-azetidinyl)ethyl)-
C0078761|zetidoline
C0055929|clopenthixol decanoate
C0055929|clopentixol decanoate
C0058537|DN 1417
C0058537|DN-1417
C0058537|L-Prolinamide, N-((tetrahydro-5-oxo-2-furanyl)carbonyl)-L-histidyl-
C0217937|benzamide, 5-chloro-2-methoxy-4-(methylamino)-N-(2-methyl-1-(phenylmethyl)-3-pyrrolidinyl)-
C0217937|nemonapride
C0073502|4H-Pyrrolo(2,3-g)isoquinolin-4-one, 3-ethyl-1,4a,5,6,7,8,8a,9-octahydro-2,6-dimethyl-, trans-(+-)-
C0073502|Ro 22-1319
C0073502|Ro-22-1319
C0062103|haloperidol decanoate
C0062103|Haloperidol deconoate
C0062103|haloperidol decanoate (discontinued) (medication)
C0062103|haloperidol decanoate (discontinued)
C0062103|haloperidol decanoate [Chemical/Ingredient]
C0062103|Haloperidol decanoate (product)
C0062103|Haloperidol decanoate (substance)
C0062103|Haloperidol deconoate (substance)
C0140593|cis-9-(3-(3,5-dimethyl-1-piperazinyl)propyl)carbazole
C0140593|rimcazole
C0057143|1,2,4-Triazolo(4,3-a)pyridine, 5,6,7,8-tetrahydro-3-(2-(4-(2-methylphenyl)-1-piperazinyl)ethyl)-
C0057143|dapiprazole
C0057143|dapiprazole [Chemical/Ingredient]
C0057143|Dapiprazole (product)
C0057143|Dapiprazole (substance)
C0060579|3-fluoro-6-(4-methylpiperazinyl)-11H-dibenz(b,e)azepine
C0060579|fluperlapine
C0051747|amperozide
C1099053|Ecopipam
C1099053|5H-Benzo(d)naphth(2,1-b)azepin-12-ol, 11-chloro-6,6a,7,8,9,13b-hexahydro-7-methyl-, trans-(-)-
C0378456|3,4,4a,10b-tetrahydro-4-propyl-2H,5H-(1)benzopyrano(4,3-b)-1,4-oxazin-9-ol
C0378456|PBPO
C0378456|PBTO
C0084572|2-(4-(4-(1,2-benzisothiazol-3-yl)-1-piperazinyl)butyl)hexahydro-1H-isoindole-1,3-(2H)-dione
C0084572|Perospirone
C0084528|1-(2-(4-(5-chloro-1-(4-fluorophenyl)-1H-indol-3-yl)-1-piperidinyl)ethyl)-2-imidazolidinone
C0084528|sertindole
C0084528|sertindole (medication)
C0084528|sertindole [Chemical/Ingredient]
C0084528|Sertindole (product)
C0084528|Sertindole (substance)
C0526908|2-(3-(4-(4-fluorophenyl)-1-piperazinyl)propyl)-2H-naphth(1,8-cd)isothiazole 1,1-dioxide
C0526908|fananserin
C0526908|fananserine
C0211640|DuP-734
C0211640|Ethanone, 2-(1-(cyclopropylmethyl)-4-piperidinyl)-1-(4-fluorophenyl)-, hydrobromide
C0211640|DuP 734
C0248068|Benzeneethanamine, 4-methoxy-3-(2-phenylethoxy)-N,N-dipropyl-, hydrochloride
C0248068|N,N-dipropyl-2-(4-methoxy-3-(2-phenylethoxy)phenyl)ethylamine monohydrochloride
C0293258|SR 142801
C0293258|SR-142801
C0293258|SR142801
C0389977|3-((4-(4-chlorophenyl)piperazin-1-yl)methyl)-1H-pyrrolo(2,3-b)pyridine
C0389977|CPMPP-3
C0057820|2,3,4,4a,5,9b-hexahydro-2,8-dimethyl-1H-pyrido(4,3-b)indole
C0057820|carbidine
C0057820|dicarbine
C0057820|1H-Pyrido(4,3-b)indole, 2,3,4,4a,5,9b-hexahydro-2,8-dimethyl-
C1443761|Benzimidazolinone derivative antipsychotic preparation (product)
C1443761|Benzimidazolinone derivative antipsychotic preparation
C1443762|Benzimidazolinone derivative antipsychotic agent (substance)
C1443762|Benzimidazolinone derivative antipsychotic agent
C0031434|phenothiazine
C0031434|phenosan
C0031434|Phenothiazine (product)
C0031434|Thiodiphenylamine
C0031434|Phenothiazine (substance)
C0031434|Phenothiazine, NOS
C0060580|fluphenazine decanoate
C0060580|fluphenazine depot
C0060580|ftorphenazine decanoate
C0060580|Flufenazine Decanoate
C0060580|fluphenazine decanoate (medication)
C0060580|fluphenazine depot [Chemical/Ingredient]
C0060580|Fluophenazine decanoate
C0060580|Fluophenazine decanoate (substance)
C0060580|Fluphenazine decanoate (product)
C0060580|Fluphenazine decanoate (substance)
C0304386|Thiothixene Hydrochloride
C0304386|CP 12252-1
C0304386|9H-Thioxanthene-2-sulfonamide, N,N-dimethyl-9-(3-(4-methyl-1-piperazinyl)propylidene)-, Dihydrochloride, Dihydrate
C0304386|antipsychotics thiothixene hydrochloride
C0304386|thiothixene hydrochloride (medication)
C0304386|Thiothixene hydrochloride (substance)
C0304386|Tiotixene hydrochloride
C1170754|Ziprasidone Mesylate
C1170754|ziprasidone mesylate (medication)
C1170754|Ziprasidone mesylate (substance)
C0242518|Thiethylperazine Maleate
C0242518|Thiethylperazine Malate
C0242518|thiethylperazine malate (discontinued)
C0242518|thiethylperazine malate (discontinued) (medication)
C0242518|thiethylperazine maleate (medication)
C0242518|Thiethylperazine Malate [Chemical/Ingredient]
C0242518|10H-Phenothiazine, 2-(ethylthio)-10-(3-(4-methyl-1-piperazinyl)propyl)-, (Z)-2-butenedioate
C0242518|Thiethylperazine malate (substance)
C0242518|Thiethylperazine maleate (substance)
C0033473|propiomazine
C0033473|1-Propanone, 1-(10-(2-(dimethylamino)propyl)-10H-phenothiazin-2-yl)-
C0033473|Dropiomazine
C0033473|Propiomazine -RETIRED-
C0033473|propiomazine [Chemical/Ingredient]
C0033473|Propiomazine (product)
C0033473|Propiomazine (substance)
C1721449|bifeprunox
C1721449|1-(2-Oxo-benzoxazolin-7-yl)-4-(3-biphenyl)methylpiperazinemesylate
C0601644|Imiclopazine
C0601644|1-(2-(4-(3-(2-chloro-10H-phenothiazin-10-yl)propyl)-1-piperazinyl)ethyl)-3- methyl-2-imidazolidinone
C0601644|1-(2-(3-(2-chlorophenothiazin- 10-yl)propyl)-1-piperazinylethyl)-3-methyl-2- imidazolidinone
C0601644|chlorimiphenine
C1883076|Spiclomazine
C0125997|lithium citrate
C0125997|lithium citrate (medication)
C0125997|LITHIUM (AS CITRATE)
C0125997|lithium citrate [Chemical/Ingredient]
C0125997|Lithium citrate (product)
C0125997|Lithium citrate (substance)
C0024057|Loxapine Succinate
C0024057|Butanedioic Acid, compound with 2-Chloro-11-(4-methyl-1-piperazinyl)dibenz(b,f)(1,4)oxazepine(1:1)
C0024057|2-Chloro-11-(4-methyl-1-piperazinyl)dibenz(b,f)(1,4)oxazepine Succinate(1:1)
C0024057|Cloxazepin
C0024057|loxapine succinate (medication)
C0024057|Loxapinsuccinate
C0024057|Daxolin
C0024057|Succinate, Loxapine
C0024057|Loxapine Succinate [Chemical/Ingredient]
C0024057|Loxipine Succinate
C0024057|Oxilapine succinate
C0024057|Loxapine succinate (substance)
C1880734|Farampator
C1880823|Fluspiperone
C0065505|4'-((3-(4-(2-fluorophenyl)-1-piperazinyl)propyl)oxy)-3'-methoxyacetanilide
C0065505|mafoprazine
C0700543|Mesoridazine Besylate
C0700543|Mesoridazine benzenesulphonate
C0700543|Mesoridazine benzenesulfonate
C0700543|Mesoridazine besylate (substance)
C0301379|Mebutamate
C0301379|mebutamate (discontinued)
C0301379|mebutamate (discontinued) (medication)
C0301379|Mebutamate (substance)
C0013015|Domperidone
C0013015|2H-Benzimidazol-2-one, 5-chloro-1-(1-(3-(2,3-dihydro-2-oxo-1H-benzimidazol-1-yl)propyl)-4-piperidinyl)-1,3-dihydro-
C0013015|Domperidon
C0013015|Domperidone [Chemical/Ingredient]
C0013015|Domperidone(motility) [see chapter d for preparations] (product)
C0013015|Domperidone(motility) [see chapter d for preparations]
C0013015|Domperidone [nausea]
C0013015|Domperidone [nausea] (product)
C0013015|GI prokinetic motility agents domperidone (medication)
C0013015|GI prokinetic motility agents domperidone
C0013015|antinauseants domperidone (medication)
C0013015|antinauseants domperidone
C0013015|Domperidone (product)
C0013015|Domperidone (substance)
C0013015|Domperidone [nausea] (substance)
C0013015|Domperidone(motility) [see chapter d for preparations] (substance)
C1880846|Fosenazide
C0546875|Hydrochloride, Promazine
C0546875|Promazine Hydrochloride
C0546875|Starazin
C0546875|Talofen
C0546875|10-(3-(Dimethylamino)propyl)phenothiazine Monohydrochloride
C0546875|10H-Phenothiazine-10-propanamine, N,N-dimethyl-, Monohydrochloride
C0546875|promazine hydrochloride (discontinued) (medication)
C0546875|antipsychotics promazine hydrochloride (discontinued)
C0546875|promazine hydrochloride (discontinued)
C0546875|Promazine Hydrochloride [Chemical/Ingredient]
C0546875|Promazine hydrochloride (substance)
C0546875|Promazine hydrochloride [dup] (substance)
C0085217|Carbonate, Lithium
C0085217|Lithium Carbonate
C0085217|Carbonate, Dilithium
C0085217|Carbonic acid, dilithium salt
C0085217|lithium carbonate (medication)
C0085217|Lithium Carbonate [Chemical/Ingredient]
C0085217|Dilithium Carbonate
C0085217|Lithium carbonate preparation
C0085217|Lithium carbonate (product)
C0085217|Lithium carbonate (substance)
C0023044|Propiomazine Hydrochloride
C0023044|Propiomazine hydrochloride (substance)
C0066492|2-methylamino-4-N-methylpiperazino-5-thiomethyl-6-chloropyrimidine
C0066492|2-pyridinamine, 4-chloro-N-methyl-6-(4-methyl-1-piperazinyl)-5-(methylthio)-
C0066492|mezilamine
C0075006|8-(3-(4-fluorophenoxy)propyl)-1-phenyl-1,3,8-triazaspiro(4.5)decan-4-one
C0075006|spiramide
C0075006|8-(3-(4-Fluorophenoxy) propyl)-1-phenyl-1,3,8-triazaspiro(4, 5)decan-4-one
C0058805|(4-fluorophenyl)(1-(3-(2-(trifluoromethyl)-10H-phenothiazine-10-yl)propyl)-4-piperidinyl)methanone
C0058805|duoperone
C0304376|Triflupromazine Hydrochloride
C0304376|triflupromazine hydrochloride (discontinued) (medication)
C0304376|antipsychotics triflupromazine hydrochloride (discontinued)
C0304376|triflupromazine hydrochloride (discontinued)
C0304376|Triflupromazine hydrochloride (substance)
C0663536|Panamesine
C0663536|(5S)-5-((4-Hydroxy-4-(3,4-(methylenedioxy)phenyl)piperidino)methyl)-3-(p-methoxyphenyl)-2-oxazolidinone
C0282249|Hydrochloride, Molindone
C0282249|Molindone Hydrochloride
C0282249|4H-Indol-4-one, 3-ethyl-1,5,6,7-tetrahydro-2-methyl-5-(4-morpholinylmethyl)-, Monohydrochloride
C0282249|Lidone
C0282249|molindone hydrochloride (medication)
C0282249|Molindone Hydrochloride [Chemical/Ingredient]
C0282249|Molindone Monohydrochloride
C0282249|Monohydrochloride, Molindone
C0282249|Molindone hydrochloride (substance)
C0386741|4-amino-2-butoxy-5-chloro-N-(1-(1,3-dioxolan-2-ylmethyl)piperid-4-yl)benzamide
C0386741|dobupride
C0376160|Zuclopenthixol
C0376160|Zuclopenthixol (substance)
C0376160|Zuclopenthixol (product)
C0376160|Clopentixol cis-(Z)-
C0376160|(Z)-4-(3-(2-Chlorothioxanthen-9-ylidene)propyl)-1-piperazineethanol
C0376160|alpha-Clopenthixol
C0376160|alpha Clopenthixol
C1882247|Oxypendyl
C0355077|Chlorpromazine hydrochloride
C0355077|2-Chloro-10-(3-(dimethylamino)propyl)phenothiazine Monohydrochloride
C0355077|chlorpromazine hydrochloride (medication)
C0355077|Chlorpromazine Hydrochloride [Chemical/Ingredient]
C0355077|Hydrochloride, Chlorpromazine
C0355077|ChlorproMAZINE Hydrochloride (obsolete)
C0355077|Chlorpromazine hydrochloride [anesthesia]
C0355077|Chlorpromazine hydrochloride [anesthesia] (product)
C0355077|Chlorpromazine hydrochloride (product)
C0355077|Chlorpromazine hydrochloride [nausea] [see dh2..]
C0355077|Chlorpromazine hydrochloride [nausea] [see dh2..] (product)
C0355077|Chlorpromazine hydrochloride [anaesthesia]
C0355077|Chlorpromazine hydrochloride (substance)
C0355077|Chlorpromazine hydrochloride [anesthesia] (substance)
C0355077|Chlorpromazine hydrochloride [nausea] [see dh2..] (substance)
C0031954|piperacetazine
C0031954|1-(10-(3-(4-(2-hydroxyethyl)-1-piperidinyl)propyl)-10H-phenothiazin-2-yl)ethanone
C0031954|piperacetazine (discontinued)
C0031954|piperacetazine (discontinued) (medication)
C0031954|piperacetazine [Chemical/Ingredient]
C0031954|Piperacetazine (substance)
C0304378|Acetophenazine Maleate
C0304378|acetophenazine maleate (discontinued)
C0304378|acetophenazine maleate (discontinued) (medication)
C0304378|Acetophenazine maleate (substance)
C1880547|Erizepine
C1881437|Lofendazam
C0070425|1-(3-(2-methoxyphenothiazin-10-yl)-2-methylpropyl)-4-piperidinol
C0070425|perimetazine
C0304381|Trifluoperazine Hydrochloride
C0304381|Trifluoperazine Dihydrochloride
C0304381|10-(3-(4-Methyl-1-piperazinyl)propyl)-2-(trifluoromethyl)-10H-phenothiazine Dihydrochloride
C0304381|trifluoperazine hydrochloride (medication)
C0304381|antipsychotics trifluoperazine hydrochloride
C0304381|Trifluoperazine HCL
C0304381|Trifluoperazine hydrochloride (product)
C0304381|Trifluoperazine Hydrochloride [Chemical/Ingredient]
C0304381|Trifluoperazine hydrochloride (substance)
C0700499|Thioridazine Hydrochloride
C0700499|thioridazine hydrochloride (medication)
C0700499|antipsychotics thioridazine hydrochloride
C0700499|Thioridazine HCL
C0700499|Thioridazine Hydrochloride [Chemical/Ingredient]
C0700499|Thioridazine hydrochloride (substance)
C0700499|Thioridazine hydrochloride [dup] (substance)
C0700567|Hydrochloride, Fluphenazine
C0700567|Fluphenazine Hydrochloride
C0700567|fluphenazine hydrochloride (medication)
C0700567|Fluphenazine Hydrochloride [Chemical/Ingredient]
C0700567|Fluphenazine hydrochloride (substance)
C0700567|Fluphenazine hydrochloride [dup] (substance)
C0062101|halopemide
C0062101|N-(2-(4-(5-chloro-2-oxo-1-benzimidazolinyl)piperidino)ethyl)-p-fluorobenzamide
C1997166|Benzamide derivative antipsychotic agent (product)
C1997166|Benzamide derivative antipsychotic agent (substance)
C1997166|Benzamide derivative antipsychotic agent
C1997166|Benzamide antipsychotic
C0080138|SCH 23390
C0080138|SCH-23390
C0080138|SCH23390
C2348790|Tilozepine
C2348297|Dimeprozan
C2348661|Terbequinil
C0075494|2-((3-(2-chloroethyl)tetrahydro-2H-1,3,2-oxazaphosphorin-2-yl)amino)ethanol, methanesulfonate (ester), P-oxide
C0075494|3-(2-chloroethyl)-2-(2-mesyloxyethylamino)tetrahydro-2H-1,3,2-oxazaphosphorine 2-oxide
C0075494|cytimun
C0075494|sufosfamide
C2347049|Brazergoline
C2346736|Amicarbalide
C2347353|Nifursemizone
C0762225|Abaperidone
C0762225|7-(3-(4-(6-fluoro-1,2-benzisoxazol-3-yl)piperidin-1-yl)propoxy)-3-(hydroxymethyl)chromen-4-one
C2346888|Axamozide
C0052743|azabuperone
C0052743|azabutyrone
C2346967|Batoprazine
C0771221|Carphenazine
C0039936|thioproperazine
C0039936|10H-Phenothiazine-2-sulfonamide, N,N-dimethyl-10-(3-(4-methyl-1-piperazinyl)propyl)-
C1451709|Sonepiprazole
C1451709|isoChr-EtPip-PhSO2NH2
C1451709|4-(4-(2-(isochroman-1-yl)ethyl)piperazin-1-yl)benzenesulfonamide
C1451709|4-(4-(2-(3,4-dihydro-1H-2-benzopyran-1-yl)ethyl)-1-piperazinyl)benzenesulfonamide monomethanesulfonate
C2348431|Alpertine
C0256089|quinagolide
C0256089|dopamine agonists CV 205-502
C0256089|quinagolide (medication)
C0256089|N,N-diethyl-N'-(1,2,3,4,4a,5,10,10a-octahydro-6-hydroxy-1-propyl-3-benzo(g)quinolinyl)sulfamide, (3alpha,4aalpha,10abeta)-(+-)-isomer
C0256089|quinagolide, (3alpha,4aalpha,10abeta)-(+-)-isomer
C0256089|Quinagolide (product)
C0256089|Quinagolide (substance)
C2348812|Traboxopine
C0071968|3-piperidino-1,1-diphenylpropanol
C0071968|3-piperidinyl-1,1-diphenylpropan-1-ol
C0071968|alpha,alpha-diphenyl-1-piperidinepropanol
C0071968|pridinol
C0071968|ridinol
C2347680|Prinomide Tromethamine
C2346887|Avitriptan Fumarate
C2346887|1H-Indole-5-methanesulfonamide, 3-(3-(4-(5-methoxy-4-pyrimidinyl)-1-piperazinyl)propyl)-N-methyl-, (E)-2-butenedioate (1:1)
C2348400|Elopiprazole
C2346998|Benzindopyrine Hydrochloride
C2348601|Sulmepride
C2347211|Broclepride
C2346718|Acaprazine
C0115127|Duoperone Fumarate
C2347032|Bisorcic
C2346745|Amiperone
C2346894|Azaquinzole
C2346785|Anisopirol
C0002333|Alprazolam
C0002333|4H-(1,2,4)Triazolo(4,3-a)(1,4)benzodiazepine, 8-chloro-1-methyl-6-phenyl-
C0002333|alprazolam (medication)
C0002333|Alprazolan
C0002333|Alprazolam [Chemical/Ingredient]
C0002333|Alprazolam - chemical
C0002333|Alprazolam - chemical (substance)
C0002333|Alprazolam (product)
C0002333|Alprazolam (substance)
C0008188|Chlordiazepoxide
C0008188|7 Chloro N methyl 5 phenyl 3H 1,4 benzodiazepin 2 amine 4 oxide
C0008188|3H-1,4-Benzodiazepin-2-amine, 7-chloro-N-methyl-5-phenyl-, 4-oxide
C0008188|3H-1,4-Benzodiazepin-2-amine, 7-chloro-N-methyl-5-phenyl, 4-oxide
C0008188|chlordiazepoxide (discontinued)
C0008188|chlordiazepoxide (discontinued) (medication)
C0008188|7-Chloro-N-methyl-5-phenyl-3H-1,4-benzodiazepin-2-amine 4-oxide
C0008188|Chlordiazepoxide [Chemical/Ingredient]
C0008188|Methaminodiazepoxide
C0008188|Chlordiazepoxide (product)
C0008188|Chlordiazepoxide (substance)
C0009011|Clonazepam
C0009011|2H-1,4-Benzodiazepin-2-one, 5-(2-chlorophenyl)-1,3-dihydro-7-nitro-
C0009011|clonazepam (medication)
C0009011|Clonazepam [Chemical/Ingredient]
C0009011|Clonazepam [status epilepsy]
C0009011|Clonazepam [status epilepsy] (product)
C0009011|Clonazepam [epilepsy control]
C0009011|Clonazepam [epilepsy control] (product)
C0009011|Clonazepam (product)
C0009011|Clonazepam (substance)
C0009011|Clonazepam [epilepsy control] (substance)
C0009011|Clonazepam [status epilepsy] (substance)
C0012010|Diazepam
C0012010|2H-1,4-Benzodiazepin-2-one, 7-chloro-1,3-dihydro-1-methyl-5-phenyl-
C0012010|7-Chloro-1,3-dihydro-1-methyl-5-phenyl-2H-1,4-benzodiazepin-2-one
C0012010|diazepam (medication)
C0012010|diazepam as anxiolytic (medication)
C0012010|diazepam as anxiolytic
C0012010|Diazepam [Chemical/Ingredient]
C0012010|Diazepam [anxiolytic]
C0012010|Diazepam [anesthesia]
C0012010|Diazepam [skeletal muscle relaxant] (product)
C0012010|Diazepam [anxiolytic] (product)
C0012010|Diazepam [epilepsy use] (product)
C0012010|Diazepam [epilepsy use]
C0012010|Diazepam [skeletal muscle relaxant]
C0012010|Diazepam [anaesthesia]
C0012010|Diazepam [anesthesia] (product)
C0012010|Diazepam product
C0012010|Diazepam (product)
C0012010|Diazepam (substance)
C0012010|Diazepam [anesthesia] (substance)
C0012010|Diazepam [anxiolytic] (substance)
C0012010|Diazepam [epilepsy use] (substance)
C0012010|Diazepam [skeletal muscle relaxant] (substance)
C0016375|Flurazepam
C0016375|2H-1,4-Benzodiazepin-2-one, 7-chloro-1-(2-(diethylamino)ethyl)-5-(2-fluorophenyl)-1,3-dihydro-
C0016375|Flurazepam [Chemical/Ingredient]
C0016375|7-Chloro-1-(2-(diethylamino)ethyl)-5-(2-fluorophenyl)-1,3-dihydro-2H-1,4-benzodiazepin-2-one
C0016375|Flurazepam (product)
C0016375|Flurazepam (substance)
C0024002|Lorazepam
C0024002|2H-1,4-Benzodiazepin-2-one, 7-chloro-5-(2-chlorophenyl)-1,3-dihydro-3-hydroxy-
C0024002|7-Chloro-5-(2-chlorophenyl)-1, 3-Dihydro-3-Hydroxy-1,4- Benzodiazepin-2-one
C0024002|lorazepam (medication)
C0024002|Lorazepam [Chemical/Ingredient]
C0024002|Lorazepam [epilepsy] (product)
C0024002|Lorazepam [anesthesia]
C0024002|Lorazepam [anesthesia] (product)
C0024002|Lorazepam [anxiolytic] (product)
C0024002|Lorazepam [anaesthesia]
C0024002|Lorazepam [epilepsy]
C0024002|Lorazepam [anxiolytic]
C0024002|Lorazepam (product)
C0024002|Lorazepam (substance)
C0024002|Lorazepam [anesthesia] (substance)
C0024002|Lorazepam [anxiolytic] (substance)
C0024002|Lorazepam [epilepsy] (substance)
C0026056|Midazolam
C0026056|4H-Imidazo(1,5-a)(1,4)benzodiazepine, 8-chloro-6-(2-fluorophenyl)-1-methyl-
C0026056|8-Chloro-6-(2-fluorophenyl)-1-Methyl- 4H- Imidazo(1,5a)(1,4)Benzodiazepine
C0026056|midazolam (medication)
C0026056|sedatives midazolam
C0026056|Midazolam [Chemical/Ingredient]
C0026056|Midazolam (product)
C0026056|Midazolam (substance)
C0029997|Oxazepam
C0029997|2H-1,4-Benzodiazepin-2-one, 7-chloro-1,3-dihydro-3-hydroxy-5-phenyl-
C0029997|Ro 5-6789
C0029997|Seresta
C0029997|oxazepam (medication)
C0029997|Oxazepam [Chemical/Ingredient]
C0029997|WY-3498
C0029997|Oxazepam (product)
C0029997|Oxazepam (substance)
C0040879|Triazolam
C0040879|4H-(1,2,4)Triazolo(4,3-a)(1,4)benzodiazepine, 8-chloro-6-(2-chlorophenyl)-1-methyl-
C0040879|clorazolam
C0040879|triazolam (medication)
C0040879|sedatives triazolam
C0040879|Triazolam [Chemical/Ingredient]
C0040879|8-Chloro-6-(2-chlorophenyl)-1-methyl-4H-(1,2,4)triazolo(4,3-a)(1,4)benzodiazepine
C0040879|Triazolam (product)
C0040879|Triazolam (substance)
C0055891|1-phenyl-5-methyl-8-chloro-1,2,4,5- tetrahydro-2,4-diketo-3H-1,5-benzodiazepine
C0055891|clobazam
C0055891|clobazam (medication)
C0055891|clobazam [Chemical/Ingredient]
C0055891|Clobazam [epilepsy only]
C0055891|Clobazam [epilepsy only] (product)
C0055891|Clobazam (product)
C0055891|Clobazam (substance)
C0055891|Clobazam [epilepsy only] (substance)
C0682884|short-acting benzodiazepines
C0682884|short-acting benzodiazepines (medication)
C0008174|clorazepate
C0008174|anxiolytics clorazepate
C0008174|clorazepate (medication)
C0008174|Clorazepate (substance)
C0008174|Clorazepate product (product)
C0008174|Clorazepate product
C0008174|Chlorazepate
C0917859|Hydrochloride, Zolazepam
C0917859|Zolazepam Hydrochloride
C0917859|Zolazepam hydrochloride (substance)
C0552500|Hydroxyalprazolam
C0552500|Hydroxyalprazolam (product)
C0552500|Hydroxyalprazolam (substance)
C0064304|11-chloro-8,12b-dihydro-2,8-dimethyl-12b-phenyl-4H-(1,3)oxazino(3,2-d)(1,4)benzodiazepine-4,7(6H)-dione
C0064304|ketazolam
C0064304|ketazolam (medication)
C0064304|Ketazolam (product)
C0064304|Ketazolam (substance)
C0006213|Bromazepam
C0006213|2H-1,4-Benzodiazepin-2-one, 7-bromo-1,3-dihydro-5-(2-pyridinyl)-
C0006213|bromazepam (medication)
C0006213|Bromazepam [Chemical/Ingredient]
C0006213|7-Bromo-1,3-Dihydro-5-(2-Pyridyl)-2H-1,4-Benzodiazepin-2-One
C0006213|Bromazepam - chemical
C0006213|Bromazepam - chemical (substance)
C0006213|Bromazepam (product)
C0006213|Bromazepam (substance)
C0065185|7-chloro-5-(2-chlorophenyl)-1,3-dihydro-3-hydroxy-1-methyl-2H-1,4-benzodiazepin-2-one
C0065185|lormetazepam
C0065185|sedatives lormetazepam
C0065185|lormetazepam (medication)
C0065185|7-Chloro-5-(O-Chlorophenyl)-1,3-Dihydro-3-Hydroxy-1-Methyl-2h-1,4-Benzodiazepin-2-One
C0065185|2H-1,4-Benzodiazepin-2-One, 7-Chloro-5-(2-Chlorophenyl)-1,3-Dihydro-3-Hydroxy-1-Methyl-
C0065185|Lormetazepam (product)
C0065185|Lormetazepam (substance)
C0072828|7-chloro-5-(2-fluorophenyl)-1,3-dihydro-1-(2,2,2-trifluoroethyl)-2H-1,4-benzodiazepine-2-thione
C0072828|quazepam
C0072828|2H-1,4-Benzodiazepine-2-thione, 7-chloro-5-(2-fluorophenyl)-1,3-dihydro-1-(2,2,2-trifluoroethyl)-
C0072828|quazepam (medication)
C0072828|quazepam [Chemical/Ingredient]
C0072828|Quazepam (substance)
C0072828|Quazepam product (product)
C0072828|Quazepam product
C0014892|Estazolam
C0014892|4H-(1,2,4)Triazolo(4,3-a)(1,4)benzodiazepine, 8-chloro-6-phenyl-
C0014892|8-Chloro-6-phenyl-4H-(1,2,4)triazolo-(4,3-a)(1,4)benzodiazepine
C0014892|sedatives estazolam
C0014892|estazolam (medication)
C0014892|Estazolam [Chemical/Ingredient]
C0014892|Estazolam (substance)
C0014892|Estazolam product (product)
C0014892|Estazolam product
C0011279|N Descyclopropylmethyl Prazepam
C0011279|N Descyclopropylmethylprazepam
C0011279|N Destrifluoroethylhalazepam
C0011279|Nordazepam
C0011279|2H-1,4-Benzodiazepin-2-one, 7-chloro-1,3-dihydro-5-phenyl-
C0011279|Desmethyldiazepam
C0011279|Demethyldiazepam
C0011279|N-Descyclopropylmethyl-Prazepam
C0011279|N-Descyclopropylmethylprazepam
C0011279|N-Destrifluoroethylhalazepam
C0011279|Nordazepam [Chemical/Ingredient]
C0011279|Deoxydemoxepam
C0011279|Nordiazepam
C0011279|Norprazepam
C0011279|7-Chloro-1,3-Dihydro-5-Phenyl-2H-1,4-Benzodiazepin-2-One
C0011279|Nordazepam (substance)
C0304401|Benzodiazepine nucleus
C0304401|Benzodiazepine nucleus (substance)
C0028126|Nitrazepam
C0028126|2H-1,4-Benzodiazepin-2-one, 1,3-dihydro-7-nitro-5-phenyl-
C0028126|nitrazepam (medication)
C0028126|sedatives nitrazepam
C0028126|Nitrazepam [Chemical/Ingredient]
C0028126|Nitrodiazepam
C0028126|1,3-Dihydro-7-Nitro-5-Phenyl-2H-1,4-Benzodiazepin-2-One
C0028126|Nitrazepam (product)
C0028126|Nitrazepam (substance)
C0525768|7-amino-flunitrazepam
C0525768|7-aminoflunitrazepam
C0525768|7-Aminoflunitrazepam (substance)
C0039468|Temazepam
C0039468|3 Hydroxydiazepam
C0039468|2H-1,4-Benzodiazepin-2-one, 7-chloro-1,3-dihydro-3-hydroxy-1-methyl-5-phenyl-
C0039468|Oxydiazepam
C0039468|10-chloro-4-hydroxy-6-methyl-2-phenyl-3,6-diazabicyclo[5.4.0]undeca-2,8,10,12-tetraen-5-one
C0039468|temazepam (medication)
C0039468|Hydroxydiazepam
C0039468|3-Hydroxydiazepam
C0039468|Temazepam [Chemical/Ingredient]
C0039468|Methyloxazepam
C0039468|Temazepam [anaesthesia]
C0039468|Temazepam [anesthesia] (product)
C0039468|Temazepam [anesthesia]
C0039468|Temazepam [hypnotic]
C0039468|Temazepam [hypnotic] (product)
C0039468|Temazepam (product)
C0039468|Temazepam (substance)
C0039468|Temazepam [anesthesia] (substance)
C0039468|Temazepam [hypnotic] (substance)
C0016296|Flunitrazepam
C0016296|2H-1,4-Benzodiazepin-2-one, 5-(2-fluorophenyl)-1,3-dihydro-1-methyl-7-nitro-
C0016296|flunitrazepam (medication)
C0016296|Fluridrazepam
C0016296|Flunitrazepam [Chemical/Ingredient]
C0016296|5-(O-Fluorophenyl)-1,3-Dihydro-1-Methyl-7-Nitro-2H-1,4-Benzodiazepin-2-One
C0016296|Flunitrazepam (product)
C0016296|Flunitrazepam (substance)
C1289963|Desmethylclobazam (substance)
C1289963|Desmethylclobazam
C0063132|hydroxyethylflurazepam
C0063132|Hydroxyethylflurazepam (substance)
C0077013|6-(2-chlorophenyl)-2,4-dihydro-2-((4-methyl-1-piperazinyl)methylene)-8-nitro-1H-imidazo(1,2-a) (1,4)benzodiazepin-1-one
C0077013|loprazolam
C0077013|triazulenone
C0077013|Loprazolam (product)
C0077013|Loprazolam (substance)
C0032910|Prazepam
C0032910|2H-1,4-Benzodiazepin-2-one, 7-chloro-1-(cyclopropylmethyl)-1,3-dihydro-5-phenyl-
C0032910|prazepam (discontinued) (medication)
C0032910|prazepam (discontinued)
C0032910|Prazepam [Chemical/Ingredient]
C0032910|Prazepam (product)
C0032910|Prazepam (substance)
C0025051|Medazepam
C0025051|1H-1,4-Benzodiazepine, 7-chloro-2,3-dihydro-1-methyl-5-phenyl-
C0025051|Medazapam
C0025051|Medazepam [Chemical/Ingredient]
C0025051|Medazapam (substance)
C0025051|Medazepam (product)
C0025051|Medazepam (substance)
C0062092|7-chloro-1,3-dihydro-5-phenyl-1- (2,2,2-trifluoroethyl)-2H-1,4-benzodiazepin-2-one
C0062092|halazepam
C0062092|halazepam (medication)
C0062092|halazepam [Chemical/Ingredient]
C0062092|Halazepam (substance)
C0062092|Halazepam product (product)
C0062092|Halazepam product
C0552501|Hydroxytriazolam
C0552501|Hydroxytriazolam (substance)
C0057377|7-chloro-1,3-dihydro-5-phenyl-2H-1,4-benzodiazepin-2-one 4-oxide
C0057377|demoxepam
C0057377|Demoxepam (substance)
C0690642|Triazolam 0.125 MG Oral Tablet
C0690642|Triazolam 0.125mg Oral tablet
C0690642|Triazolam, 0.125 mg oral tablet
C0690642|TRIAZOLAM 0.125MG TAB
C0690642|Triazolam 0.125 MILLIGRAM In 1 TABLET ORAL TABLET
C0690642|Triazolam Tab 0.125 MG
C0690642|TRIAZOLAM 0.125MG TAB [VA Product]
C0690642|TRIAZOLAM 0.125 mg ORAL TABLET [Triazolam]
C0690642|Triazolam 0.125mg tablet (product)
C0690642|Triazolam 0.125mg tablet
C0690643|Triazolam 0.25 MG Oral Tablet
C0690643|Triazolam 0.25mg Oral tablet
C0690643|Triazolam, 0.25 mg oral tablet
C0690643|TRIAZOLAM 0.25MG TAB
C0690643|Triazolam 0.25 MILLIGRAM In 1 TABLET ORAL TABLET
C0690643|Triazolam Tab 0.25 MG
C0690643|TRIAZOLAM 0.25MG TAB [VA Product]
C0690643|triazolam 0.25 mg ORAL TABLET [Triazolam]
C0690643|Triazolam 0.25mg tablet (product)
C0690643|Triazolam 0.25mg tablet
C4048284|benzodiazepine
C4048284|Benzodiazepine (product)
C4048284|Benzodiazepine (substance)
C4048284|Benzodiazepine, NOS
C0071082|7-chloro-5-phenyl-1-propargyl-1,4-benzodiazepin-2- one
C0071082|pinazepam
C0071082|propazepam
C0071082|Pinazepam (substance)
C0071082|Pinazepam (product)
C0009073|clotiazepam
C0009073|2H-Thieno(2,3-e)-1,4-diazepin-2-one, 5-(2-chlorophenyl)-7-ethyl-1,3-dihydro-1-methyl-
C0009073|Clotiazepam (substance)
C0053117|1,3,6,7,8,9-hexahydro-5-phenyl-2H-(1)benzothieno(2,3-e)-1,4-diazepin-2-one
C0053117|6,7-tetramethylene-5-phenyl-1,2-dihydro-3H-thieno(2,3-e)(1,4)diazepin-2-one
C0053117|bentazepam
C0053117|Bentazepam (substance)
C0076341|7-chloro-5-(1-cyclohexen-1- yl)-1,3-dihydro-1-methyl-2H-1,4-benzodiazepin-2-one
C0076341|tetrazepam
C0076341|tetrazepam (medication)
C0076341|Tetrazepam (substance)
C0054151|2-bromo-4-(2-chlorophenyl)-9-methyl-6H-thieno(3,2-f)(1,2,4)triazolo(4,3-a)(1,4)diazepine
C0054151|brotizolam
C0054151|sedatives brotizolam
C0054151|brotizolam (medication)
C0054151|6H-Thieno(3,2-F)(1,2,4)Triazolo(4,3-A)(1,4)Diazepine,2-Bromo-4-(2-Chlorophenyl)-9-Methyl-
C0054151|2-Bromo-4-(O-Chlorophenyl)-9-Methyl-6H-Thieno(3,2-F)-S-Triazolo(4,3-A)(1,4)Diazepine
C0054151|Brotizolam (substance)
C0005064|Benzodiazepines
C0005064|BENZODIAZEPINE CPDS
C0005064|benzodiazepines (medication)
C0005064|Benzodiazepines [Chemical/Ingredient]
C0005064|Benzodiazepine Compounds
C0005064|Benzodiazepine
C0360114|Benzodiazepine sedative
C0360114|Benzodiazepine sedative (product)
C0360114|Benzodiazepine sedative (substance)
C0053218|Benzodiazepine antiepileptic (product)
C0053218|Benzodiazepine antiepileptic
C0242293|Flurazepam Hydrochloride
C0242293|Hydrochloride, Flurazepam
C0242293|flurazepam hydrochloride (medication)
C0242293|Flurazepam Hydrochloride [Chemical/Ingredient]
C0242293|Flurazepam Dihydrochloride
C0242293|Dihydrochloride, Flurazepam
C0242293|Insumin Dihydrochloride
C0242293|Flurazepam HCl
C0242293|Flurazepam hydrochloride (substance)
C0057905|desalkylflurazepam
C0057905|desdialkylflurazepam
C0057905|dideethylflurazepam
C0057905|didesethylflurazepam
C0057905|N-desalkylflurazepam
C0057905|Desalkylflurazepam (substance)
C0057905|N-1-desalkylflurazepam
C0005065|Benzodiazepinones
C0005065|Benzodiazepinones [Chemical/Ingredient]
C0016293|Flumazenil
C0016293|4H-Imidazo(1,5-a)(1,4)benzodiazepine-3-carboxylic acid, 8-fluoro-5,6-dihydro-5-methyl-6-oxo-, ethyl ester
C0016293|flumazenil (medication)
C0016293|Flumazenil [Chemical/Ingredient]
C0016293|Flumazepil
C0016293|Flumazenil (product)
C0016293|Flumazenil (substance)
C0031978|Pirenzepine
C0031978|6H-Pyrido(2,3-b)(1,4)benzodiazepin-6-one, 5,11-dihydro-11-((4-methyl-1-piperazinyl)acetyl)-
C0031978|Pirenzepin
C0031978|Pyrenzepine
C0031978|Pirenzepine [Chemical/Ingredient]
C0031978|Pirenzepine (product)
C0031978|Pirenzepine (substance)
C0536095|Ro 48-6791
C0536095|Ro-48-6791
C0701356|WY 4036
C0701356|WY4036
C0701356|WY-4036
C0702213|Tazepam
C0702214|Serax
C0702215|Adumbran
C2352304|RS 678
C2352304|RS678 cpd
C2352304|RS-678
C2352305|RS 779
C2352305|RS779 cpd
C2352305|RS-779
C0009033|Chlorazepate, Dipotassium
C0009033|Clorazepate Dipotassium
C0009033|Dipotassium, Clorazepate
C0009033|1H-1,4-Benzodiazepine-3-carboxylic acid, 7-chloro-2,3-dihydro-2-oxo-5-phenyl-, monopotassium salt, compd. with potassium hydroxide (K(OH)) (1:1)
C0009033|1H-1,4-Benzodiazepine-3-carboxylic acid, 7-chloro-2,3-dihydro-2-oxo-5-phenyl-, Monopotassium Salt, compound with Potassium Hydroxide
C0009033|Potassium 7-chloro-2,3-dihydro-2-oxo-5-phenyl-1H-1,4-benzodiazepine-3-carboxylate KOH
C0009033|clorazepate dipotassium (medication)
C0009033|Clorazepate Dipotassium [Chemical/Ingredient]
C0009033|Dipotassium Chlorazepate
C0009033|Potassium clorazepate
C0009033|Clorazepate dipotassium (product)
C0009033|Clorazepate dipotassium (substance)
C0009033|Dipotassium clorazepate
C2604475|GWL78 cpd
C2604475|GWL 78
C2604475|GWL-78
C2604604|COCOBOO-acetamide
C2604604|2-(5-cyclohexyl-1-(2-cyclopentyl-2-oxoethyl)-2-oxo-1,2-dihydro-3H-1,3,4-benzotriazepin-3-yl)-N-(3-(5-oxo-2,5-dihydro-(1,2,4)oxadiazol-3-yl)phenyl)acetamide
C2604810|ethyl FNIBC
C2604810|ethyl 8-fluoro-6-(3-nitrophenyl)-4H-imidazo(1,5-a)(1,4)benzodiazepine-3-carboxylate
C2606964|PWZ-029
C2606902|quino(7,8-b)benzodiazepine
C0050844|adinazolam
C0167214|adinazolam mesylate
C0009034|Monopotassium, Clorazepate
C0009034|clorazepate monopotassium
C0009034|clorazepate monopotassium (medication)
C2699536|Cyprazepam
C2697918|Levotofisopam
C0068774|1-methyl-7-nitro-5-phenyl-1,3-dihydro-2H-1,4- benzodiazepin-2-one
C0068774|nimetazepam
C2698499|Nortetrazepam
C2699964|Tolufazepam
C2699964|1-(4'-Methylphenylsulfonyl)ethyl-5-(2-chlorophenyl)-7-chloro-2H-1,4-benzodiazepin-2-one
C2698992|Carburazepam
C0055715|8-bromo-6-(ortho-chlorophenyl)-1-cyclohexyl-4H-5-triazolo(3,4-c)thieno(2,4-e)-1,4-diazepine
C0055715|ciclotizolam
C0164835|7-chloro-5-(2-fluorophenyl)-2,3-dihydro-3-hydroxy-2-oxo-1H-1,4-benzodiazepine-1-propionitrile
C0164835|cinolazepam
C0110063|4H-Imidazo(1,5-a)(1,4)benzodiazepine, 8-chloro-6-(2-chlorophenyl)-1-methyl-
C0110063|8-chloro-6-(2-chlorophenyl)-1-methyl-4H-imidazo(1,5a)(1,4)benzodiazepine
C0110063|climazolam
C2714934|7-chloro-4-(cyclohexylmethyl)-1-methyl-3,4-dihydro-1H-1,4-benzodiazepine-2,5-dione
C2714934|BNZ-1 cpd
C2714935|4-cyclohexylmethyl-1-methyl-3,4-dihydro-1H-1,4-benzodiazepine-2,5-dione
C2714935|BNZ-2 cpd
C2715396|iodophenyl-MOPDBDU
C2715396|1-(3-iodophenyl)-3-(1-methyl-2-oxo-5-phenyl-2,3-dihydro-1H-benzo(e)(1,4)diazepin-3-yl)urea
C2715729|limazepine B1
C2715731|limazepine D
C2717477|RO4938581
C2717477|3-bromo-10-difluoromethyl-9H-imidazo(1,5-a)(1,2,4)triazolo(1,5-d)(1,4)benzodiazepine
C2744849|RO 4882224
C2744849|RO4882224
C2744849|RO-4882224
C0604102|7-chloro-2,3-dihydro-1-(2,2,2-trifluoroethyl)-5-(o-fluorophenyl)-1H-1,4-benzodia zepine
C0604102|fletazepam
C0065179|2H-pyrido(3,2-e)-1,4-diazepin-2-one, 7-chloro-5-(2-chlorophenyl)-1,3-dihydro-3-hydroxy-
C0065179|3-hydroxy-5-(o-chlorophenyl)-7-chloro-1,2-dihydro-2H-pyrido(3,2-e)-1,4-diazepin-2-one
C0065179|lopirazepam
C0089958|10-chloro-2,3,7,11b-tetrahydro-3-methyl-11b-(2-chlorophenyl)oxazolo(3,2-d)(1,4)benzodiazepin-6(5H)-one
C0089958|Mexazolam
C0089958|10-chloro-11b-(2-chlorophenyl)-2,3,7,11b-tetrahydro-3-methyloxazolo(3,2-d)(1,4)benzodiazepin-6(5H)-one
C0120735|10-bromo-11b-(2-fluorophenyl)-2,3,7,11b-tetrahydrooxazolo(3,2-d)(1,4)benzodiazepin-6(5H)-one
C0120735|haloxazolam
C0065842|3-methylclonazepam
C0065842|5-(2-chlorophenyl)-1,3-dihydro-3-methyl-7-nitro- 2H-1,4-benzodiazepin-2-one
C0065842|meclonazepam
C1619621|1H-1,4-Benzodiazepine, 7-bromo-5-(2-chlorophenyl)-2,3-dihydro-2-(methoxymethyl)-1-methyl-
C1619621|1H-1,4-Benzodiazepine, 7-bromo-5-(2-chlorophenyl)-2,3-dihydro-2-methoxy-1-methyl-
C1619621|metaclazepam
C0066040|Metaclazepam hydrochloride
C0066040|7-Bromo-5-(O-Chlorophenyl)-2,3-Dihydro-2-(Methoxymethyl)-1-Methyl-1H-1,4-Benzodiazepine Hydrochloride
C0066040|7-Bromo-5-(2-Chlorophenyl)-2,3-Dihydro-2-(Methoxymethyl)-1-Methyl-1H-1,4-Benzodiazepine Hydrochloride
C0066040|Brometazepam Hydrochloride
C0066040|Metuclazepam Hydrochloride
C0066040|7-bromo-5-(2'-chlorophenyl)-2,3-dihydro-2-(methoxyl)-1-methyl-1H-1,4-benzodiazepine.HCl
C0027556|Nefopam
C0027556|1H-2,5-Benzoxazocine, 3,4,5,6-tetrahydro-5-methyl-1-phenyl-
C0027556|Nefopam [Chemical/Ingredient]
C0027556|Benzoxazocine
C0027556|Nefopam (product)
C0027556|Nefopam (substance)
C0015820|Hydrochloride, Nefopam
C0015820|nefopam hydrochloride
C0015820|nefopam hydrochloride (medication)
C0015820|3,4,5,6-Tetrahydro-5-Methyl-1-Phenyl-1H-2,5-Benzoxazocine Hydrochloride
C0015820|Nefopam hydrochloride product (substance)
C0015820|Nefopam hydrochloride product
C0015820|Fenazoxine
C0015820|Nefopam hydrochloride (substance)
C0055964|10-chloro-2,3,5,6,7,11b-hexahydro-11b-(o- chlorophenyl)benzo(6,7)-1,4-diazepino-(5,4-b)-oxazol-6-one
C0055964|cloxazolam
C0055964|cloxazolam (medication)
C0055964|Betavel
C0055964|10-Chloro-11b-(o-chlorophenyl)-2,3,7,11b-tetrahydro-oxazolo(3,2-d) (1,4)benzodiazepin-6(5H)-one
C0055964|Enadel
C0055964|Tolestan
C0059772|1H-1,4-benzodiazepine-3-carboxylic acid, 7-chloro-5-(2-fluorophenyl)-2,3-dihydro-2-oxo-, ethyl ester
C0059772|ethyl flucozepate
C0059772|ethyl loflazepate
C0059772|ethyl loflazepate (medication)
C0059862|Etizolam
C0059862|etizolam (medication)
C2932012|4-(3,5-dihydroxybenzyl)-N-(2-methyl-4-((1-methyl-4,10-dihydropyrazolo(3,4-b)(1,5)benzodiazepin-5(1H)-yl)carbonyl)benzyl)piperazine-1-carboxamide
C2933864|EVT 201
C2933864|EVT201
C2933864|EVT-201
C2934398|2-amino-PPBI
C2934398|2-amino-4-(piperidin-1-yl)-11H-pyrimido(4,5-b)(1,5)benzodiazepin-6-ium
C2934400|2-amino-4-(methyl(2-methylphenyl)amino)-11H-pyrimido(4,5-b)(1,5)benzodiazepin-6-ium
C2934400|2-amino-MMAPBI
C2935069|benzopyrano(4,3-c)-1,5-benzodiazepine
C2935196|TKM0150
C2976597|5-(2-chlorophenyl)-7-fluoro-1,2-dihydro-8-methoxy-3-methylpyrazol(3,4b)(1,4)benzodiazepine
C1527794|Diazepinomicin
C1527794|11h-dibenzo(B,E)(1,4)diazepin-11-one, 5,10-dihydro-4,6,8-trihydroxy-10-((2E,6E)-3,7,11-trimethyl-2,6,10-dodecatrien-1-yl)-
C0117998|7-chloro-1-cyclopropylmethyl-1,3-dihydro-5-(2-fluorophenyl)-2H-1,4-benzodiazepin-2-one
C0117998|flutoprazepam
C1881907|Motrazepam
C1881907|2,3-Dihydro-1-(methoxymethyl)-7-nitro-5-phenyl-1H-1,4-benzodiazepin-2-on
C0605583|7-chloro-1,3-dihydro-5-phenyl-1H-2-oxo-3-pivalyloxy- 1,4-benzodiazepine
C0605583|pivoxazepam
C0605583|7-Chloro-1,3-dihydro-3-hydroxy-5-phenyl-2H-1,4-benzodiazepin-2-one Pivalate (Ester)
C2348591|Sulazepam
C0059029|7-chloro-1-(2-(ethylsulfonyl)ethyl)-5-(2-fluorophenyl)-1,3-dihydro-2H-1,4-benzodiazep in-2-one
C0059029|elfazepam
C2347902|Reclazepam
C2347902|2-(7-Chloro-5-(o-chlorophenyl)-2,3-dihydro-1H-1,4-benzodiazepin-1-yl)-2-oxazolin-4-one
C2347902|4(5H)-Oxazolone, 2-(7-chloro-5-(2-chlorophenyl)-2,3-dihydro-1H-1,4-benzodiazepin-1-yl)-
C3272985|3-(11-Dimethylheptyl)-7,8,9,10-tetrahydro-6,6,9-trimethyl-6H-dibenzo(b,d)pyran-1-yl 4-(1-azepanyl)butyrat
C3272985|1H-Azepine-1-butanoic acid, hexahydro-, 3-(1,2-dimethylheptyl)-7,8,9,10-tetrahydro-6,6,9-trimethyl-6H-dibenzo(b,d)pyran-1-yl ester
C3272985|SP 175
C3272985|Nabazenil
C3272985|SP-175
C0006795|camazepam
C0006795|Carbamic acid, dimethyl-, 7-chloro-2,3-dihydro-1-methyl-2-oxo-5-phenyl-1H-1,4-benzodiazepin-3-yl ester
C0006795|3-N,N-Dimethylcarbamoyloxy-7-chloro-5-phenyl-1-methyl-1,3-dihydro-2H-1,4-benzodiazepin-2-one
C0055353|2'-chloronordiazepam
C0055353|2H-1,4-Benzodiazepin-2-one, 7-chloro-5-(2-chlorophenyl)-1,3-dihydro-
C0055353|7-chloro-5-(2-chlorophenyl) 1,3-dihydro-2H-1,4-benzodiazepin-2-one
C0055353|chlordemethyldiazepam
C0055353|chlordesmethyldiazepam
C0055353|chlorodesmethyldiazepam
C0055353|Delorazepam
C0055353|2-Chloronordiazepam
C0055353|B1, Benzodiazepine
C0055353|Cl-DMDZ
C0055353|1,3-Dihydro-7-chloro-5-(o-chlorophenyl)-2H-1,4-benzodiazepin-2-one
C3273839|7-Chloro-1,3-dihydro-1-methyl-5-phenyl-2H-benzo-1,4-diazepin-2-onemonohydrochloride
C3273839|Diazepam Hydrochloride
C3273839|Diazepam HCl
C0887259|Monohydrochloride, Flurazepam
C0887259|Flurazepam Monohydrochloride
C0887259|2H-1,4-Benzodiazepin-2-one, 7-chloro-1-(2-(diethylamino)ethyl)-5-(2-fluorophenyl)-1,3-dihydro-, Monohydrochloride
C0060689|7-chloro-1-(dimethylphosphinmethyl)-5-phenyl-1,3- dihydro-2H-1,4-benzodiazepin-2-one
C0060689|fosazepam
C0060689|2H-1,4-Benzodiazepin-2-one, 7-chloro-1-((dimethylphosphinyl)methyl)-1,3-dihydro-5-phenyl-
C0060689|7-Chloro-1-((dimethylphosphinyl)methyl)-1,3-dihydro-5-phenyl-2H-1,4-benzodiazepin-2-one
C0172965|(1-hydrazinocarbonyl)-7-bromo-5-phenyl-1,2-dihydro-3H-1,4-benzodiazepine-2-one
C0172965|gidazepam
C0069747|butanedioic acid, mono(7-chloro-2,3-dihydro-2-oxo-5-phenyl-1H-1,4-benzodiazepin-3-yl) ester
C0069747|oxazepam hemisuccinate
C0069747|(RS)-Oxazepam H
C0069747|( -)-Oxazepam succinate
C0069747|7-Chloro-1,3-dihydro-3-hemisuccinyloxy-2H-1,4-benzodiazepin-2-one
C3273842|Oxazepam Monosodium Succinate
C0070543|7-bromo-5-(2-chlorphenyl)-1,2-dihydro-3H-1,4-benzodiazepin-2-one
C0070543|fenazepam
C0070543|phenazepam
C0070543|7-bromo-5-(2-chlorophenyl) 1,3-dihydro-2H-1,4-benzodiazepin-2-one
C0070543|2H-1,4-Benzodiazepin-2-one, 1,3-dihydro-7-bromo-5-(2-chlorophenyl)-
C0073389|1-ethyl-4,6-dihydro-3-methyl-8-phenylpyrazolo(4,3-e)(1,4)diazepin-5(lH)-one
C0073389|pyrazapon
C0073389|ripazepam
C0073389|1-Ethyl-4,6-dihydro-3-methyl-8-phenylpyrazolo(4,3-e)(1,4)diazepin-5(1H)-one
C0073389|Pyrazolo(4,3-e)(1,4)diazepin-5(1H)-one, 1-ethyl-4,6-dihydro-3-methyl-8-phenyl-
C3273843|Tuclazepam
C3273843|7-Chlor-5-(2-chlorphenyl)-2,3-dihydro-1-methyl-1H-1,4-benzodiazepin-2-methanol
C0077789|2-(allyloxy)amino 7-chloro-5-(o-chlorophenyl)-3H-1, 4-benzodiazepine
C0077789|uldazepam
C0077789|2-((Allyloxy)amino)-7-chloro-5-(o-chlorophenyl)-3H-1,4-benzodiazepine
C1982372|Benzodiazepines &#x7C; vitreous fluid
C1982367|Benzodiazepines &#x7C; gastric fluid
C1982371|Benzodiazepines &#x7C; urine
C1982364|Benzodiazepines &#x7C; bld-ser-plas
C1982365|Benzodiazepines &#x7C; body fluid
C2600781|Benzodiazepines.other &#x7C; Urine
C3534272|Benzodiazepines &#x7C; Saliva
C1972398|Quazepam &#x7C; bld-ser-plas
C1982369|Benzodiazepines &#x7C; meconium
C1982363|Benzodiazepine metabolites &#x7C; urine
C1982370|Benzodiazepines &#x7C; stool
C1982368|Benzodiazepines &#x7C; hair
C1982373|Benzodiazepines &#x7C; XXX
C3711897|R1498 compound
C3252279|evacetrapib
C3712514|olanzapine propan-2-ol hemisolvate monohydrate
C2975231|I-BET compound
C2975231|GSK525762A
C2975231|GSK 525762A
C2975231|GSK-525762A
C2975231|GSK525762
C2975231|IBET compound
C2975231|BET Inhibitor GSK525762
C2975231|I-BET762
C3713096|7-chloro-2-methylamino-5-phenyl-3H-1,4-benzodiazepine-4-oxide
C3712513|olanzapine propan-2-one hemisolvate monohydrate
C3491461|PF-184563
C3177676|7-methoxy-8-(5-(4-(1,3-benzothiazol-2-yl)-2-methoxyphenoxy)pentyl)oxy-(11aS)1,2,3,11a-tetra-hydro-5H-pyrrolo(2,1-c)(1,4)benzodiazepin-5-one
C3177676|7-MB-MP-PB cpd
C3712515|2-methyl-4-(4-methylpiperazin-1-yl)-10H-thieno(2,3-b)(1,5)benzodiazepine
C3181149|8-ethynyl-6-(2'-pyridine)-4H-2,5,10b-triazabenzo(e)azulene-3-carboxylic acid ethyl ester
C3829073|Midazolam-containing Buccal Liquid
C3851482|limazepine h
C3851484|limazepine G
C3886229|N-p-tosyl-1,5-benzodiazepin-2-one
C3886414|PGW5 compound
C3884716|oxoprothracarcin
C3884297|JM-20 compound
C3884297|3-ethoxycarbonyl-2-methyl-4-(2-nitrophenyl)-4,11-dihydro-1H-pyrido(2,3-b)(1,5)benzodiazepine
C3885219|QH-II-66
C4079047|diethyl-(Z)-2-(5,7-diphenyl-1,3,4-oxadiazepin-2-yl)-2-butenedioate
C0699927|Rohypnol
C0699927|Rohypnol (not approved for use in U.S.)
C0699927|Rohypnol (not approved for use in U.S.) (medication)
C0699927|Rohipnol
C0699927|Roche Brand of Flunitrazepam
C0699927|Narcozep
C0069749|10-chloro-2,3,7,11b-tetrahydro-2-methyl-11b-phenylbenzo(6,7)(1,4)diazepino(5,4-b) oxazol-6-one
C0069749|oxazolam
C0069749|oxazolazepam
C0060485|1-methyl-5-(2-fluorophenyl)-7-chloro-1,3-dihydro-2H-(1,4)benzodiazepin-2-one
C0060485|7-chloro-5-(2-fluorophenyl)-1,3-dihydro-1-methyl-2H-1,4-benzodiazepin-2-one
C0060485|fludiazepam
C0060485|fludiazepan
C0054826|5-(3-(4-piperidino-4-carbamoylpiperidino)propyl)- 10,11-dihydro-5(h)-dibenz(b,f)azepine
C0054826|carbadipimidine
C0054826|carpipramine
C0114875|1-(2-hydroxyethyl)-3-hydroxy-7-chloro-1,3-dihydro-5-(o-fluorophenyl)-2H-1,4-benzodiazepin-2-one
C0114875|doxefazepam
C0603384|7-chloro-5-(2-chlorophenyl)-1,3--dihydro-3-hydroxy-1-(2-hydroxyethyl)-2H-1,4-benzodiazepin-2-one
C0603384|N-(2-hydroxyethyl)lorazepam
C0604445|7-chloro-5-(2-fluorophenyl)-1,3-dihydro-1-(2-(methylsulfonyl)ethyl)-2H-1,4-benzodiazepin-2-one
C0604445|ID 622
C0604445|ID-622
C0604760|2H-1,5-Benzodiazepin-2-one, 8-chloro-1,3,4,5-tetrahydro-1-phenyl-
C0604760|8-chloro-1-phenyl-2,3,4,5-tetrahydro-1H-1,5-benzodiazepin-2-one
C0076784|1-(3,4-dimethoxyphenyl)-5-ethyl-7,8-dimethoxy- 4-methyl-5H-2,3-benzodiazepine
C0076784|tofisopam
C0076784|tofizopam
C0076784|1-(3,4-dimethoxyphenyl)-5-ethyl-7,8-dimethoxy-4-methyl-5H-2,3-benzodiazepine
C0060593|10-chloro-11b-(2'-fluorophenyl)-2,3,5,6,7,11b-hexahydro-7-(2''-hydroxyethyl)benzo(6,7)-1,4-diazepino(5,4-b)oxazol-6-one
C0060593|10-chloro-11b-(2-fluorophenyl)-2,3,7,11b-tetrahydro-7-(2-hydroxyethyl)oxazolo(3,2-d)(1,4)benzodiazepin-6(5H)-one
C0060593|flutazolam
C0076658|2-methyldiethylaminoethyl-4-p-phenylthiophenyl-3H- (1,5)benzodiazepine iodide
C0076658|thiabenzonium iodide
C0076658|tibenzonium iodide
C0076658|tibezonium
C0076658|Diethylmethyl(2-((4-(P-(Phenylthio)Phenyl)-3H-1,5-Benzodiazepin-2-yl)Thio)Ethyl)Ammonium
C0063325|ID 690
C0063325|ID-690
C0606744|7-chloro-5-(2-chlorophenyl)-1,3-dihydro-1-methyl-3-(4-morpholinylmethylene)-2H-1,4-benzodiazepin-2-one
C0606744|AX-A411-BS
C0055866|2H-1,4-Benzodiazepin-2-one, 7-chloro-1-(2-(cyclopropylmethoxy)ethyl)-1,3-dihydro-5-phenyl-
C0055866|7-chloro-1,3-dihydro-1-((2-cyclopropylmethoxy)ethyl)-5-phenyl-2H-1,4-benzodiazepin-2-one
C0055866|clazepam
C0073449|2H-1,4-Benzodiazepin-2-one, 1,3-dihydro-1-(methoxymethyl)-7-nitro-5-phenyl-
C0073449|Ro 06-9098-000
C0132831|N-desalkyl-2-oxoquazepam
C0132831|7-chloro-5-(2-fluorophenyl)-1,3-dihydro-2H-1,4- benzodiazepin-2-one
C0132831|norflutoprazepam
C0132831|norfludiazepam
C0132831|norflurazepam
C0073528|5-(2-fluorophenyl)-1,3-dihydro-1-methyl-2H-1,4- benzodiazepin-2-one
C0073528|Ro 5-3438
C0092802|2-chlorodiazepam
C0092802|2H-1,4-Benzodiazepin-2-one, 7-chloro-5-(2-chlorophenyl)-1,3-dihydro-1-methyl-
C0067928|1H-1,5-benzodiazepine-2,4(3H,5H)-dione, 8-chloro-1-phenyl-
C0067928|demethylclobazam
C0067928|N-desmethylclobazam
C0067928|norclobazam
C0611677|SAS 646
C0611797|Ka 2547
C0611797|Ka-2547
C0056431|CP 1414 S
C0056431|CP 1414S
C0056431|CP-1414 S
C0616152|4,5-dihydro-2,3-dimethyl-4-phenyl-3H-1,3-benzodiazepine
C0616486|psyton
C0076670|1-methyl-2-(3-thienylcarbonyl)aminomethyl-5-(2-fluorophenyl)-H-2,3-dihydro-1,4-benzodiazepine
C0076670|3-Thiophenecarboxamide, N-((5-(2-fluorophenyl)-2,3-dihydro-1-methyl-1H-1,4-benzodiazepin-2-yl)methyl)-
C0076670|tifluadom
C0076670|titfluadom
C0074103|SC 32855
C0074103|SC-32855
C0617110|5H-Pyrrolo(2,1-c)(1,4)benzodiazepin-5-one, 2-ethylidene-1,2,3,11a-tetrahydro-, (+)-
C0617110|prothracarcin
C0052237|1,3,4,14b-tetrahydro-2-methyl-10H-pyrazino-(1,2-a)pyrrolo(2,1-c)(1,4)benzodiazepine
C0052237|aptazapine
C0052237|2H,10H-Parazino(1,2-a)pyrrolo(2,1-c)(1,4)benzodiazepine,1,3,4,14b-tetrahydro-2-methyl-
C0047483|3-hydroxyphenazepam
C0047483|3-oxyfenazepam
C0061841|GP 55-129
C0061841|GP 55129
C0061841|GP-55129
C0073469|Ro 14-7437
C0073469|Ro-14-7437
C0093602|2-oxoquazepam
C0093602|2oxoquaz
C0093602|7-chloro-1-(2,2,2-trifluoroethyl)-1,3-dihydro-5-(2-fluorophenyl)-2H-1,4-benzodiazepin-2-one
C0619423|Sch 23-324
C0619423|Sch-23-324
C0619423|Sch 23324
C0147987|1-methyl-4-carbamoyl-5-phenyl-7-chloro-1,3,4,5-tetrahydro-2H-1,4-benzodiazepine-2-one
C0147987|4H-1,4-Benzodiazepine-4-carboxamide, 7-chloro-1,2,3,5-tetrahydro-1-methyl-2-oxo-5-phenyl-
C0147987|uxepam
C0099755|7-chloro-5-(2-fluorophenyl) 2,3-dihydro-2-oxo-1H-1,4-benzodiazepine-3-carboxylic acid
C0099755|loflazepic acid
C0621265|lepirazepam
C0055302|1,2,3,11a-tetrahydro-2,8-dihydroxy-7-methoxy-5H-pyrrolo(2,1-c)(1,4)-benzodiazepin-5-one
C0055302|5H-Pyrrolo(2,1-c)(1,4)benzodiazepin-5-one, 1,2,3,11a-tetrahydro-2,8-dihydroxy-7-methoxy-, (2S-trans)-
C0055302|chicamycin B
C0055301|1,2,3,10,11a-pentahydro-2,8-dihydroxy-7,11-dimethoxy-5H-pyrrolo(2,1-c)(1,4)-benzodiazepin-5-one
C0055301|5H-Pyrrolo(2,1-c)(1,4)benzodiazepin-5-one, 1,2,3,10,11,11a-hexahydro-2,8-dihydroxy-7,11-dimethoxy-, (2S-(2alpha,11alpha,11abeta))-
C0055301|chicamycin A
C0129948|N,N-dimethyl-6-phenyl-11H-pyrido(2,3-b)(1,4)benzodiazepin-11-propanamine
C0129948|11H-Pyrido(2,3-b)(1,4)benzodiazepine-11-propanamine, N,N-dimethyl-6-phenyl-, (E)-2-butenedioate (1:1)
C0129948|tampramine fumarate
C0073477|4H-Imidazo(1,5-a)(1,4)benzodiazepine-3-carboxylic acid, 8-azido-5,6-dihydro-5-methyl-6-oxo-, (Z,E,E,E,E)-
C0073477|Ro 15-4513
C0073477|RO-154513
C0073477|Ro15-4513
C0623223|7-chloro 5-(2-chlorophenyl)-1,3-dihydro-2H-(1,4)-benzodiazepine-2-thione
C0623223|7-CCDBT
C0073670|1H-Imidazo(1,2-a)(1,4)benzodiazepin-1-one, 6-(2-chlorophenyl)-2-((4-ethyl-1-piperazinyl)methylene)-2,4-dihydro-8-nitro-, (R-(R*,R*))-2,3-dihydroxybutanedioate (1:1)
C0073670|RU 32007
C0073670|RU-32007
C0623725|Pyrazino(1,2-a)(1,4)benzodiazepine, 1,2,3,4,4a,5-hexahydro-3-methyl-7-(2-thienyl)-
C0623725|KC 5944
C0623725|KC-5944
C0623750|Agarose, ((N,N'-1,2-ethanediylbis(N-(carboxymethyl)glycinato))(4-)-N,N',O,O',ON,ON')-, (2S-trans)-
C0623750|1012-S-acetamide adipic hydrazide Sepharose 4B
C0623750|BAAHS
C0164299|1-(3-chlorophenyl)-4-methyl-7,8-dimethoxy-5H-2,3-benzodiazepine
C0164299|girisopam
C0060496|7-fluoro-2-methyl-4(4-methyl-1-piperazinyl)-10H-thieno(2,3b)(1,5)benzodiazepine
C0060496|flumezapine
C0067931|N-desmethylmetaclazepam
C0073481|Ro 16-0521
C0073481|Ro-16-0521
C0073481|Urea, N-(6-bromo-5-(2-chlorophenyl)-2,3-dihydro-1,3-dimethyl-2-oxo-1H-1,4-benzodiazepin-7-yl)-N'-(2-hydroxy-1-(hydroxymethyl)-1-methylethyl)-, (S)-
C0628287|N-desmethylquazepam
C0066721|mono-N-demethyladinazolam
C0066721|mono-N-desmethyladin azolam
C0066721|N-desmethyladinazolam
C0066721|N-desmethyladinazolam mesylate
C0066721|N-desmethyladinozolam
C0066721|mono-N-demethyladinazolam mesylate
C0073534|Ro 7-0213
C0073534|Ro-7-0213
C0049851|7-BPDBD
C0049851|7-bromo-5-phenyl-1,2-dihydro-2H-1,4-benzodiazepin-2-one
C0085056|ZIMET 54-79
C0085056|ZIMET 5479
C0073510|Ro 23-0364
C0073510|Ro-23-0364
C0632104|N-demethyltimelotem
C0632104|N-desmethyltimelotem
C0635312|5H-Pyrrolo(2,1-c)(1,4)benzodiazepin-5-one, 7-((4,6-dideoxy-3-C-methyl-4-(methylamino)-alpha-L-mannopyranosyl)oxy)-1,2,3,11a-tetrahydro-2-propylidene-
C0635312|sibanomicin
C0636784|AHR 11797
C0636784|AHR-11797
C0044701|1012S
C0044701|compound 1012S
C0526445|Nerisopam
C0526445|1-(4-aminophenyl)-4-methyl-7,8-dimethoxy-5H-2,3-benzodiazepine
C0638880|6H-Imidazo(1,5-a)(1,4)benzodiazepin-6-one, 3-(5-cyclopropyl-1,2,4-oxadiazol-3-yl)-4,5-dihydro-5-methyl-
C0638880|FG 8119
C0638880|FG-8119
C0062021|Benzenamine, 4-(8-methyl-9H-1,3-dioxolo(4,5-h)(2,3)benzodiazepin-5-yl)-
C0062021|GYKI 52466
C0062021|GYKI-52466
C0639138|Acetamide, 2-(7-bromo-5-(2-fluorophenyl)-1,3-dihydro-1-methyl-2H-1,4-benzodiazepin-2-ylidene)-, (E)-
C0639138|KC 2846
C0639138|KC-2846
C0072934|R 82150
C0072934|R-82150
C0072934|R82150
C0083173|6H-Imidazo(1,5-a)(1,4)benzodiazepin-6-one, 7-chloro-4,5-dihydro-5-methyl-3-(5-(1-methylethyl)-1,2,4-oxadiazol-3-yl)-
C0083173|L 663581
C0083173|L-663581
C0641973|GYKI 52713
C0641973|GYKI-52713
C0643367|2-hydroxy-4-methylpyrimido(4,5-b)(1,5)benzodiazepin-5-one
C0643367|HMPBD
C0084281|Imidazo(4,5,1-jk)(1,4)benzodiazepine-2(1H)-thione, 9-chloro-4,5,6,7-tetrahydro-5-methyl-6-(3-methyl-2-butenyl)-, (S)-
C0084281|R 82913
C0084281|R-82913
C0084281|R82913
C0645521|Quinazolino(3',2':1,6)pyrido(2,3-b)(1,4)benzodiazepine-9,16-dione, 6,7,7a,8-tetrahydro-, (-)-
C0645521|auranthine
C0140776|Ro 24-7429
C0140776|Ro-24-7429
C0109226|CGS 15040A
C0109226|CGS-15040A
C0109226|2H,10H-Indolo(2,1-c)pyrazino(1,2-a)(1,4)benzodiazepine-16-carboxylic acid, 1,3,4,16b-tetrahydro-2-methyl-, methyl ester, monohydrochloride
C0147541|U-46,195
C0147541|U46,195
C0147541|U-46195
C0147541|U 46195
C0649797|7-(4-bromophenyl)-8-phenoxy-4,5-benzo-3-aza-2-nonem
C0649797|7-BPPBAN
C0168533|BIM-18216
C0168533|BIM 18216
C0653743|biotin-(N-(2-aminoethyl)-8-chloro-6-(2-chlorophenyl)-4H(1,2,4)triazolo(3,4-a)(1,4)benzodiazepine-2-carboxamide) conjugate
C0653743|biotinylated 1012-S conjugate
C0653743|biotin-1012-S
C0656355|12,13,14,14a-tetrahydro-9H,11H-pyrazino(2,1-c)pyrrolo(1,2-a)(1,4)benzodiazepine
C0656355|isonoraptazepine
C0213386|GYKI-53655
C0213386|GYKI 53655
C0660404|U-51477
C0660404|U 51477
C0660406|U-34599
C0660406|U 34599
C0660406|4H-(1,2,4)Triazolo(4,3-a)(1,4)diazepine, 8-chloro-1,4-dimethyl-6-phenyl-
C0219102|6-(2-bromophenyl)-8-fluoro-4-H-imidazo(1,5-a)(1-4)benzodiazepine-3-carboxamide
C0219102|imidazenil
C0661222|4-BDBDT
C0661222|4-(3-bromophenyl)-1,3-dihydro-2H-1,5-benzodiazepin-2-thione
C0249301|tripitramine
C0250723|GYKI 53405
C0250723|GYKI-53405
C0252422|9a,9b,14b,14c-tetraphenylbenzo(1,2-h-4,5-h')dicyclohepta(1,2,3-bc)glycoluril
C0252422|TPB-DCHU
C0252468|R 86183
C0252468|R-86183
C0252468|R86183
C0254734|L 368935
C0254734|L-368,935
C0254734|Urea, N-(2,3-dihydro-1-(2-methylpropyl)-2-oxo-5-phenyl-1H-1,4-benzodiazepin-3-yl)-N'-(3-(1H-tetrazol-5-yl)phenyl)-, (R)-
C0254783|YM 022
C0254783|YM-022
C0254783|YM022
C0254783|Urea, N-(2,3-dihydro-1-(2-(2-methylphenyl)-2-oxoethyl)-2-oxo-5-phenyl-1H-1,4-benzodiazepin-3-yl)-N'-(3-methylphenyl)-, (R)-
C0257405|benzomalvin A
C0257406|benzomalvin B
C0257407|benzomalvin C
C0289297|1,1-bis(((5,11-dihydro-6-oxo-6H-pyrido(2,3-b)(1,4)benzodiazepin-11-yl)carbonyl)methyl)-8,17-dimethyl-1,8,17,24-tetraazatetracosane
C0289297|dipitramine
C0290224|BZA 5B
C0290224|BZA-5B
C0294497|R 79882
C0294497|R-79882
C0294497|R79882
C0383534|Ro 14-5974
C0383534|Ro 145974
C0383534|Ro-14-5974
C0383534|Ro-145974
C0383538|Ro 19-0528
C0383538|Ro 190528
C0383538|Ro-19-0528
C0383538|Ro-190528
C0385516|8-chloro-TIBO
C0385516|8-chlorotetrahydroimidazo(4,5,1-jk)(1,4)-benzodiazepin-2(1H)-thione
C0385516|Tivirapine
C0385516|(S)-8-Chloro-4,5,6,7-tetrahydro-5-methyl-6-(3-methyl-2-butenyl)imidazo(4,5,1-jk)(1,4)benzodiazepine-2(1H)-thione
C0077112|1-methyl-5-phenyl-7-trifluoromethyl-(1H)-1,5-benzodiazepine-2,4-(3H,5H)dione
C0077112|triflubazam
C0391429|NNC 13-8241
C0391429|NNC-13-8241
C0531537|9-amino-11-ethyl-6-methylpyrido(2,3-b)(1,4)benzodiazepin-5-one
C0531537|9-aminonevirapine
C0532436|sarmazenil
C0532436|Ethyl 7-chloro-5,6-dihydro-5-methyl-6-oxo-4H-imidazo-(1,5-a)(1,4)benzodiazepine-3-carboxylate
C0536423|1-(3-(N'-(4-(2-(N-aminosulfonylamidino)ethylthiomethyl)thiazol-2-yl)guanidinomethyl)phenyl)-3-(1-methyl-2-oxo-5-phenyl-2,3-dihydro-1H-1,4-benzodiazepin-3-yl)urea
C0536423|AETGPMOPDBU
C0537435|GYKI 53665
C0537435|GYKI-53665
C0538541|EGIS 7649
C0538541|EGIS-7649
C0538838|S 8510
C0538838|S-8510
C0540410|7-chloro-1,3-dihydro-3-hemisuccinyloxy-5-phenyl-1,4-benzodiazepin-2-one
C0541175|Ro 48-6792
C0541355|4,5,6,7-tetrahydro-5-methylimidazo(4,5,1-jk)(1,4)benzodiazepin-2(1H)-one
C0541355|4567-TMB
C0667114|7-chloro-1,3-dihydro-1-(1,1-dimethylethyl)-5-(2-fluorophenyl)-2H-1,4-benzodiazepin-2-one
C0667114|7-CDDFB
C0667714|RY80
C0667714|RY 80
C0670249|Ro 48-8684
C0670792|BDA 452
C0670792|BDA-452
C0670792|BDA452
C0670796|BDA 250
C0670796|BDA-250
C0670796|BDA250
C0755389|L-364,373
C0755389|L 364373
C0755389|L364373
C0756415|RY-008, imidazobenzodiazepine
C0756415|RY 008
C0756868|1-(4'-aminophenyl)-3,5-dihydro-7,8-dimethoxy-4H-2m3-benzodiazepine-4-thione
C0756868|1-NHPh-DDBT
C0759918|RL 218
C0759918|RL-218
C0759921|RL 236
C0759921|RL-236
C0760184|TS 941
C0760184|TS-941
C0760184|TS941
C0760535|L 735,821
C0760535|L-735,821
C0760535|L 735821
C0760535|L-735821
C0761079|CR 2945
C0761079|CR-2945
C0761079|CR2945
C0764989|tarazepide
C0764989|(-)-N-((S)-2,3-Dihydro-1-methyl-2-oxo-5-phenyl-1H-1,4-benzodiazepin-3-yl)-5,6-dihydro-4H-pyrrolo(3,2,1-ij)quinoline-2-carboxamide
C0765506|DMP 406
C0765506|DMP-406
C0766295|GYKI 53784
C0766295|GYKI-53784
C0768431|LE 511
C0768431|LE-511
C0768431|LE511
C0907968|1-(4'-aminophenyl)-3,5-dihydro-7,8--dimethoxy-2,3-benzodiazepine
C0907968|2,3-BZ cpd
C0908355|VP 339
C0908355|VP-339
C0908356|VP 365
C0908356|VP-365
C0908672|7-bromo-5-phenyl-dihydro-3H-1,4-benzodiazepine
C0908672|7-bromo-PhHBDZ
C0909356|CL 385,004
C0909356|CL 385004
C0909356|CL-385,004
C0909356|CL-385004
C0914661|tetrazolo(1,5-a)(1,4)benzodiazepine
C0914662|triazolo(4,3-d)benzodiazepine
C0960422|Lotrafiban
C0961688|4-phenyl-2-trichloromethyl-3H-1,5-benzodiazepine
C1306120|7-cyano-2,3,4,5-tetrahydro-1-(1H-imidazol-4-ylmethyl)-3-(phenylmethyl)-4-(2-thienylsulfonyl)-1H-1,4-benzodiazepine
C0963297|1,5-benzodiazepin-2-one
C0963508|GYKI 47261
C0963508|GYKI-47261
C0967164|1,2,3,4-tetrahydrobenzo(e)(1,4)diazepin-5-one
C0967164|TH-BDAO
C0969588|8-fluoro-12-(4-methylpiperazin-1-yl)-6H-(1)benzothieno(2,3-b)(1,5)benzodiazepine
C0969588|8-fluoro-12-(4-methylpiperazin-1-yl)-6H-(1)benzothieno(2,3-b)(1,5)benzodiazepine maleate
C0969588|Y 931
C1097584|ethyl-8-ethyl-5,6-dihydro-5-methyl-6-oxo-4H-imidazo(1,5a)(1,4)benzodiazepine-3-carboxylate
C1097588|ETADOAIB cpd
C1097588|ethyl-8-trimethylsilyl-2-acetyl-12,12a-dihydro-9-oxo-9H,11H-azeto(2,1-c)imidazo(1,5a)-1,4-benzodiazepine
C1098285|BZA-2B
C1098285|Cys-(N-methyl)-3-amino-1-carboxymethyl-2,3-dihydro-5-phenyl-1H-1,4-benzodiazepin-2-one-Met
C1098621|circumdatin C
C1434719|PBDS cpd
C1434719|pyrrolo(2,1-c)(1,4)benzodiazepine
C1136832|BD-1158
C1143145|RY 024
C1143145|RY024
C1143677|3-tert-butoxycarbonylamino-2-oxo-2,3,4,5-tetrahydro-1,5-benzodiazepine-1-acetic acid methyl ester
C1143677|BTOTBAM ester
C1143762|1-M-6P-TBD
C1143762|1-methyl-6-phenyl-4H-s-triazo-(4,3-alpha)(1,4)benzodiazepinone
C1172344|1,4-benzodiazepine
C1172344|Bz-423
C1172477|6-chloro-PPPBD
C1172477|8-chloro-6-(4-phenethyl-1-piperazinyl)-11H-pyrido(2,3-b)(1,4)benzodiazepine
C1173066|Indiplon
C1174538|5-P-3-U-BDA
C1174538|5-phenyl-3-ureido-1,5-benzodiazepine
C1311127|(11aS)-8-hydroxy-7-methoxy-1,2,3,11a-tetrahydro-5H-pyrrolo(2,1-c)(1,4)benzodiazepin-5-one
C1311268|TIBO cpd
C1311268|4,5,6,7-tetrahydroimidazo-(4,5,1- jk)(1,4)benzodiazepin-2 (1 H)-one
C1311387|8,9-dimethoxy-6-(4-bromophenyl)-11H-(1,2,4)triazolo(4,5-c)(2,3)benzodiazepin-3(2H)-one
C1311387|8,9-dimethoxy-BTBDO
C1313512|1-(4-dimethylaminomethylphenyl)-8,9-dihydro-7H-2,7,9a-benzo(cd)azulen-6-one
C1435117|2,3,4,5-tetrahydro-1-(1H-imidazol-4-ylmethyl)-4-(2-biphenylylcarbonyl)-1H-1,4-benzodiazepine
C1454299|BMS-225975
C1454299|BMS225975
C1505431|GI 181771X
C1505431|GI-181771X
C1505431|GI181771X
C1608551|FLUOXETINE/OLANZAPINE
C1608551|Fluoxetine / olanzapine
C1608551|FLUoxetine-OLANZapine
C1608551|Olanzapine + fluoxetine (product)
C1608551|Olanzapine + fluoxetine
C1608551|olanzapine-fluoxetine combination
C1570489|mmy-SJG compound
C1571352|FQP-BD cpd
C1571352|fluoroquinolone-pyrrolo(2,1-c)(1,4)benzodiazepine
C1611910|2,3-dimethyl-6-phenyl-12H-(1,3)dioxolo(4,5-h)imidazo(1,2-c)(2,3)benzodiazepine
C1615028|EGIS-10608
C1614477|EGIS-8332
C1687864|RY 023
C1686352|6-fluoro-10-(3-(2-methoxyethyl)-4-methylpiperazin-1-yl)-2-methyl-4H-3-thia-4,9-diazabenzo(f)azulene
C1698804|RWJ-351647
C1700769|DPBDA cpd
C1700769|5,11-dihydro-pyrido(2,3-b)(1,5)benzodiazepine
C1721896|alpha5IA-II
C1871751|RO0281501
C1871751|RO 0281501
C1872487|2-hydroxymethylolanzapine
C1870086|DRH-417
C1870086|NSC 709119
C1880572|Ethyl Carfluzepate
C1880826|Flutemazepam
C1882473|Proflazepam
C0209249|2-benzoyl-6-ethyl-7-methoxy-5-methylimidazol(1,2-a)pyrimidine
C0209249|Methanone, (6-ethyl-7-methoxy-5-methylimidazo(1,2-a)pyrimidin-2-yl)phenyl-
C0209249|divaplon
C0700528|Hydrochloride, Chlordiazepoxide
C0700528|Chlordiazepoxide Hydrochloride
C0700528|chlordiazepoxide hydrochloride (medication)
C0700528|Chlordiazepoxide Hydrochloride [Chemical/Ingredient]
C0700528|Chlordiazepoxide Monohydrochloride
C0700528|Monohydrochloride, Chlordiazepoxide
C0700528|Chlordiazepoxide hydrochloride (substance)
C0700528|Chlordiazepoxide hydrochloride (product)
C0770393|CLORAZEPIC ACID
C1881125|Iclazepam
C1881782|Menitrazepam
C0071879|3,7-dihydro-5-phenyl-6,7-dimethylpyrrole(3,4-e)(1,4)diazepin-2-(1H)-one
C0071879|premazepam
C0035766|Hydrochloride, Medazepam
C0035766|Medazepam Hydrochloride
C0035766|Monohydrochloride, Medazepam
C0035766|Medazepam Monohydrochloride
C1880574|Ethyl Dirazepate
C0700457|Hydrochloride, Midazolam
C0700457|Midazolam Hydrochloride
C0700457|anxiolytics midazolam hydrochloride
C0700457|midazolam hydrochloride (medication)
C0700457|Midazolam Hydrochloride [Chemical/Ingredient]
C0700457|midazolam (as hydrochloride)
C0700457|Midazolam hydrochloride (product)
C0700457|Midazolam hydrochloride (substance)
C3179470|remimazolam
C2000107|4-(2-hydroxyphenyl)-2-phenyl-2,3-dihydro-1H-1,5-benzodiazepine
C2000107|4-(2-hydroxyphenyl)-PDBDZ
C0065086|lithium bromide
C0065086|Lithium bromide (substance)
C0978225|Lithium Carbonate 150 MG Oral Capsule
C0978225|Lithium Carbonate 150mg Oral capsule
C0978225|Lithium Carbonate, 150 mg oral capsule
C0978225|lithium 150 mg oral capsule
C0978225|LITHIUM CARBONATE 150MG CAP
C0978225|LITHIUM CARBONATE 150MG CAP UD
C0978225|lithium carbonate 150 MILLIGRAM In 1 CAPSULE ORAL CAPSULE
C0978225|Lithium Carbonate Cap 150 MG
C0978225|LITHIUM CARBONATE 150 mg ORAL CAPSULE, GELATIN COATED
C0978225|LITHIUM CARBONATE 150MG CAP,UD [VA Product]
C0978225|LITHIUM CARBONATE 150MG CAP,UD
C0978225|LITHIUM CARBONATE 150MG CAP [VA Product]
C0978225|LITHIUM CARBONATE 150 mg ORAL CAPSULE [LITHIUM CARBONATE]
C0978225|LiCO3 150 MG Oral Capsule
C0978225|Lithium carbonate 150mg capsule (product)
C0978225|Lithium carbonate 150mg capsule
C0689383|Lithium Carbonate 300 MG Oral Capsule
C0689383|Lithium Carbonate 300mg Oral capsule
C0689383|Lithium Carbonate, 300 mg oral capsule
C0689383|lithium 300 mg oral capsule
C0689383|LITHIUM CARBONATE 300MG CAP
C0689383|lithium carbonate 300 MILLIGRAM In 1 CAPSULE ORAL CAPSULE
C0689383|Lithium Carbonate Cap 300 MG
C0689383|LITHIUM CARBONATE 300 mg ORAL CAPSULE, GELATIN COATED
C0689383|LITHIUM CARBONATE 300MG CAP [VA Product]
C0689383|LITHIUM CARBONATE 300 mg ORAL CAPSULE [LITHIUM CARBONATE]
C0689383|LiCO3 300 MG Oral Capsule
C0689383|Lithium carbonate 300mg capsule (product)
C0689383|Lithium carbonate 300mg capsule
C0689384|Lithium Carbonate 300 MG Oral Tablet
C0689384|Lithium Carbonate 300mg Oral tablet
C0689384|Lithium Carbonate, 300 mg oral tablet
C0689384|lithium 300 mg oral tablet
C0689384|LITHIUM CARBONATE 300MG TAB
C0689384|Lithium Carbonate Tab 300 MG
C0689384|LITHIUM CARBONATE 300MG TAB [VA Product]
C0689384|LiCO3 300 MG Oral Tablet
C0689384|Lithium carbonate 300mg tablet (product)
C0689384|Lithium carbonate 300mg tablet
C0689385|Lithium Carbonate 300 MG Oral Tablet, Extended Release
C0689385|Lithium Carbonate 300mg Oral tablet, extended release
C0689385|lithium 300 mg oral tablet, extended release
C0689385|LITHIUM CARBONATE 300MG SA TAB
C0689385|Lithium Carbonate Tab CR 300 MG
C0689385|Lithium carbonate 300mg slow release tablet
C0689385|LITHIUM CARBONATE 300 mg ORAL TABLET, FILM COATED, EXTENDED RELEASE
C0689385|LITHIUM CARBONATE 300MG TAB,SA
C0689385|LITHIUM CARBONATE 300MG TAB,SA [VA Product]
C0689385|LITHIUM CARBONATE 300 mg ORAL TABLET, EXTENDED RELEASE [LITHIUM CARBONATE]
C0689385|LITHIUM CARBONATE 300 mg ORAL TABLET, FILM COATED, EXTENDED RELEASE [Lithium Carbonate]
C0689385|Lithium Carbonate 300 MG Extended Release Oral Tablet
C0689385|LiCO3 300 MG Extended Release Oral Tablet
C0689385|Lithium Carbonate, 300 mg oral tablet, extended release
C0689385|Lithium carbonate 300mg m/r tablet
C0689385|Lithium carbonate 300mg m/r tablet (product)
C0689386|Lithium Carbonate 450 MG Oral Tablet, Extended Release
C0689386|Lithium Carbonate 450mg Oral tablet, extended release
C0689386|Lithium carbonate 450mg tablet
C0689386|lithium 450 mg oral tablet, extended release
C0689386|LITHIUM CARBONATE 450MG SA TAB
C0689386|Lithium Carbonate Tab CR 450 MG
C0689386|LITHIUM CARBONATE 450MG TAB,SA [VA Product]
C0689386|LITHIUM CARBONATE 450MG TAB,SA
C0689386|LITHIUM CARBONATE 450 mg ORAL TABLET, EXTENDED RELEASE [LITHIUM CARBONATE]
C0689386|Lithium carbonate cr 450mg tablet (product)
C0689386|Lithium carbonate cr 450mg tablet
C0689386|lithium carbonate 450 MG Extended Release Oral Tablet
C0689386|LiCO3 450 MG Extended Release Oral Tablet
C0689386|LITHIUM CARBONATE 450 mg ORAL TABLET [Lithium Carbonate ER]
C0689386|Lithium carbonate 450mg m/r tablet
C0689386|Lithium carbonate 450mg m/r tablet (product)
C0689386|Lithium Carbonate, 450 mg oral tablet, extended release
C0689386|Lithium carbonate 450mg m/r tablet (substance)
C0689386|Lithium carbonate 450mg tablet (product)
C0689387|Lithium Carbonate 600 MG Oral Capsule
C0689387|Lithium Carbonate 600mg Oral capsule
C0689387|Lithium Carbonate, 600 mg oral capsule
C0689387|lithium 600 mg oral capsule
C0689387|LITHIUM CARBONATE 600MG CAP
C0689387|lithium carbonate 600 MILLIGRAM In 1 CAPSULE ORAL CAPSULE
C0689387|Lithium Carbonate Cap 600 MG
C0689387|LITHIUM CARBONATE 600 mg ORAL CAPSULE, GELATIN COATED
C0689387|LITHIUM CARBONATE 600MG CAP [VA Product]
C0689387|LiCO3 600 MG Oral Capsule
C0689387|Lithium carbonate 600mg capsule (product)
C0689387|Lithium carbonate 600mg capsule
C0700189|Lithonate
C0771417|Lithium Salicylate
C0700753|Eskalith
C0700753|Escalith
C0700751|Lithobid
C0700752|Lithane
C0065091|lithium orotate
C2716130|potassium lithium titanate
C1966347|Lithium Aspartate
C1966347|antimanics lithium aspartate
C1966347|lithium aspartate (medication)
C0689381|Lithium 8 MEQ/5 ML Oral Solution
C0689381|Lithium Citrate 8mEq/5mL Oral solution
C0689381|lithium citrate 60 MG/ML Oral Solution
C0689381|LITHIUM CITRATE 8MEQ/5ML SF SYRUP
C0689381|Lithium Hydroxide Monohydrate 8 meq in 5 mL ORAL SOLUTION
C0689381|Lithium Citrate 8mEq/5mL Oral syrup
C0689381|Lithium Citrate 8 MEQ/5 ML Oral Solution
C0689381|LITHIUM CITRATE 8MEQ/5ML SYRUP
C0689381|LITHIUM CITRATE 8MEQ/5ML (SF) SYRUP
C0689381|LITHIUM CITRATE 8MEQ/5ML (SF) SYRUP [VA Product]
C0689381|LITHIUM CITRATE 8MEQ/5ML SYRUP [VA Product]
C0689381|LITHIUM CARBONATE 8 meq in 5 mL ORAL SOLUTION [Lithium]
C0689381|Lithium Citrate 8mEq/5ml Solution
C0689381|Lithium 8mEq/5mL Oral solution
C0689381|Lithium 8mEq/5ml Solution
C0689381|LITHIUM 8MEQ/5ML SOLN,ORAL
C0689381|LITHIUM 8MEQ/5ML ORAL SOLN
C0689381|LITHIUM 8MEQ/5ML SOLN,ORAL [VA Product]
C0689381|lithium ion 8 MEQ per 5 ML Oral Syrup
C0689381|lithium citrate eqv to lithium carbonate 300 MG per 5 ML (lithium ion 8 MEQ per 5 ML) Oral Syrup
C0689381|Lithium carbonate 300 mg in 5 mL ORAL SOLUTION [Lithium]
C0689381|LITHIUM CITRATE 8 meq in 5 mL ORAL SOLUTION
C0689381|Lithium Oral Solution 8 mEq/5ML
C0689381|Lithium Citrate 300 MG/5 ML Oral Syrup
C0689381|Lithium Citrate, 300 mg/5 mL oral syrup
C0689381|lithium 300 mg/5 mL oral syrup
C0693401|Lithium Carbonate 400 MG Oral Tablet, Extended Release
C0693401|LiCO3 400 MG Extended Release Oral Tablet
C0693401|lithium carbonate 400 MG Extended Release Oral Tablet
C0693401|Lithium carbonate 400mg m/r tablet
C0693401|Lithium carbonate 400mg m/r tablet (product)
C0693401|Lithium carbonate 400mg m/r tablet (substance)
C0350511|Lithium Carbonate 104 MG/ML Oral Solution
C0350511|lithium carbonate 520 MG per 5 ML Oral Solution
C0350511|LiCO3 104 MG/ML Oral Solution
C0350511|Lithium carbonate 520mg/5mL sugar free liquid (product)
C0350511|Lithium carbonate 520mg/5mL sugar free liquid
C0350511|Lithium carbonate 520mg/5mL sugar free liquid (substance)
C0692744|Lithium Carbonate 250 MG Oral Tablet
C0692744|LiCO3 250 MG Oral Tablet
C0692744|Lithium carbonate 250mg tablet
C0692744|Lithium carbonate 250mg tablet (product)
C0692744|Lithium carbonate 250mg tablet (substance)
C0789694|Lithium Carbonate 200 MG Extended Release Oral Tablet
C0789694|LiCO3 200 MG Extended Release Oral Tablet
C0789694|Lithium carbonate 200mg m/r tablet
C0789694|Lithium carbonate 200mg m/r tablet (product)
C0789694|Lithium carbonate 200mg m/r tablet (substance)
C0302213|LITHIUM SALTS
C0302213|[CN750] LITHIUM SALTS
C0302213|Lithium salt
C0302213|Lithium salt (substance)
C0302213|Lithium salt, NOS
C0065093|lithium succinate
C0065093|Lithium succinate (product)
C0065093|lithium succinate (medication)
C0065093|antimanics lithium succinate
C0065093|Lithium succinate (substance)
C1991690|Lithium &#x7C; body fluid
C1991692|Lithium &#x7C; red blood cells
C2738318|Lithium &#x7C; Gastric fluid
C0366526|Lithium:Mass:Pt:Dose:Qn
C0366526|Lithium Dose
C0366526|Lithium [Mass] of Dose
C0366526|Lithium:Mass:Point in time:Dose med or substance:Quantitative
C1991694|Lithium &#x7C; Tissue and Smears
C1991695|Lithium &#x7C; urine
C1991691|Lithium &#x7C; hair
C1991696|Lithium &#x7C; Urine and Serum or Plasma
C1991693|Lithium &#x7C; saliva
C1991688|Lithium &#x7C; bld-ser-plas
C3495095|Lithium Cation
C3495095|Li+
C3495095|Lithium Ion
C0303507|Lithium isotope
C0303507|Lithium isotope (substance)
C0078149|Veinobiase
C1121051|noolith
C1122689|dysprosium lithium borate glass
C1175911|LiTaO3
C1175911|lithium tantalate oxide
C1175913|LiFePO4
C1311954|Li2ZrO3
C1311954|lithium zirconate
C1455455|LiMn2O4
C1455455|lithium manganese oxide
C0287163|Seroquel
C0287163|quetiapine (Seroquel)
