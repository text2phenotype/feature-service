C0948762|Absolute neutrophil count
C1168174|Absolute neutrophil count decreased
C1262264|Absolute neutrophil count abnormal
C1699112|Absolute neutrophil count increased
C0362968|Neutrophils # Bld Auto
C0948762|Absolute neutrophil count
C0948762|ANC
C0948762|blood absolute neutrophil count (ANC)
C0948762|blood absolute neutrophil count (ANC) (lab test)
C0948762|blood ANC
C0948762|blood absolute neutrophil count
C0948762|blood absolute granulocyte count
C0948762|blood ANC (absolute neutrophil count)
C0948762|blood absolute neutrophil count (lab test)
C0948762|Neutrophils
C0948762|NEUT
C1168174|Decreased ANC
C1168174|Decreased Absolute Neutrophil Count
C1168174|Absolute neutrophil count decreased
C1262264|Absolute neutrophil count abnormal
C1699112|Absolute neutrophil count increased
C0362968|Neutrophils # Bld Auto
C0362968|Neutrophils:NCnc:Pt:Bld:Qn:Automated count
C0362968|Neutrophils [#/volume] in Blood by Automated count
C0362968|Neutrophils:Number Concentration (count/vol):Point in time:Whole blood:Quantitative:Automated count
