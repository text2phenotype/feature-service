C2239176|Liver carcinoma
C2239176|Liver cell carcinoma
C2239176|Carcinoma, Hepatocellular
C2239176|Carcinomas, Hepatocellular
C2239176|Hepatocellular Carcinomas
C2239176|Hepatoma
C2239176|Hepatomas
C2239176|hepatocellular carcinoma
C2239176|LCC
C2239176|carcinoma of liver (diagnosis)
C2239176|hepatocellular carcinoma of liver (diagnosis)
C2239176|hepatocellular carcinoma of liver
C2239176|liver neoplasm malignant carcinoma
C2239176|carcinoma of liver
C2239176|Liver carcinoma
C2239176|Liver Cell Cancer (Hepatocellular Carcinoma)
C2239176|Carcinoma, Hepatocellular [Disease/Finding]
C2239176|Cancers, Adult Liver
C2239176|Adult Liver Cancer
C2239176|Cancer, Adult Liver
C2239176|Adult Liver Cancers
C2239176|Liver Cancers, Adult
C2239176|Liver Cancer, Adult
C2239176|Liver Cell Carcinoma, Adult
C2239176|Liver Cell Carcinomas
C2239176|Cell Carcinoma, Liver
C2239176|Cell Carcinomas, Liver
C2239176|Carcinoma, Liver Cell
C2239176|Carcinomas, Liver Cell
C2239176|Hepatic cell carcinoma
C2239176|Primary carcinoma of liver
C2239176|liver neoplasm malignant carcinoma primary
C2239176|Primary carcinoma of liver (diagnosis)
C2239176|HCC
C2239176|CARCINOMA, HEPATOCELLULAR, MALIGNANT
C2239176|[M]Hepatocellular carcinoma NOS
C2239176|Carcinoma of the Liver Cells
C2239176|Primary Carcinoma of the Liver Cells
C2239176|Carcinoma of Liver Cells
C2239176|Primary Carcinoma of Liver Cells
C2239176|Liver cell carcinoma (clinical)
C2239176|Hepatocellular carcinoma (clinical)
C2239176|Carcinoma liver
C2239176|Carcinoma hepatocellular
C2239176|Hepatocarcinoma
C2239176|Hepatoma, malignant
C2239176|Malignant hepatoma
C2239176|LCC - Liver cell carcinoma
C2239176|HCC - Hepatocellular carcinoma
C2239176|Hepatocellular carcinoma (morphologic abnormality)
C2239176|Liver cell carcinoma (disorder)
C2239176|Primary carcinoma of liver (disorder)
C2239176|carcinoma; hepatic cell
C2239176|carcinoma; hepatocellular
C2239176|hepatic cell; carcinoma
C2239176|hepatocellular; carcinoma
C2239176|Hepatocellular carcinoma, NOS
C2239176|Hepatoma, NOS
C2239176|Carcinoma of liver, specified as primary
C2239176|Carcinoma of liver cell
C2205336|malignant epithelioma of liver
C2205336|liver neoplasm malignant carcinoma epithelioma
C2205336|malignant epithelioma of liver (diagnosis)
C2111635|large cell carcinoma of liver
C2111635|large cell carcinoma of liver (diagnosis)
C2012092|glassy cell carcinoma of liver (diagnosis)
C2012092|glassy cell carcinoma of liver
C2205337|anaplastic carcinoma of liver (diagnosis)
C2205337|anaplastic carcinoma of liver
C2205337|liver neoplasm malignant carcinoma anaplastic
C2082443|pleomorphic carcinoma of liver
C2082443|pleomorphic carcinoma of liver (diagnosis)
C2011254|giant cell carcinoma of liver (diagnosis)
C2011254|giant cell carcinoma of liver
C2018394|spindle cell carcinoma of liver
C2018394|spindle cell carcinoma of liver (diagnosis)
C2011218|giant cell and spindle cell carcinoma of liver (diagnosis)
C2011218|liver neoplasm malignant carcinoma giant cell & spindle cell
C2011218|giant cell and spindle cell carcinoma of liver
C2142923|pseudosarcomatous carcinoma of liver (diagnosis)
C2142923|pseudosarcomatous carcinoma of liver
C2111805|polygonal cell carcinoma of liver (diagnosis)
C2111805|polygonal cell carcinoma of liver
C0334286|Biliary Cystadenocarcinoma
C0334286|cystadenocarcinoma of bile duct
C0334286|cystadenocarcinoma of bile duct (diagnosis)
C0334286|liver neoplasm malignant bile duct cystadenocarcinoma
C0334286|Bile Duct Mucinous Cystic Neoplasm with an Associated Invasive Carcinoma
C0334286|Bile Duct Cystadenocarcinoma
C0334286|Bile duct cystadenocarcinoma (morphologic abnormality)
C0334286|bile duct; cystadenocarcinoma
C0334286|cystadenocarcinoma; bile duct
C0334286|Cystadenocarcinoma of the Bile Duct
C2076526|infiltrating ductal carcinoma of liver (diagnosis)
C2076526|infiltrating ductal carcinoma of liver
C2106546|comedocarcinoma of liver
C2106546|liver neoplasm malignant carcinoma comedocarcinoma
C2106546|comedocarcinoma of liver (diagnosis)
C2078053|intracystic carcinoma of liver (diagnosis)
C2078053|intracystic carcinoma of liver
C2047535|hypersecretory cystic carcinoma of liver (diagnosis)
C2047535|liver neoplasm malignant carcinoma cystic hypersecretory
C2047535|hypersecretory cystic carcinoma of liver
C2064401|undifferentiated carcinoma of liver (diagnosis)
C2064401|undifferentiated carcinoma of liver
C2064401|Undifferentiated Liver Carcinoma
C2064401|Undifferentiated Primary Liver Carcinoma
C0334287|fibrolamellar hepatocellular carcinoma of liver (diagnosis)
C0334287|fibrolamellar hepatocellular carcinoma of liver
C0334287|Fibrolamellar variant of hepatocellular carcinoma
C0334287|Fibrolamellar hepatocellular carcinoma
C0334287|Hepatocellular carcinoma (fibrolamellar variant)
C0334287|FLC
C0334287|Fibrolamellar Carcinoma
C0334287|[M]Hepatocellular carcinoma, fibrolamellar
C0334287|[M] Hepatocellular carcinoma, fibrolamellar
C0334287|Hepatocellular carcinoma, fibrolamellar
C0334287|Fibrolamellar hepatocellular carcinoma (disorder)
C0334287|Hepatocellular carcinoma, fibrolamellar (morphologic abnormality)
C0334287|carcinoma; hepatocellular, fibrolamellar
C0334287|fibrolamellar; hepatocellular carcinoma
C0334287|hepatocellular; carcinoma, fibrolamellar
C0334287|Fibrolamellar Carcinoma of Liver Cells
C0334287|Fibrolamellar Carcinoma of the Liver Cells
C0334287|Hepatocellular Fibrolamellar Carcinoma
C0334287|Liver Cell Fibrolamellar Carcinoma
C0334287|Oncocytic Hepatocellular Tumor
C0334287|Polygonal Cell Type Hepatocellular Carcinoma with Fibrous Stroma
C2205338|scirrhous hepatocellular carcinoma of liver (diagnosis)
C2205338|scirrhous hepatocellular carcinoma of liver
C1266019|spindle cell hepatocellular carcinoma of liver
C1266019|spindle cell hepatocellular carcinoma of liver (diagnosis)
C1266019|Hepatocellular carcinoma, sarcomatoid
C1266019|Hepatocellular carcinoma, spindle cell variant (morphologic abnormality)
C1266019|Hepatocellular carcinoma, spindle cell variant
C1266020|clear cell hepatocellular carcinoma of liver (diagnosis)
C1266020|clear cell hepatocellular carcinoma of liver
C1266020|Hepatocellular carcinoma, clear cell type (morphologic abnormality)
C1266020|Hepatocellular carcinoma, clear cell type
C2082477|pleomorphic hepatocellular carcinoma of liver
C2082477|pleomorphic hepatocellular carcinoma of liver (diagnosis)
C0221287|hepatocellular carcinoma and cholangiocarcinoma
C0221287|liver neoplasm hepatocellular carcinoma & cholangiocarcinoma
C0221287|hepatocellular carcinoma and cholangiocarcinoma (diagnosis)
C0221287|Mixed hepatocellular cholangiocarcinoma
C0221287|[M]Combined hepatocellular carcinoma and cholangiocarcinoma
C0221287|Combined hepatocellular and cholangiocarcinoma
C0221287|Hepatocholangiocarcinoma
C0221287|Mixed hepatocellular and bile duct carcinoma
C0221287|Combined hepatocellular carcinoma and cholangiocarcinoma
C0221287|Combined hepatocellular carcinoma and cholangiocarcinoma (disorder)
C0221287|Combined hepatocellular carcinoma and cholangiocarcinoma (morphologic abnormality)
C0221287|cholangiocarcinoma; with hepatocellular carcinoma
C0221287|cholangiohepatoma
C0221287|hepatocellular carcinoma; cholangiocarcinoma
C0221287|Liver and Intrahepatic Biliary Tract Carcinoma
C0221287|Carcinoma of Liver and Intrahepatic Biliary Tract
C0221287|Carcinoma of the Liver and Intrahepatic Biliary Tract
C0279607|hepatoma, adult primary
C0279607|adult primary hepatocellular carcinoma
C0279607|hepatocellular carcinoma, adult primary
C0279607|Adult Hepatocellular Carcinoma
C0279607|Adult Hepatoma
C0279607|Adult Liver Carcinoma
C0279607|Adult Primary Carcinoma of Liver Cell
C0279607|Adult Primary Carcinoma of the Liver Cell
C0279607|Adult Primary Hepatoma
C0279607|Adult Primary Liver Carcinoma
C0279607|Adult Primary Liver Cell Carcinoma
C2983709|Hepatocellular Carcinoma by AJCC v6 Stage
C2984092|Hepatocellular Carcinoma by AJCC v7 Stage
C3273019|Early Hepatocellular Carcinoma
C3273032|Lymphoepithelioma-Like Hepatocellular Carcinoma
C3273033|Well Differentiated Hepatocellular Carcinoma
C3273034|Moderately Differentiated Hepatocellular Carcinoma
C3273035|Poorly Differentiated Hepatocellular Carcinoma
C0345904|Liver, unspecified
C0345904|Malignant neoplasm of liver, unspecified
C0345904|malignant neoplasm of liver
C0345904|liver cancer
C0345904|liver cancer (diagnosis)
C0345904|liver neoplasm malignant
C0345904|malignant neoplasm of liver (diagnosis)
C0345904|Hepatic neoplasms malignant
C0345904|Cancer, Hepatic
C0345904|Cancers, Hepatic
C0345904|Hepatic Cancers
C0345904|Cancers, Liver
C0345904|Liver Cancers
C0345904|malignant tumor of liver
C0345904|Malignant neo liver NOS
C0345904|Malignant neoplasm of liver, not specified as primary or secondary
C0345904|hepatic cancer
C0345904|Cancer, Liver
C0345904|Malig neoplasm of liver, not specified as primary or sec
C0345904|Cancers, Hepatocellular
C0345904|Hepatocellular Cancers
C0345904|Malignant neoplasm of liver unspecified (disorder)
C0345904|Malignant tumor of liver (disorder)
C0345904|Malignant neoplasm of liver unspecified
C0345904|Malignant tumour of liver
C0345904|Liver--Cancer
C0345904|CANCER, HEPATOCELLULAR
C0345904|Hepatic neoplasm malignant NOS
C0345904|Malignant hepatic neoplasm
C0345904|Malignant liver tumor
C0345904|Hepatic tumour malignant
C0345904|Liver, cancer of
C0345904|Malignant liver tumour
C0345904|Hepatic neoplasm malignant
C0345904|Hepatic tumor malignant
C0345904|Hepatocellular Cancer
C0345904|Cancer of the Liver
C0345904|CA - Liver cancer
C0345904|Malignant neoplasm of liver (disorder)
C0345904|Malignant neoplasm of liver, NOS
C0345904|Cancer of Liver
C0345904|Neoplasm malig;liver
C0345904|malignant neosplasm of the liver
C0564703|Ca liver/biliary system NOS (disorder)
C0564703|Carcinoma liver/biliary system NOS
C0564703|Ca liver/biliary system
C0564703|Carcinoma liver/biliary system NOS (disorder)
C0564703|Ca liver/biliary system NOS
C0564703|carcinoma of liver and biliary system (diagnosis)
C0564703|neoplasm malignant carcinoma of liver and biliary system
C0564703|carcinoma of liver and biliary system
C0564703|Carcinoma liver/biliary system
C0564703|Carcinoma liver and/or biliary system (disorder)
C0564703|Carcinoma liver and/or biliary system
C0564703|Carcinoma liver/biliary system (disorder)
C2676033|HEPATOBLASTOMA CAUSED BY SOMATIC MUTATION
C1969388|hepatocellular carcinoma, somatic (diagnosis)
C1969388|hepatocellular carcinoma, somatic
C3898888|Hepatocellular Carcinoma Barcelona Clinic Liver Cancer Staging
C3898888|Hepatocellular Carcinoma by BCLC Stage
C3898888|BCLC Staging for Hepatocellular Carcinoma
C3898888|Hepatocellular Carcinoma by Barcelona Clinic Liver Cancer Stage
C3898888|Hepatocellular Carcinoma BCLC Staging
C3898888|Barcelona Clinic Liver Cancer Staging for Hepatocellular Carcinoma
C4030880|biopsy of liver showed carcinoma
C4030880|biopsy of liver showed carcinoma (procedure)
C4030854|biopsy of liver showed carcinoma primary
C4030854|biopsy of liver showed carcinoma primary (procedure)
C0744869|Metastatic hepatocellular carcinoma (morphologic abnormality)
C0744869|Metastatic hepatocellular carcinoma
C0348340|Other specified carcinomas of liver
C0348340|[X]Other specified carcinomas of liver
C0348340|Other specified carcinoma of liver
C0348340|Other specified carcinoma of liver (disorder)
C0348340|[X]Other specified carcinomas of liver (disorder)
C1391911|bile duct; carcinoma, with hepatocellular carcinoma
C1391911|carcinoma; bile duct, with hepatocellular carcinoma
C1391911|carcinoma; hepatocellular, with bile duct carcinoma
C1391911|hepatocellular; carcinoma, with bile duct carcinoma
C1391914|carcinoma; hepatocholangiolitic
C1391914|hepatocholangiolitic; carcinoma
C0206624|Hepatoblastoma
C0206624|Hepatoblastomas
C0206624|hepatoblastoma of liver
C0206624|hepatoblastoma of liver (diagnosis)
C0206624|Hepatoblastoma [Disease/Finding]
C0206624|HBL
C0206624|HEPATOBLASTOMA, MALIGNANT
C0206624|Pediatric Hepatoblastoma
C0206624|Pediatric Embryonal Hepatoma
C0206624|Hepatoblastoma NOS
C0206624|Embryonal hepatoma
C0206624|HBL - Hepatoblastoma
C0206624|Hepatoblastoma (clinical)
C0206624|Hepatoblastoma (disorder)
C0206624|Hepatoblastoma (morphologic abnormality)
C0206624|childhood hepatoblastoma
C0206624|hepatoblastoma, childhood
C0206624|embryonal; hepatoma
C0206624|hepatoma; embryonal
C1396365|embryoma; liver
C1396365|liver; embryoma
C1396366|embryoma; malignant, liver
C1396366|malignant; embryoma, liver
C1336811|Transplant-Related Hepatocellular Carcinoma
C1333067|Clear Cell Carcinoma of Liver Cells
C1333067|Clear Cell Carcinoma of the Liver Cells
C1333067|Clear Cell Hepatocellular Carcinoma
C1333067|Hepatocellular Clear Cell Carcinoma
C1333067|Liver Cell Clear Cell Carcinoma
C0279606|childhood hepatocellular carcinoma
C0279606|carcinoma, hepatocellular, childhood
C0279606|hepatocellular carcinoma, childhood
C0279606|pediatric hepatocellular carcinoma
C0279606|Childhood Hepatoma
C0279606|Childhood Liver Cell Carcinoma
C0279606|Pediatric Carcinoma of Liver Cell
C0279606|Pediatric Carcinoma of the Liver Cell
C0279606|Pediatric Hepatoma
C0279606|Pediatric Liver Cell Carcinoma
C0279606|Childhood Carcinoma of Liver Cell
C0279606|Childhood Carcinoma of the Liver Cell
C1112459|Liver cell carcinoma non-resectable
C1112459|Hepatocellular carcinoma non-resectable
C1112459|Non-Resectable Hepatocellular Carcinoma
C0861876|Liver carcinoma recurrent
C0861876|Carcinoma liver recurrent
C0861876|Hepatoma recurrent
C0861876|Hepatocellular carcinoma recurrent
C0861876|Liver cell carcinoma recurrent
C0861876|Malignant hepatoma recurrent
C0861876|Hepatocellular Carcinoma, Recurrent
C0861876|Recurrent Carcinoma of Liver Cell
C0861876|Recurrent Carcinoma of the Liver Cell
C0861876|Recurrent Hepatocellular Carcinoma
C0861876|Recurrent Hepatoma
C0861876|Recurrent Liver Cell Carcinoma
C0861876|Relapsed Carcinoma of Liver Cell
C0861876|Relapsed Carcinoma of the Liver Cell
C0861876|Relapsed Hepatocellular Carcinoma
C0861876|Relapsed Hepatoma
C0861876|Relapsed Liver Cell Carcinoma
C1332222|Aflatoxins-Related Hepatocellular Carcinoma
C1710014|Sarcomatoid Hepatocellular Carcinoma
C1710014|Sarcomatous Hepatocellular Carcinoma
C1709568|Pleomorphic Hepatocellular Carcinoma
C1266018|Sclerosing Hepatocellular Carcinoma
C1266018|Scirrhous Hepatocellular Carcinoma
C1266018|Hepatocellular carcinoma, scirrhous (morphologic abnormality)
C1266018|Hepatocellular carcinoma, scirrhous
C1266018|Sclerosing hepatic carcinoma
C1332228|Alcohol-Related Hepatocellular Carcinoma
C1333979|Hepatitis Virus Related Hepatocellular Carcinoma
C1333979|Hepatitis Virus-Related Hepatocellular Carcinoma
C0863194|Carcinoma liver resectable
C0863194|Liver cell carcinoma resectable
C0863194|Malignant hepatoma resectable
C0863194|Hepatoma resectable
C0863194|Liver carcinoma resectable
C0863194|Hepatocellular carcinoma resectable
C0863194|Hepatocellular Carcinoma, Resectable
C0863194|Resectable Carcinoma of Liver Cell
C0863194|Resectable Carcinoma of the Liver Cell
C0863194|Resectable Hepatocellular Carcinoma
C0863194|Resectable Hepatoma
C0863194|Resectable Liver Cell Carcinoma
C2111636|large cell carcinoma of liver with rhabdoid phenotype
C2111636|large cell carcinoma of liver with rhabdoid phenotype (diagnosis)
C2075624|liver neoplasm malignant clear cell type
C2075624|clear cell type neoplasm of liver (diagnosis)
C2075624|clear cell type neoplasm of liver
C2111730|large cell neuroendocrine carcinoma of liver
C2111730|large cell neuroendocrine carcinoma of liver (diagnosis)
