C2367785|hepatitis C genotype testing documented
C1533728|Hepatitis C virus genotype determination
C1148363|Hepatitis C virus genotype (finding)
C4272868|hepatitis c viral genotype
C3532919|Hepatitis C virus genotype 1
C3532920|Hepatitis C virus genotype 2
C3532921|Hepatitis C virus genotype 3
C3532922|Hepatitis C virus genotype 4
C3532923|Hepatitis C virus genotype 5
C3532924|Hepatitis C virus genotype 6
C3532919|HCV genotype 1
C3532920|HCV genotype 2
C3532921|HCV genotype 3
C3532922|HCV genotype 4
C3532923|HCV genotype 5
C3532924|HCV genotype 6
C3805156|Chronic hepatitis C virus genotype 1
C4049392|Chronic hepatitis C genotype 1
C4049393|Chronic hepatitis C genotype 1a
C4049394|Chronic hepatitis C genotype 1b
C4049395|Chronic hepatitis C genotype 2
C4049396|Chronic hepatitis C genotype 2a
C4049397|Chronic hepatitis C genotype 2b
C4049416|Chronic hepatitis C genotype 4i
C4049417|Chronic hepatitis C genotype 4j
C4049418|Chronic hepatitis C genotype 5
C4049419|Chronic hepatitis C genotype 5a
C4049420|Chronic hepatitis C genotype 6
C4049421|Chronic hepatitis C genotype 6a
C4049422|Chronic hepatitis C genotype 4c
C4049423|Chronic hepatitis C genotype 4d
C4049424|Chronic hepatitis C genotype 4e
C4049425|Chronic hepatitis C genotype 4f
C4049426|Chronic hepatitis C genotype 4g
C4049427|Chronic hepatitis C genotype 4h
C4049428|Chronic hepatitis C genotype 3d
C4049429|Chronic hepatitis C genotype 3e
C4049430|Chronic hepatitis C genotype 3f
C4049431|Chronic hepatitis C genotype 4
C4049432|Chronic hepatitis C genotype 4a
C4049433|Chronic hepatitis C genotype 2c
C4049434|Chronic hepatitis C genotype 2d
C4049435|Chronic hepatitis C genotype 3
C4049436|Chronic hepatitis C genotype 3a
C4049437|Chronic hepatitis C genotype 3b
C4049438|Chronic hepatitis C genotype 3c
C4049588|Chronic hepatitis C genotype 4b
C3805156|Chronic HCV genotype 1
C4049392|Chronic HCV genotype 1
C4049393|Chronic HCV genotype 1a
C4049394|Chronic HCV genotype 1b
C4049395|Chronic HCV genotype 2
C4049396|Chronic HCV genotype 2a
C4049397|Chronic HCV genotype 2b
C4049416|Chronic HCV genotype 4i
C4049417|Chronic HCV genotype 4j
C4049418|Chronic HCV genotype 5
C4049419|Chronic HCV genotype 5a
C4049420|Chronic HCV genotype 6
C4049421|Chronic HCV genotype 6a
C4049422|Chronic HCV genotype 4c
C4049423|Chronic HCV genotype 4d
C4049424|Chronic HCV genotype 4e
C4049425|Chronic HCV genotype 4f
C4049426|Chronic HCV genotype 4g
C4049427|Chronic HCV genotype 4h
C4049428|Chronic HCV genotype 3d
C4049429|Chronic HCV genotype 3e
C4049430|Chronic HCV genotype 3f
C4049431|Chronic HCV genotype 4
C4049432|Chronic HCV genotype 4a
C4049433|Chronic HCV genotype 2c
C4049434|Chronic HCV genotype 2d
C4049435|Chronic HCV genotype 3
C4049436|Chronic HCV genotype 3a
C4049437|Chronic HCV genotype 3b
C4049438|Chronic HCV genotype 3c
C4049588|Chronic HCV genotype 4b
C4272862|hepatitis c viral genotype 6
C4272863|hepatitis c viral genotype 5
C4272864|hepatitis c viral genotype 4
C4272865|hepatitis c viral genotype 3
C4272866|hepatitis c viral genotype 2
C4272867|hepatitis c viral genotype 1
C4272862|HCV viral genotype 6
C4272863|HCV viral genotype 5
C4272864|HCV viral genotype 4
C4272865|HCV viral genotype 3
C4272866|HCV viral genotype 2
C4272867|HCV viral genotype 1
C4284773|Hepatitis C virus genotype panel
C4284909|Hepatitis C virus genotype panel
C3655061|Hepatitis C virus resistance panel
C0973340|Infectious agent genotype analysis by nucleic acid (DNA or RNA); Hepatitis C virus
C1971440|Hepatitis C genotype testing documented as performed prior to initiation of antiviral treatment for Hepatitis C (HEP C)
C2030676|hepatitis C virus genotype analysis by nucleic acid
C4064267|probe and target amplification for hepatitis C virus genotype
C1742607|Reagents, Molecular Assay, Infection, Virus, Hepatitis C, Genotype
C3690224|IVD Test Reagent/Kits, Molecular Assay, Infection, Virus, Hepatitis C, Genotype
C4284773|HCV genotype panel
C4284909|HCV genotype panel
C3655061|HCV resistance panel
C0973340|Infectious agent HCV genotype analysis
C1971440|HCV genotype testing 
C2030676|HCV genotype analysis by nucleic acid
C4064267|HCV probe and target amplification
C1742607|HCV Molecular Assay
C3495939|Hepatitis C virus genotype 1a positive
C3495940|Hepatitis C virus genotype 1b positive
C3495941|Hepatitis C virus genotype 3a positive
C3495942|Hepatitis C virus genotype 3b positive
C3495943|Hepatitis C virus genotype 1 positive
C3495944|Hepatitis C virus genotype 3 positive
C3495939|HCV genotype 1a positive
C3495940|HCV genotype 1b positive
C3495941|HCV genotype 3a positive
C3495942|HCV genotype 3b positive
C3495943|HCV genotype 1 positive
C3495944|HCV genotype 3 positive
C3854557|Hepatitis C virus genotype 2b positive
C3854558|Hepatitis C virus genotype 2 positive
C3889043|Hepatitis C virus genotype 4 positive
C3889044|Hepatitis C virus genotype 5 positive
C3889045|Hepatitis C virus genotype 6 positive
C4049398|Hepatitis C virus genotype 6a positive
C4049399|Hepatitis C virus genotype 4f positive
C4049400|Hepatitis C virus genotype 4g positive
C4049401|Hepatitis C virus genotype 4h positive
C4049402|Hepatitis C virus genotype 4i positive
C4049403|Hepatitis C virus genotype 4j positive
C4049404|Hepatitis C virus genotype 5a positive
C4049405|Hepatitis C virus genotype 3f positive
C4049406|Hepatitis C virus genotype 4a positive
C4049407|Hepatitis C virus genotype 4b positive
C4049408|Hepatitis C virus genotype 4c positive
C4049409|Hepatitis C virus genotype 4d positive
C4049410|Hepatitis C virus genotype 4e positive
C4049411|Hepatitis C virus genotype 2a positive
C4049412|Hepatitis C virus genotype 2c positive
C4049413|Hepatitis C virus genotype 2d positive
C4049414|Hepatitis C virus genotype 3c positive
C4049415|Hepatitis C virus genotype 3e positive
C4049587|Hepatitis C virus genotype 3d positive
C1954138|Hepatitis C virus genotype
C1977372|Hepatitis C virus genotype
C4298651|Hepatitis C virus genotype 3
C4298652|Hepatitis C virus genotype 1
C4064283|probe with target amplification for hepatitis C virus genotype in serum or plasma
C1147970|Hepatitis C virus genotype
C1954139|Hepatitis C virus genotype
C4300371|Hepatitis C virus genotype 3 NS5a gene
C4300372|Hepatitis C virus genotype 1 NS5b gene
C4300373|Hepatitis C virus genotype 1 NS5a gene
C3654330|Hepatitis C virus NS5 gene mutations detected
C3654331|Hepatitis C virus NS3 gene mutations detected
C4285206|Hepatitis C virus genotype 1 NS5b gene mutations detected
C4285533|Hepatitis C virus genotype 3 NS5a gene mutations detected
C4296735|Hepatitis C virus genotype 3 NS5a gene mutations detected
C4296782|Hepatitis C virus genotype 1 NS5b gene mutations detected
C4296783|Hepatitis C virus genotype 1 NS5a gene mutations detected
C4298748|Hepatitis C virus genotype 1 NS5a gene mutations detected
C1269856|PCR positive for HCV viral RNA (genotype 1A)
C2367786|hepatitis C genotype testing performed prior to initiation of antiviral treatment
C2367786|hepatitis C genotype testing performed prior to initiation of antiviral treatment (treatment)
C2367786|hepatitis C genotype testing performed prior to initiation of antiviral treatment
C1148363|Hepatitis C virus genotype (finding)
C1148363|Hepatitis C virus genotype
C1533728|Hepatitis C virus genotype
C1533728|Hepatitis C virus genotype (procedure)
C1533728|HCV Genotyping
C1533728|Hepatitis C Virus Genotype Assay
C1533728|HCV Genotype Assay
C1533728|HCV Genotype Measurement
C1533728|HCV Genotype
C1533728|Hepatitis C virus genotype determination (procedure)
C1533728|Hepatitis C virus genotype determination
C4064267|probe with target amplification hepatitis c virus genotype
C4064267|probe with target amplification hepatitis c virus genotype (lab test)
C4064283|probe with target amplification for hepatitis C virus genotype in serum or plasma (lab test)
C4064283|probe with target amplification for hepatitis C virus genotype in serum or plasma
C4064283|probe & target amplif hepatitis c virus genotype serum / plasma
C3494966|Hepatitis C virus subtype 1a (organism)
C3494966|Hepatitis C virus subtype 1a
C3494965|Hepatitis C virus subtype 1b (organism)
C3494965|Hepatitis C virus subtype 1b
C3532925|Hepatitis C virus subtype 1c
C3532925|Hepatitis C virus subtype 1c (organism)
C3494964|Hepatitis C virus subtype 2a
C3494964|Hepatitis C virus subtype 2a (organism)
C3494963|Hepatitis C virus subtype 2b (organism)
C3494963|Hepatitis C virus subtype 2b
C3532926|Hepatitis C virus subtype 2c
C3532926|Hepatitis C virus subtype 2c (organism)
C3494962|Hepatitis C virus subtype 3a
C3494962|Hepatitis C virus subtype 3a (organism)
C3494961|Hepatitis C virus subtype 3b (organism)
C3494961|Hepatitis C virus subtype 3b
C3532918|Hepatitis C virus subtype 4a
C3532918|Hepatitis C virus subtype 4a (organism)
C3532927|Hepatitis C virus subtype 4b
C3532927|Hepatitis C virus subtype 4b (organism)
C3532928|Hepatitis C virus subtype 4c
C3532928|Hepatitis C virus subtype 4c (organism)
C3532929|Hepatitis C virus subtype 4d (organism)
C3532929|Hepatitis C virus subtype 4d
C3494960|Hepatitis C virus subtype 4e (organism)
C3494960|Hepatitis C virus subtype 4e
C3494959|Hepatitis C virus subtype 5a (organism)
C3494959|Hepatitis C virus subtype 5a
C3494958|Hepatitis C virus subtype 6a (organism)
C3494958|Hepatitis C virus subtype 6a
C3805156|Chronic hepatitis C virus genotype 1
C4049392|Chronic hepatitis C genotype 1
C4049393|Chronic hepatitis C genotype 1a
C4049394|Chronic hepatitis C genotype 1b
C4049395|Chronic hepatitis C genotype 2
C4049396|Chronic hepatitis C genotype 2a
C4049397|Chronic hepatitis C genotype 2b
C4049416|Chronic hepatitis C genotype 4i
C4049417|Chronic hepatitis C genotype 4j
C4049418|Chronic hepatitis C genotype 5
C4049419|Chronic hepatitis C genotype 5a
C4049420|Chronic hepatitis C genotype 6
C4049421|Chronic hepatitis C genotype 6a
C4049422|Chronic hepatitis C genotype 4c
C4049423|Chronic hepatitis C genotype 4d
C4049424|Chronic hepatitis C genotype 4e
C4049425|Chronic hepatitis C genotype 4f
C4049426|Chronic hepatitis C genotype 4g
C4049427|Chronic hepatitis C genotype 4h
C4049428|Chronic hepatitis C genotype 3d
C4049429|Chronic hepatitis C genotype 3e
C4049430|Chronic hepatitis C genotype 3f
C4049431|Chronic hepatitis C genotype 4
C4049432|Chronic hepatitis C genotype 4a
C4049433|Chronic hepatitis C genotype 2c
C4049434|Chronic hepatitis C genotype 2d
C4049435|Chronic hepatitis C genotype 3
C4049436|Chronic hepatitis C genotype 3a
C4049437|Chronic hepatitis C genotype 3b
C4049438|Chronic hepatitis C genotype 3c
C4049588|Chronic hepatitis C genotype 4b
C3655061|Hepatitis C virus resistance panel by Genotype method
C3655061|HCV resis panell Islt Genotyp
C3655061|Hepatitis C virus resistance panel:-:Point in time:Isolate:-:Genotyping
C3655061|Hepatitis C virus resistance panel:-:Pt:Isolate:-:Genotyping
C3655064|Boceprevir:Susc:Pt:Isolate:OrdQn:Genotyping
C3655064|Boceprevir [Susceptibility] by Genotype method
C3655064|Boceprevir Islt Genotyp
C3655064|Boceprevir:Susceptibility:Point in time:Isolate:Quantitative or Ordinal:Genotyping
C3655063|Telaprevir Islt Genotyp
C3655063|Telaprevir [Susceptibility] by Genotype method
C3655063|Telaprevir:Susc:Pt:Isolate:OrdQn:Genotyping
C3655063|Telaprevir:Susceptibility:Point in time:Isolate:Quantitative or Ordinal:Genotyping
C0973340|NFCT AGNT GENOTYP NUCLEIC ACID HEPATITIS C VIRUS
C0973340|Infectious agent genotype analysis by nucleic acid (DNA or RNA); Hepatitis C virus
C0973340|GENOTYPE DNA/RNA HEP C
C0973340|Analysis of infectious agent genotype of Hepatitis C virus
C1971440|Hepatitis C genotype testing documented as performed prior to initiation of antiviral treatment for Hepatitis C (HEP C)
C1971440|HEPC GN TSTNG DOCD B/4TXMNT
C1971440|HEPATITIS C GENOTYPE PRIOR ANTIVIRAL TREATMENT
C3495939|Hepatitis C virus genotype 1a positive
C3495940|Hepatitis C virus genotype 1b positive
C3495941|Hepatitis C virus genotype 3a positive
C3495942|Hepatitis C virus genotype 3b positive
C3495943|Hepatitis C virus genotype 1 positive
C3495944|Hepatitis C virus genotype 3 positive
C4049415|Hepatitis C virus genotype 3e positive
C3854557|Hepatitis C virus genotype 2b positive
C3854558|Hepatitis C virus genotype 2 positive
C3889043|Hepatitis C virus genotype 4 positive
C3889044|Hepatitis C virus genotype 5 positive
C3889045|Hepatitis C virus genotype 6 positive
C4049398|Hepatitis C virus genotype 6a positive
C4049399|Hepatitis C virus genotype 4f positive
C4049400|Hepatitis C virus genotype 4g positive
C4049401|Hepatitis C virus genotype 4h positive
C4049402|Hepatitis C virus genotype 4i positive
C4049403|Hepatitis C virus genotype 4j positive
C4049404|Hepatitis C virus genotype 5a positive
C4049405|Hepatitis C virus genotype 3f positive
C4049406|Hepatitis C virus genotype 4a positive
C4049407|Hepatitis C virus genotype 4b positive
C4049408|Hepatitis C virus genotype 4c positive
C4049409|Hepatitis C virus genotype 4d positive
C4049410|Hepatitis C virus genotype 4e positive
C4049411|Hepatitis C virus genotype 2a positive
C4049412|Hepatitis C virus genotype 2c positive
C4049413|Hepatitis C virus genotype 2d positive
C4049414|Hepatitis C virus genotype 3c positive
C4049587|Hepatitis C virus genotype 3d positive
C1954138|Hepatitis C virus genotype:Prid:Pt:Bld:Nom:Probe.amp.tar
C1954138|HCV Gentyp Bld PCR
C1954138|Hepatitis C virus genotype:Presence or Identity:Point in time:Whole blood:Nominal:DNA Nucleic Acid Probe.amp.tar
C1954138|Hepatitis C virus genotype [Identifier] in Blood by Probe and target amplification method
C1977372|Hepatitis C virus genotype:Prid:Pt:Tiss:Nom:Probe.amp.tar
C1977372|HCV Gentyp Tiss PCR
C1977372|Hepatitis C virus genotype:Presence or Identity:Point in time:Tissue, unspecified:Nominal:DNA Nucleic Acid Probe.amp.tar
C1977372|Hepatitis C virus genotype [Identifier] in Tissue by Probe and target amplification method
C1147970|Hepatitis C virus genotype:Prid:Pt:Ser/Plas:Nom:Probe.amp.tar
C1147970|HCV Gentyp SerPl PCR
C1147970|Hepatitis C virus genotype:Presence or Identity:Point in time:Serum/Plasma:Nominal:DNA Nucleic Acid Probe.amp.tar
C1147970|Hepatitis C virus genotype [Identifier] in Serum or Plasma by Probe and target amplification method
C1954139|Hepatitis C virus genotype:Prid:Pt:XXX:Nom:Probe.amp.tar
C1954139|HCV Gentyp XXX PCR
C1954139|Hepatitis C virus genotype:Presence or Identity:Point in time:To be specified in another part of the message:Nominal:DNA Nucleic Acid Probe.amp.tar
C1954139|Hepatitis C virus genotype [Identifier] in Unspecified specimen by Probe and target amplification method
C3654330|Hepatitis C virus NS5 gene mutations detected:Prid:Pt:Isolate:Nom:Genotyping
C3654330|Hepatitis C virus NS5 gene mutations detected:Presence or Identity:Point in time:Isolate:Nominal:Genotyping
C3654330|HCV NS5 Mut Det Islt Genotyp
C3654330|Hepatitis C virus NS5 gene mutations detected [Identifier] by Genotype method
C3654331|HCV NS3 Mut Det Islt Genotyp
C3654331|Hepatitis C virus NS3 gene mutations detected:Presence or Identity:Point in time:Isolate:Nominal:Genotyping
C3654331|Hepatitis C virus NS3 gene mutations detected:Prid:Pt:Isolate:Nom:Genotyping
C3654331|Hepatitis C virus NS3 gene mutations detected [Identifier] by Genotype method
