C0524662|Opiate Addiction
C0494376|Mental and behavioral disorders due to use of opioids, dependence syndrome
C0261864|Opiate antagonists causing adverse effects in therapeutic use
C0261817|Other opiates and related narcotics causing adverse effects in therapeutic use
C0747024|OPIATE ABUSE OPIUM
C0025605|Methadone
C2874436|Opioid dependence, uncomplicated
C2874436|opioid dependence uncomplicated
C2874436|opioid dependence uncomplicated (diagnosis)
C0338781|opioid dependence in remission (diagnosis)
C0338781|opioid dependence in remission
C0338781|Opioid dependence, in remission
C0338781|Opioid dependence in remission (disorder)
C2874441|Opioid dependence with intoxication
C2874441|Opioid dependence with intoxication, unspecified
C2874441|opioid dependence with intoxication (diagnosis)
C2874442|Opioid dependence with withdrawal
C2874442|opioid dependence with withdrawal (diagnosis)
C2874443|Opioid dependence with opioid-induced mood disorder
C2874443|opioid dependence with opioid-induced mood disorder (diagnosis)
C2874447|Opioid dependence with opioid-induced psychotic disorder
C2874447|Opioid dependence with opioid-induced psychotic disorder, unspecified
C2874447|Opioid dependence w opioid-induced psychotic disorder, unsp
C2874447|opioid dependence with opioid-induced psychotic disorder (diagnosis)
C2874448|Opioid dependence with other opioid-induced disorder
C2874451|Opioid dependence with unspecified opioid-induced disorder
C0338779|opioid dependence with continuous use (diagnosis)
C0338779|opioid dependence with continuous use
C0338779|Continuous opioid dependence
C0338779|Continuous opioid dependence (disorder)
C0338780|opioid dependence with episodic use
C0338780|opioid dependence with episodic use (diagnosis)
C0338780|Episodic opioid dependence
C0338780|Episodic opioid dependence (disorder)
C0338734|opioid dependence in combination with another drug (diagnosis)
C0338734|opioid dependence in combination with another drug
C0338734|Combined opioid with non-opioid drug dependence (disorder)
C0338734|Combined opioid with other drug dependence (disorder)
C0338734|Combined opioid with non-opioid drug dependence
C0338734|Combined opioid with other drug dependence, unspecified
C0338734|Combined opioid with other drug dependence, unspecified (disorder)
C0338734|Combined opioid with other drug dependence NOS
C0338734|Combined opioid with other drug dependence NOS (disorder)
C0338734|Combined opioid with other drug dependence
C3472691|Opioid dependence, on agonist therapy (disorder)
C3472691|Opioid dependence, on agonist therapy
C3472691|opioid dependence, on agonist therapy (diagnosis)
C0524662|Opioid dependence
C0524662|Dependence, Opiate
C0524662|Opiate Addiction
C0524662|opioid dependence (diagnosis)
C0524662|Addiction, Opiate
C0524662|Opioid dependence-unspec
C0524662|Opioid type dependence, unspecified use
C0524662|Opioid type dependence, unspecified
C0524662|[X]Drug addiction - opioids
C0524662|Unspecified opioid dependence
C0524662|Unspecified opioid dependence (disorder)
C0524662|Opioid type drug dependence
C0524662|Dependence on opiates
C0524662|Opioid type dependence
C0524662|Narcotism
C0524662|Opioid dependence (disorder)
C0524662|dependence; opiate
C0524662|dependence; opioids
C0524662|opioids; dependence
C0524662|Opiate Dependence
C3509112|opioid dependence with opioid-induced disorder
C3509112|opioid dependence with opioid-induced disorder (diagnosis)
C0338782|Opioid drug dependence NOS (disorder)
C0338782|Opioid drug dependence NOS
C0019337|Heroin Dependence
C0019337|Addiction, Heroin
C0019337|Dependence, Heroin
C0019337|Heroin Addiction
C0019337|Heroin Dependence [Disease/Finding]
C0019337|Addiction;drug(s);heroin
C0019337|[X]Heroin addiction
C0019337|Heroin dependence (diagnosis)
C0019337|opioid dependence heroin
C0019337|Heroin dependence (disorder)
C0019337|dependence; heroin
C0019337|heroin; dependence
C1960518|Fentanyl dependence (disorder)
C1960518|Fentanyl dependence
C1960518|Fentanyl dependence (diagnosis)
C1960518|opioid dependence fentanyl
C0026552|Morphine Dependence
C0026552|Addiction, Morphine
C0026552|Dependence, Morphine
C0026552|Morphine Addiction
C0026552|Morphine Dependence [Disease/Finding]
C0026552|opioid dependence morphine
C0026552|Morphine dependence (diagnosis)
C0026552|Morphine dependence (disorder)
C0026552|dependence; morphine
C0026552|morphine; dependence
C0026552|morphinism
C0338776|Methadone dependence
C0338776|opioid dependence methadone
C0338776|Methadone dependence (diagnosis)
C0338776|Methadone dependence (disorder)
C0338776|dependence; methadone
C0338776|methadone; dependence
C0338777|Opium dependence
C0338777|Opium dependence (diagnosis)
C0338777|opioid dependence opium
C0338777|Opium dependence (disorder)
C0338777|dependence; opium
C3840144|Buprenorphine dependence (disorder)
C3840144|Buprenorphine dependence
C0154478|Opioid dependence-contin
C0154478|Opioid type dependence, continuous
C0154478|Opioid type dependence, continuous use
C0154479|Opioid dependence-episod
C0154479|Opioid type dependence, episodic
C0154479|Opioid type dependence, episodic use
C0154480|Opioid dependence-remiss
C0154480|Opioid type dependence, in remission
C0494376|Mental and behavioral disorders due to use of opioids, dependence syndrome
C0494376|Mental and behavioural disorders due to use of opioids, dependence syndrome
C0494376|[X]Mental and behavioral disorders due to use of opioids: dependence syndrome
C0494376|[X]Mental and behavioral disorders due to use of opioids: dependence syndrome (disorder)
C0494376|[X]Mental and behavioural disorders due to use of opioids: dependence syndrome
C0494376|opiumism
C0865342|Opium alkaloids and their derivatives dependence
C1386557|codeine; dependence
C1386557|dependence; codeine
C1386560|dependence; dextromethorphan
C1386560|dextromethorphan; dependence
C1386561|dependence; dextromoramide
C1386561|dextromoramide; dependence
C1386562|dependence; dextrorphan
C1386562|dextrorphan; dependence
C1386566|dependence; ethylmorphine
C1386566|ethylmorphine; dependence
C1386570|dependence; drug, synthetic, with morphine-like effect
C1386577|dependence; laudanum
C1386577|laudanum; dependence
C1386588|dependence; methyl morphine
C1386588|methyl morphine; dependence
C1386594|dependence; paregoric
C1386594|paregoric; dependence
C1404354|morphinomania
C0261864|Adv eff opiat antagonist
C0261864|Opiate antagonists causing adverse effects in therapeutic use
C0868345|Levallorphan causing adverse effects in therapeutic use
C0868346|Nalorphine causing adverse effects in therapeutic use
C0868347|Naloxone causing adverse effects in therapeutic use
C0261817|Adv eff opiates
C0261817|Other opiates and related narcotics causing adverse effects in therapeutic use
C0868267|Codeine causing adverse effects in therapeutic use
C0868267|Methylmorphine causing adverse effects in therapeutic use
C0868268|Meperidine causing adverse effects in therapeutic use
C0868268|Pethidine causing adverse effects in therapeutic use
C0868269|Morphine causing adverse effects in therapeutic use
C0868270|Opium causing adverse effects in therapeutic use
C0868271|Opium alkaloids causing adverse effects in therapeutic use
C0025607|Methadyl Acetate
C0025607|methadylacetate
C0025607|Benzeneethanol, beta-(2-(dimethylamino)propyl)-alpha-ethyl-beta-phenyl-, acetate (ester)
C0025607|acetylmethadol
C0025607|Methadyl Acetate [Chemical/Ingredient]
C0025607|6-(Dimethylamino)-4,4-Diphenyl-3-Heptanol Acetate
C0057880|3-Hexanone, 4,4-diphenyl-6-(1-piperidinyl)-, hydrochloride, mixt. with 1-(diphenylmethyl)-4-methylpiperazine monohydrochloride
C0057880|diconal
C0058410|4,4-diphenyl-6-piperidino-3-heptanone
C0058410|dipipanone
C0058410|Phenylpiperone
C0058410|Dipipanone (product)
C0058410|Dipipanone (substance)
C0064006|6-(dimethylamino)-5-methyl-4,4-diphenyl-3-hexanone
C0064006|isomethadone
C0049312|5-methylmethadone
C0699057|Dolophine
C0699057|Roxane Brand of Methadone Hydrochloride
C0699058|Adanon
C0699059|Althose
C0699061|Amidone
C0699061|Amidine
C0699061|Amidone brand of methadone
C0260007|Phenadone
C0730805|Pinadone
C0730805|Pinewood Brand of Methadone Hydrochloride
C0788510|normethadone 10 MG/ML / oxilofrine 20 MG/ML Oral Solution
C0116497|erythro-5-methylmethadone
C0145747|threo-5-methylmethadone
C0592779|Methadose
C0592779|Mallinckrodt Brand of Methadone Hydrochloride
C0592779|Rosemont Brand of Methadone Hydrochloride
C0594373|Methex
C0594373|Generics Brand of Methadone Hydrochloride
C0025605|Methadone
C0025605|3-Heptanone, 6-(dimethylamino)-4,4-diphenyl-
C0025605|Methadone [Chemical/Ingredient]
C0025605|Methadone (product)
C0025605|Methadone (substance)
C0981584|Methadone Hydrochloride 5mg Oral tablet
C0981584|Methadone Hydrochloride, 5 mg oral tablet
C0981584|methadone 5 mg oral tablet
C0981584|METHADONE HCL 5MG EFFERVSC TAB
C0981584|METHADONE HCL 5MG TAB
C0981584|Methadone HCl Tab 5 MG
C0981584|METHADONE HYDROCHLORIDE 5 mg ORAL TABLET
C0981584|METHADONE HCL 5MG TAB [VA Product]
C0981584|METHADONE HCL 5MG TAB,EFFERVSC
C0981584|METHADONE HCL 5MG TAB,EFFERVSC [VA Product]
C0981584|methadone HCl 5 MG Oral Tablet
C0981584|Methadone hydrochloride 5mg tablet
C0981584|Methadone hydrochloride 5mg tablet (product)
C0981584|Methadone hydrochloride 5mg tablet (substance)
C0721688|Methadone Hydrochloride
C0721688|methadone hydrochloride (medication)
C0721688|Hydrochloride, Methadone
C0721688|Methadone Hydrochloride [Chemical/Ingredient]
C0721688|Methadone HCl [analgesic]
C0721688|Methadone HCl [cough] (product)
C0721688|Methadone HCl [analgesic] (product)
C0721688|Methadone HCl [cough]
C0721688|Methadone hydrochloride (substance)
C0721688|Methadone HCl [analgesic] (substance)
C0721688|Methadone HCl [cough] (substance)
C2093101|methadone hydrochloride (Dolophine) injection
C2093101|methadone hydrochloride injection
C2093101|methadone hydrochloride injection (medication)
C0806932|Methadone.long acting metabolite
C0806932|Long acting metabolite of methadone (substance)
C0806932|Long acting metabolite of methadone
C0033493|Propoxyphene
C0033493|D Propoxyphene
C0033493|Benzeneethanol, alpha-(2-(dimethylamino)-1-methylethyl)-alpha-phenyl-, propanoate (ester), (S-(R*,S*))-
C0033493|PROPOXYPHENE D
C0033493|Dextropropoxyphene
C0033493|Propoxyphene (product)
C0033493|Dextropropoxyphene (product)
C0033493|synthetic narcotics propoxyphene preparations
C0033493|propoxyphene preparations (medication)
C0033493|propoxyphene preparations
C0033493|D-Propoxyphene
C0033493|Dextropropoxyphene [Chemical/Ingredient]
C0033493|4-Dimethylamino-3-methyl-1,2-diphenyl-2-propoxybutane
C0033493|Propoxyphene (substance)
C0033493|Dextropropoxyphene (substance)
C1992369|Methadone &#x7C; bld-ser-plas
C1992375|Methadone &#x7C; stool
C1992378|Methadone &#x7C; XXX
C1992373|Methadone &#x7C; meconium
C1626306|Methadone+Metabolite
C1992383|Methadone.R &#x7C; bld-ser-plas
C1992377|Methadone &#x7C; vitreous fluid
C1992374|Methadone &#x7C; milk
C1992368|Methadone &#124; bile fluid
C1992368|Methadone &#x7C; bile fluid
C3534187|Methadone &#x7C; Saliva
C0366544|Methadone Dose
C0366544|Methadone:Mass:Pt:Dose:Qn
C0366544|Methadone [Mass] of Dose
C0366544|Methadone:Mass:Point in time:Dose med or substance:Quantitative
C1992376|Methadone &#x7C; urine
C0046103|1,5-dimethyl-3,3-diphenyl-2-ethylidenepyrrolidine
C0046103|2-ethylidene-1,5-dimethyl-3,3-diphenylpyrrolidine
C0046103|EDPP
C0046103|2-Et-1,5-diMe-3,3-DPP
C0046103|EDDP-3,3
C1992371|Methadone &#x7C; gastric fluid
C1992372|Methadone &#x7C; hair
C0628179|6-dimethylamino-4-(4-hydroxyphenyl)-4-phenylheptan-3-one
C0628179|para-hydroxymethadone
C0624343|2-formamido-4,4-diphenyl-5-heptanone
C0624343|FADPH
C0069008|6-dimethylamino-4,4-diphenylhexan-3-one
C0069008|nor-methadone
C0069008|normethadone
C0360477|Oral methadone
C0360477|Methadone Oral Product
C0360477|Oral form methadone (product)
C0360477|Oral form methadone
C0360477|Oral methadone (product)
C0360477|Oral methadone (substance)
C0360478|Parenteral methadone
C0360478|Parenteral form methadone (product)
C0360478|Parenteral form methadone
C0360478|Parenteral methadone (product)
C0360478|Parenteral methadone (substance)
C0684217|Physeptone
C0684217|Martindale Brand of Methadone Hydrochloride
C0684217|Phymet
C0684217|GlaxoSmithKline Brand of Methadone Hydrochloride
C1563840|Biomet Brand of Methadone Hydrochloride
C1563840|Biodone
C1563841|Pharmascience Brand of Methadone Hydrochloride
C1563841|Metadol
C1563842|Esteve Brand of Methadone Hydrochloride
C1563842|Metasedin
C1563843|addiCare Brand of Methadone Hydrochloride
C1563843|Methaddict
C1563844|Yamanouchi Brand of Methadone Hydrochloride
C1563844|Symoron
C0731186|Martindale Methadone DTF
