C0004096|Asthma
C0340067|drug-induced asthma (diagnosis)
C0340067|asthma drug-induced
C0340067|drug-induced asthma
C0340067|Drug-induced asthma (disorder)
C0340067|Drug-induced asthma, NOS
C0348819|Mixed asthma
C0348819|asthma mixed
C0348819|mixed asthma (diagnosis)
C0348819|Mixed asthma (disorder)
C0348819|asthma; mixed
C0348819|mixed; asthma
C0858626|Asthmatic attack induced
C0856716|Aspirin-sensitive asthma
C0856716|Aspirin asthma
C0856716|Asthma aspirin-sensitive
C0859194|Chronic obstructive asthma (with obstructive pulmonary disease), w/o-ment of status asthmaticus
C0859194|Chronic obstructive asthma (with obstructive pulmonary disease), w/o ment of status asthmaticus
C0494660|Predominantly allergic asthma
C0494660|allergic (predominantly) asthma
C0494660|asthma; predominantly allergic
C0494660|predominantly allergic; asthma
C0236072|Bronchospasm paradoxical
C0236072|Paradoxical bronchospasm
C0236072|Paradoxical bronchospasm (finding)
C0155883|Chronic obstructive asthma
C0155883|chronic obstructive asthma (diagnosis)
C0155883|Chronic obstructive asthma (with obstructive pulmonary disease)
C0948683|Asthmatic attack atopic
C0155879|extrinsic asthma with status asthmaticus
C0155879|extrinsic asthma with status asthmaticus (diagnosis)
C0155879|Ext asthma w status asth
C0155879|Extrinsic asthma with status asthmaticus (disorder)
C0155880|Nonallergic asthma
C0155880|Intrinsic asthma
C0155880|intrinsic asthma (diagnosis)
C0155880|intrinsic nonallergic asthma
C0155880|Intrinsic asthma (disorder)
C0155880|Intrinsic asthma NOS
C0155880|Intrinsic asthma NOS (disorder)
C0155880|Non-allergic asthma
C0155880|Non-allergic asthma (diagnosis)
C0155880|asthma non-allergic
C0155880|Asthma due to internal immunological process
C0155880|Non-allergic asthma (disorder)
C0155880|asthma; intrinsic, nonallergic
C0155880|asthma; intrinsic
C0155880|asthma; nonallergic
C0155880|intrinsic; asthma, nonallergic
C0155880|intrinsic; asthma
C0155880|nonallergic; asthma
C0155880|Intrinsic asthma (disorder) [Ambiguous]
C0155882|intrinsic asthma with status asthmaticus (diagnosis)
C0155882|intrinsic asthma with status asthmaticus
C0155882|Int asthma w status asth
C0155882|Intrinsic asthma with status asthmaticus (disorder)
C0155878|Extrinsic asthma without mention of status asthmaticus
C0155878|Extrinsic asthma NOS
C0155878|Extrinsic asthma, unspecified
C0155881|Intrinsic asthma without mention of status asthmaticus
C0155881|Intrinsic asthma NOS
C0155881|Intrinsic asthma, unspecified
C0155886|Asthma, unspecified type, without mention of status asthmaticus
C0155886|Asthma NOS
C0155886|Asthma, unspecified type, unspecified
C0549336|Asthma aggravated
C0347950|Asthma attack
C0347950|Asthma attack NOS (disorder)
C0347950|Asthma attack (& NOS) (disorder)
C0347950|Asthma attack (& NOS)
C0347950|Asthma attack NOS
C0347950|asthma attack (diagnosis)
C0347950|Asthma attack (disorder)
C0347950|Acute exacerbation of asthma
C0347950|Acute exacerbation of asthma (disorder)
C0347950|Asthmatic attack
C0810292|Other and unspecified asthma
C0004096|Asthma
C0004096|Asthmas
C0004096|Asthma, unspecified
C0004096|Bronchial asthma
C0004096|asthma (diagnosis)
C0004096|Br. asthma
C0004096|Asthma NOS
C0004096|Unspecified asthma
C0004096|Asthma [Disease/Finding]
C0004096|Asthma, Bronchial
C0004096|Asthma (disorder)
C0004096|Asthma unspecified (disorder)
C0004096|Asthma NOS (disorder)
C0004096|Asthma unspecified
C0004096|-- Asthma
C0004096|Asthmatic
C0004096|Asthma bronchial
C0004096|Bronchitic asthma
C0004096|Cardio/pulm: Asthma
C0004096|Airway hyperreactivity
C0004096|Asthma, NOS
C0004096|Bronchial asthma, NOS
C0004096|Asthma (disorder) [Ambiguous]
C0038218|Asthmatic Crises
C0038218|Asthmatic Shocks
C0038218|Asthmaticus, Status
C0038218|Crises, Asthmatic
C0038218|Crisis, Asthmatic
C0038218|Shock, Asthmatic
C0038218|Shocks, Asthmatic
C0038218|Status Asthmaticus
C0038218|Status asthmaticus -RETIRED-
C0038218|Asthma w status asthmat
C0038218|Asthmatic Shock
C0038218|Status Asthmaticus [Disease/Finding]
C0038218|Asthmatic Crisis
C0038218|Status asthmaticus NOS
C0038218|(Severe asthma attack) or (status asthmaticus NOS)
C0038218|Status asthmaticus NOS (disorder)
C0038218|Status asthmaticus (disorder)
C0038218|Severe asthma attack
C0038218|(Severe asthma attack) or (status asthmaticus NOS) (disorder)
C0038218|Acute severe asthma
C0038218|Asthma with status asthmaticus
C0038218|Acute severe exacerbation of asthma
C0038218|Asthma with status asthmaticus (disorder)
C0038218|Acute severe exacerbation of asthma (disorder)
C0038218|Asthma, unspecified type, with status asthmaticus
C0038218|asthma with status asthmaticus (diagnosis)
C0038218|asthmaticus; status
C0038218|status; asthmaticus
C0004099|Asthma, Exercise Induced
C0004099|Asthma, Exercise-Induced
C0004099|Asthmas, Exercise-Induced
C0004099|Exercise Induced Asthma
C0004099|Exercise-Induced Asthmas
C0004099|EXERCISE IND ASTHMA
C0004099|ASTHMA EXERCISE IND
C0004099|exercise-induced asthma
C0004099|exercise-induced asthma (diagnosis)
C0004099|EIA (exercise-induced asthma)
C0004099|Asthma exercise induced
C0004099|Asthma, Exercise-Induced [Disease/Finding]
C0004099|Exercise-induced asthma (finding)
C0004099|EIA - Exercise-induced asthma
C0004099|Exercise-induced asthma (disorder)
C1319853|Aspirin Induced Asthmas
C1319853|Aspirin-Induced Asthmas
C1319853|NSAID-induced Asthmas
C1319853|Aspirin-Induced Asthma Syndromes
C1319853|Asthma Syndrome, Aspirin-Induced
C1319853|Asthma, NSAID induced
C1319853|Syndrome, Aspirin-Induced Asthma
C1319853|Syndromes, Aspirin-Induced Asthma
C1319853|Asthmas, Aspirin-Induced
C1319853|Asthma, Aspirin Induced
C1319853|Asthma Syndromes, Aspirin-Induced
C1319853|Asthmas, Aspirin Induced
C1319853|Induced Asthmas, Aspirin
C1319853|Asthma, Aspirin-Induced
C1319853|Asthmas, NSAID-induced
C1319853|NSAID-induced Asthma
C1319853|Aspirin Induced Asthma Syndrome
C1319853|Induced Asthma, Aspirin
C1319853|Asthma, NSAID-induced
C1319853|Asthma, Aspirin-Induced [Disease/Finding]
C1319853|Aspirin Induced Asthma
C1319853|Aspirin-Induced Asthma
C1319853|Aspirin-Induced Asthma Syndrome
C1319853|Aspirin-induced asthma (diagnosis)
C1319853|asthma drug-induced aspirin
C1319853|Aspirin-induced asthma (disorder)
C1960045|Mild intermittent asthma
C1960045|Mild intermittent asthma (disorder)
C1960045|mild intermittent asthma (diagnosis)
C1960045|Mild intermittent asthma NOS
C1960046|Mild persistent asthma (disorder)
C1960046|Mild persistent asthma
C1960046|mild persistent asthma (diagnosis)
C1960046|Mild persistent asthma NOS
C1960047|Moderate persistent asthma
C1960047|Moderate persistent asthma (disorder)
C1960047|moderate persistent asthma (diagnosis)
C1960047|Moderate persistent asthma NOS
C1960048|Severe persistent asthma (disorder)
C1960048|Severe persistent asthma
C1960048|severe persistent asthma (diagnosis)
C1960048|Severe persistent asthma NOS
C2887463|Unspecified asthma with (acute) exacerbation
C2887464|Unspecified asthma with status asthmaticus
C2887465|Unspecified asthma, uncomplicated
C2919352|Seasonal asthma (disorder)
C2919352|Seasonal asthma
C2919352|Seasonal asthma (diagnosis)
C2919352|asthma seasonal
C0349790|asthma with acute exacerbation
C0349790|asthma with acute exacerbation (diagnosis)
C0349790|Exacerbation of asthma (disorder)
C0349790|Exacerbation of asthma
C0349790|Acute exacerbation of asthma
C0694548|cough variant asthma
C0694548|cough variant asthma (diagnosis)
C0694548|Cough variant asthma (disorder)
C0264408|childhood asthma (diagnosis)
C0264408|childhood asthma
C0264408|Childhood asthma NOS
C0264408|Asthma in Children
C0264408|Childhood asthma (disorder)
C0264408|asthma; childhood
C0264408|childhood; asthma
C0264408|Asthma, childhood
C1740754|INTERMITTENT ASTHMA
C1740754|Intermittent asthma (Asthma)
C1740754|Intermittent asthma (disorder)
C1740754|intermittent asthma (diagnosis)
C0264423|occupational asthma (diagnosis)
C0264423|occupational asthma
C0264423|Asthmas, Occupational
C0264423|Asthma, Occupational
C0264423|Occupational Asthmas
C0264423|Asthma, Occupational [Disease/Finding]
C0264423|Industrial asthma
C0264423|Occupational asthma (disorder)
C0155877|Allergic asthma
C0155877|extrinsic asthma
C0155877|extrinsic asthma (diagnosis)
C0155877|atopic asthma
C0155877|extrinsic allergic asthma
C0155877|Extrinsic asthma (disorder)
C0155877|Extrinsic asthma NOS (disorder)
C0155877|Allergic atopic asthma (disorder)
C0155877|Allergic atopic asthma
C0155877|Extrinsic asthma NOS
C0155877|Allergic asthma (disorder)
C0155877|asthma allergic
C0155877|Allergic asthma (diagnosis)
C0155877|ASTHMA, ATOPIC
C0155877|Asthma extrinsic
C0155877|asthma; allergic extrinsic
C0155877|asthma; atopic
C0155877|asthma; extrinsic
C0155877|atopic; asthma
C0155877|extrinsic; asthma
C0155877|allergic; asthma, extrinsic
C0155877|allergic; extrinsic asthma
C0155877|Extrinsic asthma [Ambiguous] (disorder)
C0155877|Allergic atopic asthma [Ambiguous]
C0155877|Asthma, allergic NOS
C0264413|Asthma late onset
C0264413|Late onset asthma
C0264413|LOA - late onset asthma
C0264413|Late onset asthma (disorder)
C0264413|Late-onset asthma
C0264413|Late-onset asthma (LOA)
C0264413|asthma late-onset
C0264413|Late-onset asthma (diagnosis)
C0264413|asthma; late onset
C0264413|late onset; asthma
C0729337|asthma brittle
C0729337|asthma brittle (diagnosis)
C0729337|Brittle asthma
C0729337|Brittle asthma (disorder)
C3508931|asthma uncomplicated
C3508931|asthma uncomplicated (diagnosis)
C3508931|Uncomplicated asthma (disorder)
C3508931|Uncomplicated asthma
C0264508|Asthmatic pulmonary alveolitis
C0264508|Asthmatic pulmonary alveolitis (disorder)
C0264411|hay fever with asthma
C0264411|Extrinsic asthma - atopy
C0264411|Hay asthma (disorder)
C0264411|Pollen asthma
C0264411|Extrinsic (atopic) asthma
C0264411|Hay asthma
C0264411|hay fever with asthma (diagnosis)
C0264411|Hay fever with asthma (disorder)
C0264411|asthma; hay fever
C0264411|hay fever; asthma
C0264411|Asthma, hay
C0264451|Weavers' cough
C0264451|weavers' cough (diagnosis)
C0264451|Weavers' cough (disorder)
C0264417|Canine allergic bronchitis
C0264417|Canine allergic bronchitis (disorder)
C0684913|chemical-induced asthma
C0684913|asthma chemical-induced
C0684913|chemical-induced asthma (diagnosis)
C0684913|Chemical-induced asthma (disorder)
C0684913|Chemical-induced asthma, NOS
C1956414|Cardiac asthma
C1956414|Asthma, Cardiac
C1956414|Asthma - cardiac
C1956414|Asthma cardiac
C1956414|Cardiac asthma (disorder)
C1956414|asthma; cardiac
C1956414|cardiac; asthma
C0264404|Chronic allergic bronchitis (diagnosis)
C0264404|Chronic allergic bronchitis
C0264404|allergic bronchitis chronic
C0264404|Chronic allergic bronchitis (disorder)
C0340070|millers' asthma
C0340070|millers' asthma (diagnosis)
C0340070|asthma millers'
C0340070|Mill-workers' asthma
C0340070|Millers' cough
C0340070|Grain worker's asthma
C0340070|Millers' asthma (disorder)
C0006542|Byssinoses
C0006542|Byssinosis
C0006542|Mill fever
C0006542|cotton dust asthma
C0006542|brown lung
C0006542|cotton mill fever
C0006542|byssinosis (diagnosis)
C0006542|occupational asthma (byssinosis)
C0006542|Brown Lungs
C0006542|Brown Lung Diseases
C0006542|Byssinosis [Disease/Finding]
C0006542|Brown Lung Disease
C0006542|Mill fever (disorder)
C0006542|Cotton workers' lung disease
C0006542|Cotton-dust asthma
C0006542|Byssinosis (disorder)
C0006542|disease (or disorder); respiratory tract, due to cotton dust
C0006542|fibrosis; lung, with byssinosis
C0006542|lung; fibrosis, with byssinosis
C1563057|Work aggravated asthma
C1563057|Work aggravated asthma (disorder)
C1260881|Allergic bronchitis
C1260881|allergic bronchitis (diagnosis)
C1260881|Bronchitis;allergic
C1260881|allergic bronchitis NOS
C1260881|Feline asthma
C1260881|Feline allergic bronchitis
C1260881|Feline allergic bronchitis (disorder)
C1260881|Allergic bronchitis (disorder)
C1260881|Allergic bronchitis, NOS
C1260881|Bronchitis, allergic
C0264449|Pneumonopathy due to inhalation of dust (disorder)
C0264449|Pneumonopathy due to inhalation of dust
C0264449|Pneumonopathy due to inhalation of dust, NOS
C1319018|asthmatic bronchitis
C1319018|asthmatic bronchitis (diagnosis)
C1319018|Asthma/bronchitis
C1319018|Asthmatic bronchitis NOS
C1319018|Bronchitis;asthmatic
C1319018|Bronchitis;wheezy
C1319018|Asthmatic bronchitis (disorder)
C1319018|Wheezy bronchitis
C1319018|Bronchitis asthmatic
C1319018|Asthmatic bronchitis, NOS
C1319018|Bronchitis, asthmatic
C0032318|Pneumonopathy due to inhalation of other dust
C0032318|Pneumopathy due to inhalation of other dust
C0032318|Dust pneumonopathy NEC
C0032318|Pneumopathy due to inhalation of other dust NOS (disorder)
C0032318|Pneumopathy due to inhalation of other dust (disorder)
C0032318|Pneumopathy due to inhalation of other dust NOS
C3266628|Persistent asthma
C3266628|Persistent asthma (disorder)
C3266628|Persistent asthma (diagnosis)
C3266628|asthma persistent
C3662842|Chronic obstructive airway disease with asthma (disorder)
C3662842|Chronic obstructive airway disease with asthma
C3661951|Asthma with irreversible airway obstruction
C3661951|Asthma with irreversible airway obstruction (disorder)
C0582415|asthma acute
C0582415|Acute asthma
C0582415|Acute asthma (diagnosis)
C0582415|Acute asthma (disorder)
C0582415|asthma; acute
C0582415|acute; asthma
C1828277|Substance induced asthma
C1828277|Substance induced asthma (disorder)
C1828277|substance-induced asthma
C1828277|asthma substance-induced
C1828277|substance-induced asthma (diagnosis)
C0581124|Mild asthma (finding)
C0581124|Mild asthma (disorder)
C0581124|Mild asthma
C0581124|Mild asthma (procedure)
C0581124|asthma mild
C0581124|Mild asthma (diagnosis)
C0581123|Occasional asthma (finding)
C0581123|Occasional asthma (disorder)
C0581123|Occasional asthma
C0581123|Occasional asthma (procedure)
C0581123|asthma occasional
C0581123|Occasional asthma (diagnosis)
C0264405|Asthma without status asthmaticus (diagnosis)
C0264405|Asthma without status asthmaticus
C0264405|Asthma without status asthmaticus (disorder)
C0581125|Moderate asthma (finding)
C0581125|Moderate asthma (disorder)
C0581125|Moderate asthma
C0581125|Moderate asthma (procedure)
C0581125|asthma moderate
C0581125|Moderate asthma (diagnosis)
C0340073|Factitious asthma
C0340073|asthma factitious
C0340073|Factitious asthma (diagnosis)
C0340073|Emotional laryngeal wheezing
C0340073|Functional laryngeal stridor
C0340073|Factitious asthma (disorder)
C0581126|Severe asthma (finding)
C0581126|Severe asthma (disorder)
C0581126|Severe asthma (procedure)
C0581126|Severe asthma
C0581126|asthma severe
C0581126|Severe asthma (diagnosis)
C0581126|asthma; severe
C0581126|severe; asthma
C1859647|ASTHMA, SHORT STATURE, AND ELEVATED IgA
C1853964|DERMATITIS, ATOPIC, 3
C1853964|ATOD3
C1853964|Dermatitis, Atopic, with Asthma
C3280315|PAFAD
C3280315|PLATELET-ACTIVATING FACTOR ACETYLHYDROLASE DEFICIENCY
C1858067|ASTHMA AND NASAL POLYPS
C1869116|ASTHMA, SUSCEPTIBILITY TO
C1869116|ASTHMA, SUSCEPTIBILITY TO (finding)
C1869116|asthma susceptibility
C1869116|asthma susceptibility (diagnosis)
C1869116|ASTHMA-RELATED TRAITS, SUSCEPTIBILITY TO
C1869116|ASTHMA, BRONCHIAL
C3838502|asthma protection (diagnosis)
C3838502|asthma protection
C3838894|Asthma in mother complicating childbirth (disorder)
C3838894|Asthma in childbirth
C3838894|Asthma in mother complicating childbirth
C4038730|Asthma-chronic obstructive pulmonary disease overlap syndrome
C4038730|Asthma-chronic obstructive pulmonary disease overlap syndrome (disorder)
C4038730|Asthma-COPD overlap syndrome (ACOS)
C4038730|Asthma-COPD overlap syndrome
C0741267|Steroid dependent asthma
C0741267|Steroid dependent asthma (disorder)
C1388871|asthma; croup
C1388871|croup; asthma
C1388880|asthmatic; dyspnea
C1388880|dyspnea; asthmatic
C1388882|asthmatic; dyspnea, with bronchitis
C1388882|dyspnea; asthmatic, with bronchitis
C1403212|obstruction; airway, with asthma
C1403212|airway; obstruction, with asthma
C1260416|Other forms of asthma
C1176342|Asthma NOS w (ac) exac
C1176342|Asthma, unspecified type, with (acute) exacerbation
