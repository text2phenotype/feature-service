C2062763|benzodiazepine abuse
C2878161|underdosing of benzodiazepines
C0418282|Intentional benzodiazepine overdose
C2878162|Underdosing of benzodiazepines, initial encounter
C2878163|Underdosing of benzodiazepines, subsequent encounter
C2878164|Underdosing of benzodiazepines, sequela
C0747951|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE
C0747952|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE DEPENDENCE
C0747953|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE POTENTIAL
C0747954|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE REMISSION
C0747955|PRESCRIPTION DRUG ABUSE BENZODIAZEPINE WITHDRAWAL
C2104566|continuous benzodiazepine abuse (diagnosis)
C2104566|continuous benzodiazepine abuse
C2104567|episodic benzodiazepine abuse (diagnosis)
C2104567|episodic benzodiazepine abuse
C2104568|benzodiazepine abuse in remission (diagnosis)
C2104568|benzodiazepine abuse in remission
C2878162|Underdosing of benzodiazepines, initial encounter
C2878163|Underdosing of benzodiazepines, subsequent encounter
C2878164|Underdosing of benzodiazepines, sequela
C0572936|Intentional flunitrazepam overdose
C0572936|Intentional flunitrazepam overdose (disorder)
C0572989|Intentional prazepam overdose
C0572989|Intentional prazepam overdose (disorder)
C0572977|Intentional ketazolam overdose
C0572977|Intentional ketazolam overdose (disorder)
C0572950|Intentional nitrazepam overdose
C0572950|Intentional nitrazepam overdose (disorder)
C0572969|Intentional clobazam overdose
C0572969|Intentional clobazam overdose (disorder)
C0572962|Intentional bromazepam overdose
C0572962|Intentional bromazepam overdose (disorder)
C0572939|Intentional flurazepam overdose
C0572939|Intentional flurazepam overdose (disorder)
C0572947|Intentional lormetazepam overdose
C0572947|Intentional lormetazepam overdose (disorder)
C0572943|Intentional loprazolam overdose
C0572943|Intentional loprazolam overdose (disorder)
C0572981|Intentional medazepam overdose
C0572981|Intentional medazepam overdose (disorder)
C0418284|Intentional chlordiazepoxide overdose (disorder)
C0418284|Deliberate overdose of chlordiazepoxide
C0418284|Intentional chlordiazepoxide overdose
C0418284|Deliberate overdose of chlordiazepoxide (disorder)
C0572993|Intentional midazolam overdose
C0572993|Intentional midazolam overdose (disorder)
C0418283|self-inflicted overdose of diazepam
C0418283|self-inflicted overdose of diazepam (diagnosis)
C0418283|toxicity from diazepam due to a self-inflicted overdose
C0418283|Intentional diazepam overdose
C0418283|Deliberate overdose of diazepam (disorder)
C0418283|Deliberate overdose of diazepam
C0418283|Intentional diazepam overdose (disorder)
C0418285|Deliberate overdose of temazepam (disorder)
C0418285|Intentional temazepam overdose (disorder)
C0418285|Intentional temazepam overdose
C0418285|Deliberate overdose of temazepam
C0572954|Intentional triazolam overdose
C0572954|Intentional triazolam overdose (disorder)
C0572958|Intentional alprazolam overdose
C0572958|Intentional alprazolam overdose (disorder)
C0572973|Intentional potassium clorazepate overdose
C0572973|Intentional potassium clorazepate overdose (disorder)
C0572973|Intentional dipotassium clorazepate overdose
C0572985|Intentional oxazepam overdose
C0572985|Intentional oxazepam overdose (disorder)
C0573000|Intentional lorazepam overdose
C0573000|Intentional lorazepam overdose (disorder)
C0572892|Intentional clonazepam overdose
C0572892|Intentional clonazepam overdose (disorder)
