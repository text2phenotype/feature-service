C0027415|Narcotics
C0202273|Drug of abuse, quantitative screen, includes amphetamines, barbiturates, benzodiazepines, cannabinoids, cocaine, methadone, methaqualone, opiates, phencyclidines and propoxyphene
C0086190|Illicit Drugs
C2911101|Drug abuse counseling and surveillance of drug abuser
C0202273|Drug of abuse, quantitative screen, includes amphetamines, barbiturates, benzodiazepines, cannabinoids, cocaine, methadone, methaqualone, opiates, phencyclidines and propoxyphene
C0221793|opiate alkaloid
C0221793|Alkaloids, Opiate
C0221793|Opiate Alkaloids
C0221793|Opiate Alkaloids [Chemical/Ingredient]
C0221793|Opium alkaloid
C0221793|Opium alkaloid (product)
C0221793|Opium alkaloid (substance)
C0221793|Opium Alkaloids
C0025605|Methadone
C0025605|3-Heptanone, 6-(dimethylamino)-4,4-diphenyl-
C0025605|Methadone [Chemical/Ingredient]
C0025605|Methadone (product)
C0025605|Methadone (substance)
C0030350|Papaverine
C0030350|Isoquinoline, 1-((3,4-dimethoxyphenyl)methyl)-6,7-dimethoxy-
C0030350|Papaverine [Chemical/Ingredient]
C0030350|Papaverine (substance)
C0030350|Papaverine (product)
C0030350|PAP
C0728935|K 315
C0728935|K315
C0728935|K-315
C0205752|Endogenous Opioids
C0205752|endogenous opiate
C0205752|Endogenous Opiates
C0205752|endorphin
C0205752|endogenous opioid
C0205752|Opioids (Endogenous)
C0205752|Opiates, Endogenous
C0596008|Levorphanol Tartrate
C0596008|Tartrate, Levorphanol
C0596008|l-3-Hydroxy-N-methylmorphinan Bitartrate
C0596008|2H-10,4a-Iminoethanophenanthren-6-ol, 1,3,4,9,10,10a-hexahydro-11-methyl-, Tartrate
C0596008|Lemoran
C0596008|Morphinan-3-ol, 17-methyl-, Tartrate(1:1)(Salt)
C0596008|Morphinan-3-ol, 17-methyl-,(2R,3R)-2,3-dihydroxybutanedioate(1:1)
C0596008|NIH 4590
C0596008|Ro 1-5431/7
C0596008|levorphanol tartrate (medication)
C0596008|synthetic narcotics levorphanol tartrate
C0596008|Levorphanol Tartrate [Chemical/Ingredient]
C0596008|Levorphanol tartrate [anaesth]
C0596008|Levorphanol tartrate [anesth]
C0596008|Levorphanol tartrate (substance)
C0596008|Levorphanol tartrate [anesth] (product)
C0596008|Levorphan tartrate
C0596008|Levorphanol tartrate [anesth] (substance)
C0596008|Levorphanol tartrate [dup] (substance)
C0376196|Opiates
C0376196|opiate
C0376196|Opiate (product)
C0376196|Opium Derivatives
C0002327|Alphaprodine
C0002327|4-Piperidinol, 1,3-dimethyl-4-phenyl-, propanoate (ester), cis-
C0002327|Alphaprodine [Chemical/Ingredient]
C0002327|Alphaprodine (substance)
C0006405|Buprenorphine
C0006405|6,14-Ethenomorphinan-7-methanol, 17-(cyclopropylmethyl)-alpha-(1,1-dimethylethyl)-4,5-epoxy-18,19-dihydro-3-hydroxy-6-methoxy-alpha-methyl-, (5alpha,7alpha(S))-
C0006405|Buprenorphine [Chemical/Ingredient]
C0006405|Buprenorphine product
C0006405|Buprenorphine product (product)
C0006405|Buprenorphine (product)
C0006405|Buprenorphine (substance)
C0006491|Butorphanol
C0006491|Morphinan-3,14-diol, 17-(cyclobutylmethyl)-
C0006491|17-(Cyclobutylmethyl)morphinan-3,14-diol
C0006491|Butorphanol [Chemical/Ingredient]
C0006491|Butorphanol product
C0006491|Butorphanol product (product)
C0006491|Butorphanol (product)
C0006491|Butorphanol (substance)
C0009214|Codeine
C0009214|N Methylmorphine
C0009214|Morphinan-6-ol, 7,8-didehydro-4,5-epoxy-3-methoxy-17-methyl-, (5alpha,6alpha)-
C0009214|codeine (medication)
C0009214|narcotics codeine
C0009214|Codeine [Chemical/Ingredient]
C0009214|N-Methylmorphine
C0009214|Methyl morphine
C0009214|Methylmorphine
C0009214|Codeine (product)
C0009214|Codeine (substance)
C0011817|D Moramide
C0011817|Dextromoramide
C0011817|Pyrrolidine, 1-(3-methyl-4-(4-morpholinyl)-1-oxo-2,2-diphenylbutyl)-, (S)-
C0011817|MORAMIDE D
C0011817|Pyrrolamidol
C0011817|D-Moramide
C0011817|Dextromoramide [Chemical/Ingredient]
C0011817|SKF-5137
C0011817|4-(2-Methyl-4-Oxo-3,3-Diphenyl-4-(1-Pyrrolidinyl)Butyl)Morpholine
C0011817|R-875
C0011817|(+)-4-(2-Methyl-4-Oxo-3,3-Diphenyl-4-(1-Pyrrolidinyl)Butyl)Morpholine
C0011817|D-2,2-Diphenyl-3-Methyl-4-Morpholinobutyrylpyrrolidine
C0011817|(+)-1-(3-Methyl-4-Morpholino-2,2-Diphenylbutyryl)Pyrrolidine
C0011817|1-((3S)-3-Methyl-4-(4-Morpholinyl)-1-Oxo-2,2-Diphenylbutyl)Pyrrolidine
C0011817|Dextromoramide (product)
C0011817|Dextromoramide (substance)
C0011892|Heroin
C0011892|Morphinan-3,6-diol, 7,8-didehydro-4,5-epoxy-17-methyl- (5alpha,6alpha)-, diacetate (ester)
C0011892|diacetylmorphine
C0011892|Diamorphine
C0011892|Heroin [Chemical/Ingredient]
C0011892|heroin (Schedule I substance)
C0011892|Junk
C0011892|Smack
C0011892|Skag
C0011892|H
C0011892|Acetomorphine
C0011892|Black tar
C0011892|Heroin (product)
C0011892|Heroin (substance)
C0012305|Dihydromorphine
C0012305|Morphinan-3,6-diol, 4,5-epoxy-17-methyl-, (5alpha,6alpha)-
C0012305|Dihydromorphine [Chemical/Ingredient]
C0012305|Paramorphan
C0012305|Paramorfan
C0012306|Hydromorphone
C0012306|Morphinan-6-one, 4,5-epoxy-3-hydroxy-17-methyl-, (5alpha)-
C0012306|Dihydromorphinone
C0012306|Hydromorphon
C0012306|hydromorphone (medication)
C0012306|Hydromorphone [Chemical/Ingredient]
C0012306|(-)-Hydromorphone
C0012306|Hydromorphone (substance)
C0012306|Hydromorphone (product)
C0015109|Ethylmorphine
C0015109|Morphinan-6-ol, 7,8-didehydro-4,5-epoxy-3-ethoxy-17-methyl-, (5alpha,6alpha)-
C0015109|Ethylmorphine (product)
C0015109|Codethyline
C0015109|Ethomorphine
C0015109|Ethylmorphine [Chemical/Ingredient]
C0015109|(5Alpha,6Alpha)-7,8-Didehydro-4,5-Epoxy-3-Ethoxy-17-Methylmorphinan-6-Ol
C0015109|Ethyl morphine
C0015109|Ethyl morphine (substance)
C0015134|Etorphine
C0015134|6,14-Ethenomorphinan-7-methanol, 4,5-epoxy-3-hydroxy-6-methoxy-alpha,17-dimethyl-alpha-propyl-, (5alpha,7alpha(R))-
C0015134|Ethorphine
C0015134|Etorphine [Chemical/Ingredient]
C0015134|Etorphine (substance)
C0015846|Fentanyl
C0015846|Propanamide, N-phenyl-N-(1-(2-phenylethyl)-4-piperidinyl)-
C0015846|Fentyl
C0015846|fentanyl (medication)
C0015846|Fentanyl [Chemical/Ingredient]
C0015846|Phentanyl
C0015846|N-(1-phenethylpiperidin-4-yl)-N-phenylpropionamide
C0015846|local anesthetic fentanyl (medication)
C0015846|local anesthetic fentanyl
C0015846|Fentanyl product
C0015846|Fentanyl (product)
C0015846|Fentanyl (substance)
C0020264|Hydrocodone
C0020264|Morphinan-6-one, 4,5-epoxy-3-methoxy-17-methyl-, (5alpha)-
C0020264|Hydrocodone [Chemical/Ingredient]
C0020264|Dihydrocodeinone
C0020264|Hydrocodon
C0020264|Hydrocodone (product)
C0020264|Hydrocodone (substance)
C0023586|Levorphanol
C0023586|Morphinan-3-ol, 17-methyl-
C0023586|Levorphanol [Chemical/Ingredient]
C0023586|Levodroman
C0023586|Levorphan
C0023586|Levorphanol (product)
C0023586|Levorphanol (substance)
C0025376|Meperidine
C0025376|4-Piperidinecarboxylic acid, 1-methyl-4-phenyl-, ethyl ester
C0025376|Isonipecain
C0025376|Meperidine [Chemical/Ingredient]
C0025376|Pethidine
C0025376|narcotics meperidine
C0025376|meperidine (medication)
C0025376|Meperidine (product)
C0025376|Meperidine (substance)
C0025387|Meptazinol
C0025387|Phenol, 3-(3-ethylhexahydro-1-methyl-1H-azepin-3-yl)-
C0025387|Meptazinol [Chemical/Ingredient]
C0025387|M-(3-Ethylhexahydro-1-Methyl-1H-Azepin-3-Yl)Phenol
C0025387|Meptazinol [anesthesia] (product)
C0025387|Meptazinol [analgesic] (product)
C0025387|Meptazinol [anaesthesia]
C0025387|Meptazinol [analgesic]
C0025387|Meptazinol [anesthesia]
C0025387|Meptazinol (product)
C0025387|Meptazinol (substance)
C0025387|Meptazinol [analgesic] (substance)
C0025387|Meptazinol [anesthesia] (substance)
C0025607|Methadyl Acetate
C0025607|methadylacetate
C0025607|Benzeneethanol, beta-(2-(dimethylamino)propyl)-alpha-ethyl-beta-phenyl-, acetate (ester)
C0025607|acetylmethadol
C0025607|Methadyl Acetate [Chemical/Ingredient]
C0025607|6-(Dimethylamino)-4,4-Diphenyl-3-Heptanol Acetate
C0026549|Morphine
C0026549|Morphinan-3,6-diol, 7,8-didehydro-4,5-epoxy-17-methyl- (5alpha,6alpha)-
C0026549|Morphia
C0026549|Morphine [Chemical/Ingredient]
C0026549|narcotics morphine
C0026549|morphine (medication)
C0026549|Morphine (product)
C0026549|Morphine (substance)
C0026549|MORPH
C0027348|Nalbuphine
C0027348|Morphinan-3,6,14-triol, 17-(cyclobutylmethyl)-4,5-epoxy-, (5alpha,6alpha)-
C0027348|Nalbuphine [Chemical/Ingredient]
C0027348|Nalbuphine product (product)
C0027348|Nalbuphine product
C0027348|Nalbuphine (product)
C0027348|Nalbuphine (substance)
C0029112|Opium
C0029112|opium preparations (medication)
C0029112|opium preparations
C0029112|Opium [Chemical/Ingredient]
C0029112|Opium preparation
C0029112|Opium (substance)
C0029112|Opium preparation (substance)
C0029112|Opium preparation (product)
C0030049|Oxycodone
C0030049|Morphinan-6-one, 4,5-epoxy-14-hydroxy-3-methoxy-17-methyl-, (5alpha)-
C0030049|4,5-Epoxy-14-hydroxy-3-methoxy-17-methylmorphinan-6-one
C0030049|oxycodone (medication)
C0030049|synthetic narcotics oxycodone
C0030049|Dihydrohydroxycodeinone
C0030049|Oxycodone [Chemical/Ingredient]
C0030049|Oxycodeinon
C0030049|Dinarkon
C0030049|Dihydrone
C0030049|Oxycone
C0030049|Oxycodone product (product)
C0030049|Oxycodone product
C0030049|14-Hydroxydihydrocodeinone
C0030049|Oxycodone (substance)
C0030049|Oxycodone SR
C0030049|Oxycodone (product)
C0030073|Oxymorphone
C0030073|Morphinan-6-one, 4,5-epoxy-3,14-dihydroxy-17-methyl-, (5alpha)-
C0030073|Oxymorphone [Chemical/Ingredient]
C0030073|Morphinan-6-One, 4,5-Epoxy-3,14-Dihydroxy-17-Methyl-
C0030073|4,5Alpha-Epoxy-3,14-Dihydroxy-17-Methylmorphinan-6-One
C0030073|Oxymorphone (substance)
C0030073|Oxymorphone product (product)
C0030073|Oxymorphone product
C0030873|Pentazocine
C0030873|2,6-Methano-3-benzazocin-8-ol, 1,2,3,4,5,6-hexahydro-6,11-dimethyl-3-(3-methyl-2-butenyl)-, (2alpha,6alpha,11R*)-
C0030873|pentazocine (medication)
C0030873|synthetic narcotics pentazocine
C0030873|Pentazocine [Chemical/Ingredient]
C0030873|Pentazocine (product)
C0030873|Pentazocine (substance)
C0031376|Phenazocine
C0031376|2,6-Methano-3-benzazocin-8-ol, 1,2,3,4,5,6-hexahydro-6,11-dimethyl-3-(2-phenylethyl)-
C0031376|Phenazocine [Chemical/Ingredient]
C0031376|Phenbenzorphan
C0031376|Phenethylazocine
C0031376|Phenazocine (product)
C0031376|Phenazocine (substance)
C0031432|Phenoperidine
C0031432|4-Piperidinecarboxylic acid, 1-(3-hydroxy-3-phenylpropyl)-4-phenyl-, ethyl ester
C0031432|Fenoperidine
C0031432|Phenoperidine [Chemical/Ingredient]
C0031432|Phenoperidine (product)
C0031432|Phenoperidine (substance)
C0031982|Pirinitramide
C0031982|(1,4'-Bipiperidine)-4'-carboxamide, 1'-(3-cyano-3,3-diphenylpropyl)-
C0031982|Piritramide
C0031982|Pirinitramide [Chemical/Ingredient]
C0031982|Piritramid
C0031982|Piritramide (substance)
C0031982|1'-(3-Cyano-3,3-diphenylpropyl)-(1,4'-bipiperidine)-4'-carboxamide
C0031982|(1,4'-Bipiperidine)-4'-carboxamide, 1'-(3-Cyano-3,3-diphenylpropyl)
C0031982|R 3365
C0033400|Promedol
C0033400|4-Piperidinol, 1,2,5-trimethyl-4-phenyl-, propanoate (ester)
C0033400|Dimethylmeperidine
C0033400|Promedol [Chemical/Ingredient]
C0039746|Thebaine
C0039746|Morphinan, 6,7,8,14-tetradehydro-4,5-epoxy-3,6-dimethoxy-17-methyl-, (5alpha)-
C0039746|Thebaine [Chemical/Ingredient]
C0039746|3-O-Methyl-oripavin
C0039746|4,5alpha-Epoxy-3,6-dimethoxy-17-methyl-6,8-morphinadien
C0039746|Paramorphine
C0039746|Thebaine (substance)
C0040219|Tilidine
C0040219|3-Cyclohexene-1-carboxylic acid, 2-(dimethylamino)-1-phenyl-, ethyl ester, trans-(+-)-
C0040219|Tilidate
C0040219|Tilidine [Chemical/Ingredient]
C0040219|Tilidine (product)
C0040219|Tilidine (substance)
C0040610|Tramadol
C0040610|Cyclohexanol, 2-((dimethylamino)methyl)-1-(3-methoxyphenyl)-, cis-(+-)-
C0040610|Tramadol [Chemical/Ingredient]
C0040610|Tramadol (product)
C0040610|Tramadol (substance)
C0002026|Alfentanil
C0002026|Propanamide, N-(1-(2-(4-ethyl-4,5-dihydro-5-oxo-1H-tetrazol-1-yl)ethyl)-4-(methoxymethyl)-4-piperidinyl)-N-phenyl-
C0002026|Alfentanyl
C0002026|Alfentanil [Chemical/Ingredient]
C0002026|Alfentanil - chemical
C0002026|Alfentanil - chemical (substance)
C0002026|Alfentanil (product)
C0002026|Alfentanil (substance)
C0143993|Sufentanil
C0143993|Propanamide, N-(4-(methoxymethyl)-1-(2-(2-thienyl)ethyl)-4-piperidinyl)-N-phenyl-
C0143993|Sufentanil [Chemical/Ingredient]
C0143993|Sulfentanyl
C0143993|Sulfentanil
C0143993|Sufentanil (substance)
C0143993|Sufentanil product (product)
C0143993|Sufentanil product
C0033493|Propoxyphene
C0033493|D Propoxyphene
C0033493|Benzeneethanol, alpha-(2-(dimethylamino)-1-methylethyl)-alpha-phenyl-, propanoate (ester), (S-(R*,S*))-
C0033493|PROPOXYPHENE D
C0033493|Dextropropoxyphene
C0033493|Propoxyphene (product)
C0033493|Dextropropoxyphene (product)
C0033493|synthetic narcotics propoxyphene preparations
C0033493|propoxyphene preparations (medication)
C0033493|propoxyphene preparations
C0033493|D-Propoxyphene
C0033493|Dextropropoxyphene [Chemical/Ingredient]
C0033493|4-Dimethylamino-3-methyl-1,2-diphenyl-2-propoxybutane
C0033493|Propoxyphene (substance)
C0033493|Dextropropoxyphene (substance)
C0027415|Narcotics
C0027415|narcotic
C0027415|narcotics (medication)
C2193937|sodium iodide + niacinamide hydroiodide
C2193937|narcotics sodium iodide + niacinamide hydroiodide
C2193937|sodium iodide + niacinamide hydroiodide (medication)
C0355546|dextromoramide tartrate
C0355546|dextromoramide tartrate (medication)
C0355546|narcotics dextromoramide tartrate
C0355546|Dextromoramide tartrate (substance)
C0355546|Tartrate, Dextromoramide
C0282128|diacetylmorphine hydrochloride
C0282128|diacetylmorphine hydrochloride (medication)
C0282128|Heroin Hydrochloride
C0282128|Diamorphine Hydrochloride
C0282128|Heroine Hydrochloride
C0282128|Morphinan-3,6alpha-diol, 7,8-didehydro-4,5alpha-epoxy-17-methyl-, Morphine, Diacetate (ester), Hydrochloride
C0282128|Hydrochloride, Heroin
C0282128|Diamorphine HCl [cough]
C0282128|Diamorphine HCl [cough] (product)
C0282128|Diamorphine HCl [analgesic] (product)
C0282128|Diamorphine HCl [analgesic]
C0282128|Diamorphine hydrochloride (substance)
C0282128|Diamorphine HCl [analgesic] (substance)
C0282128|Diamorphine HCl [cough] (substance)
C0282128|Hydrochloride, Diacetylmorphine
C2194296|narcotics aspirin + caffeine + opium
C2194296|aspirin + caffeine + opium (medication)
C2194296|aspirin + caffeine + opium
C2194297|aspirin + phenobarbital
C2194297|aspirin + phenobarbital (medication)
C2194297|phenobarbital + aspirin (medication)
C2194297|phenobarbital + aspirin
C2194297|narcotics aspirin + phenobarbital
C2194297|Aspirin / Phenobarbital
C2146622|acetaminophen + ibuprofen + codeine
C2146622|narcotics acetaminophen + ibuprofen + codeine
C2146622|acetaminophen + ibuprofen + codeine (medication)
C2146622|Acetaminophen / Codeine / Ibuprofen
C2117853|acetaminophen + aspirin + meprobamate + caffeine + codeine (medication)
C2117853|acetaminophen + aspirin + meprobamate + caffeine + codeine
C1873942|ACETAMINOPHEN/ASPIRIN/CAFFEINE/CODEINE/SALICYLAMIDE
C1873942|acetaminophen + aspirin + salicylamide + caffeine + codeine
C1873942|acetaminophen + aspirin + salicylamide + caffeine + codeine (medication)
C1873942|Acetaminophen / Aspirin / Caffeine / Codeine / salicylamide
C2194298|aluminum aspirin + acetaminophen + chlorphenoxamine + phenobarbital (medication)
C2194298|aluminum aspirin + acetaminophen + chlorphenoxamine + phenobarbital
C2114801|promethazine + aspirin-phenacetin-caffeine + dihydrocodeine
C2114801|promethazine + aspirin-phenacetin-caffeine + dihydrocodeine (medication)
C2114800|narcotics promethazine + APAP + caffeine + dihydrocodeine
C2114800|promethazine + APAP + caffeine + dihydrocodeine
C2114800|promethazine + APAP + caffeine + dihydrocodeine (medication)
C1874363|ASPIRIN/CAFFEINE/DIHYDROCODEINE/PROMETHAZINE
C1874363|narcotics pomethazine + aspirin + caffeine + dihydrocodeine
C1874363|promethazine + aspirin + caffeine + dihydrocodeine
C1874363|promethazine + aspirin + caffeine + dihydrocodeine (medication)
C1874363|Aspirin / Caffeine / dihydrocodeine / Promethazine
C1302959|pentazocine hydrochloride + aspirin (discontinued) (medication)
C1302959|pentazocine hydrochloride + aspirin (discontinued)
C1302959|Aspirin + pentazocine hydrochloride (product)
C1302959|Aspirin + pentazocine hydrochloride
C2052847|pentazocine + aspirin + caffeine (medication)
C2052847|pentazocine + aspirin + caffeine
C0030131|p Chloroamphetamine
C0030131|p-Chloroamphetamine
C0030131|p Chloramphetamine
C0030131|para Chloroamphetamine
C0030131|Benzeneethanamine, 4-chloro-alpha-methyl-
C0030131|CHLOROAMPHETAMINE P
C0030131|CHLORAMPHETAMINE P
C0030131|PCA
C0030131|4-Chloroamphetamine
C0030131|alpha-Methyl-p-chlorophenethylamine
C0030131|narcotics patient controlled anesthesia (PCA) (medication)
C0030131|narcotics PCA
C0030131|narcotics patient controlled anesthesia (PCA)
C0030131|Parachloroamphetamine
C0030131|p-Chloramphetamine
C0030131|para-Chloroamphetamine
C0030131|p-Chloroamphetamine [Chemical/Ingredient]
C2047970|Imed panel locked
C2047970|narcotics Imed panel locked
C2047970|Imed panel locked (medication)
C0770427|Anileridine Hydrochloride
C0770427|anileridine hydrochloride (discontinued)
C0770427|narcotics anileridine hydrochloride (discontinued)
C0770427|anileridine hydrochloride (discontinued) (medication)
C0770428|anileridine phosphate (discontinued) (medication)
C0770428|anileridine phosphate (discontinued)
C0770428|narcotics anileridine phosphate (discontinued)
C0770428|Anileridine Phosphate
C0700525|Butorphanol Tartrate
C0700525|narcotics butorphanol tartrate
C0700525|butorphanol tartrate (medication)
C0700525|Butorphanol Tartrate [Chemical/Ingredient]
C0700525|(-)-17-(Cyclobutylmethyl)morphinan-3,14-diol D-(-)-tartrate (1:1) (salt)
C0700525|Butorphanol tartrate (substance)
C0700562|Alfentanil Hydrochloride
C0700562|alfentanil hydrochloride (medication)
C0700562|Alfentanil Hydrochloride [Chemical/Ingredient]
C0700562|Alfentanil hydrochloride - chemical
C0700562|Alfentanil hydrochloride - chemical (substance)
C0700562|Alfentanil hydrochloride (substance)
C2001271|Tapentadol
C2001271|Tapentadol (product)
C2001271|Tapentadol (substance)
C2001271|3-((1R,2R)-3-(dimethylamino)-1-ethyl-2-methylpropyl)phenol
C2001271|tapentadol (medication)
C2001271|narcotics tapentadol
C0306074|Empirin with Codeine
C0306074|narcotics aspirin + codeine (empirin with codeine)
C0306074|aspirin + codeine (Empirin with codeine) (medication)
C0306074|aspirin + codeine (Empirin with codeine)
C2351132|ACETAMINOPHEN/CODEINE
C2351132|Paracetamol +codeine
C2351132|Paracetamol +codiene
C2351132|codeine phosphate + acetaminophen
C2351132|codeine phosphate + acetaminophen (medication)
C2351132|narcotics acetaminophen + codeine
C2351132|acetaminophen + codeine (medication)
C2351132|acetaminophen + codeine
C2351132|acetaminophen-codeine
C2351132|Acetaminophen-Codeine Phosphate
C2351132|co-codamol
C2351132|acetaminophen - codeine
C2351132|acetaminophen, codeine drug combination
C2351132|cocodamol
C2351132|Acetaminophen+Codeine
C2351132|Acetaminophen / Codeine
C2351132|Paracetamol + codeine
C2351132|Paracetamol + codeine phosphate
C2351132|Acetaminophen + codeine phosphate (product)
C2351132|Acetaminophen + codeine phosphate
C2351132|Co-codamol (product)
C2351132|Acetaminophen #3
C2351132|Co-codamol (substance)
C2351132|Acetaminophen + codeine (product)
C2351132|Acetaminophen with Codeine
C0724655|Laudanum
C0724655|Opium tincture
C0724655|Tincture of opium
C0724655|narcotics tincture of opium
C0724655|tincture of opium (medication)
C0724655|Laudanum (substance)
C0724655|DTO
C0724655|Deodorized Tincture of Opium
C2013185|opiate alkaloid hydrochloride (Pantopan injectable) (medication)
C2013185|opiate alkaloid hydrochloride (Pantopan injectable)
C2066455|narcotic antitussives
C2066455|narcotic antitussives (medication)
C0282275|Oxymorphone Hydrochloride
C0282275|4,5-alpha-Epoxy-3,14-dihydroxy-17-methylmorphinan-6-one Hydrochloride
C0282275|oxymorphone hydrochloride (medication)
C0282275|narcotics oxymorphone hydrochloride
C0282275|Oxymorphone Hydrochloride [Chemical/Ingredient]
C0282275|Oxymorphone HCl
C0282275|Oxymorphone hydrochloride (substance)
C0717478|BELLADONNA/OPIUM
C0717478|narcotics opium + belladonna
C0717478|opium + belladonna (medication)
C0717478|opium + belladonna
C0717478|belladonna-opium
C0717478|Opium+belladonna (product)
C0717478|Opium+belladonna
C0700533|Hydromorphone Hydrochloride
C0700533|hydromorphone hydrochloride (medication)
C0700533|Hydromorphone Hydrochloride [Chemical/Ingredient]
C0700533|Hydromorphone HCl
C0700533|narcotics hydromorphone hcl
C0700533|Hydromorphone HCl (medication)
C0700533|Hydromorphone hydrochloride (product)
C0700533|Hydromorphone hydrochloride (substance)
C0700533|Dihydromorphinone hydrochloride
C2928489|Acetaminophen / Chlorpheniramine / Codeine
C2928489|acetaminophen/chlorpheniramine/codeine
C2928489|acetaminophen + chlorpheniramine + codeine (medication)
C2928489|acetaminophen + chlorpheniramine + codeine
C2928489|narcotics acetaminophen + chlorpheniramine + codeine
C0058763|14-hydroxydihydro-6 beta-thebainol 4-methyl ether
C0058763|3,4-dimethoxy-17-methylmorphinan-6 beta,14-diol
C0058763|drotebanol
C0058763|oxymethebanol
C0002772|Analgesics, Opioid
C0002772|OPIOID ANALGESICS
C0002772|[CN101] OPIOID ANALGESICS
C0049689|6-(0-acetyl)morphine
C0049689|6-acetylmorphine
C0049689|6-monoacetylmorphine
C0049689|6-O-monoacetylmorphine
C0049689|morphine-6-acetate
C0049689|6-MAM cpd
C0049689|Monoacetylmorphine
C0049689|6-O-monoacetylmorphine (substance)
C0049689|Acetylmorphine
C1992537|Methylfentanyl &#x7C; bld-ser-plas
C1993205|Narcotics and opioids &#x7C; urine
C0066619|16,17-didehydro-9,17-dimethoxy-17,18-seco-20-alpha-yohimban-16-carboxylic acid methyl ester
C0066619|mitragynine
C0041029|Trimeperidine
C0041029|Tripethidine
C0041029|Trimeperidine (substance)
C0058056|dihydrocodeine
C0058056|Dihydrocodeine Acid
C0058056|Morphinan-6-alpha-ol, 4,5-alpha-epoxy-3-methoxy-17-methyl-
C0058056|dihydrocodeine [Chemical/Ingredient]
C0058056|Dihydrocodeine (product)
C0058056|Dihydrocodeine (substance)
C1993204|Narcotics and opioids &#x7C; gastric fluid
C0058410|4,4-diphenyl-6-piperidino-3-heptanone
C0058410|dipipanone
C0058410|Phenylpiperone
C0058410|Dipipanone (product)
C0058410|Dipipanone (substance)
C0027410|Antagonists, Narcotic
C0027410|Narcotic Antagonists
C0027410|narcotic antagonist
C0027410|Antagonists, Opioid
C0027410|OPIOID ANTAG
C0027410|NARCOTIC ANTAG
C0027410|Receptor Antagonists, Opioid
C0027410|Antagonists, Opioid Receptor
C0027410|Opioid Antagonists
C0027410|Opioid Receptor Antagonists
C0027410|Opioid antagonist
C0027410|Opiate antagonist (product)
C0027410|Opiate antagonist (substance)
C0027410|Opiate antagonist
C0027410|Opiate antagonist, NOS
C0027410|Opiate Antagonists
C0068699|bis(nicotinyl)morphine
C0068699|morphine dinicotinate
C0068699|nicomorphine
C0068699|Nicomorphine (substance)
C0051908|anileridine
C0051908|Anileridine (substance)
C1993203|Narcotics and opioids &#x7C; bld-ser-plas
C1993202|Narcotics and opioids &#124; bile fluid
C1993202|Narcotics and opioids &#x7C; bile fluid
C3870663|Mitragynine+7-Hydroxymitragynine &#x7C; Urine
C3870618|Tapentadol glucuronide &#x7C; Urine
C0027409|Narcotic Analgesics
C0027409|narcotic agonists (medication)
C0027409|narcotic agonists
C0027409|Narcotic analgesic
C0027409|Narcotic analgesic product
C0027409|Analgesics, Narcotic
C0027409|Narcotic analgesic agent
C0058916|3 beta-hydroxy-2 beta-tropanecarboxylic acid
C0058916|ecgonine
C0058916|Ecgonine (product)
C0058916|Ecgonine (substance)
C0068953|6-(methylamino)-4,4-diphenyl-3-heptanol acetate
C0068953|alpha-ethyl-beta- (2-(methylamino)propyl)-beta-phenylbenzeneethanol, acetate (ester)
C0068953|paracymethadol
C0058841|dynorphin (1-13)
C0058917|ecgonine methyl ester
C0058917|methyl ecgonine
C0242402|Opioids
C0242402|Opiate agonist agent
C0242402|Opioid
C0242402|Opiate agonist (substance)
C0242402|Opiate agonist
C0242402|Opioid product
C0242402|Opiate agonist product
C0242402|Opiate agonist (product)
C0242402|Opioid (product)
C0242402|Opiate product
C0242402|Opiate agonist, NOS
C0242402|Opiate (substance)
C0242402|Opioid (substance)
C0242402|Opioid agent
C0242402|Opiate Agonists
C0430053|Opioid screening (procedure)
C0430053|Opioid screening
C0038388|Drugs, Street
C0038388|Street Drugs
C0086190|Abuse Drugs
C0086190|Drugs, Illicit
C0086190|Illicit Drugs
C0086190|Drugs of abuse
C0086190|Illegal drug (product)
C0086190|Illegal drug
C0086190|Illegal drug, NOS
C0086190|Illegal drug (substance)
C2911101|Drug abuse counseling and surveillance of drug abuser
