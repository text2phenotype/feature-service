C0150055|Chronic pain
C0150055|Chronic pain (finding)
C0232491|Chronic abdominal pain
C0457949|Chronic low back pain
C0232493|Epigastric pain
C0235296|Epigastric pain not food-related
C0743540|EPIGASTRIC PAIN ACUTE EXACERBATION	
C0743541|Chronic epigastric pain
C1533286|pain; abdomen, epigastric
C0267515|Chronic idiopathic anal pain
C0267515|Chronic idiopathic anal pain (disorder)
C2316723|Chronic pain due to injury (finding)
C2316723|Chronic pain due to injury
C2316650|Chronic pain in face (finding)
C2316650|Chronic facial pain
C2316650|Chronic pain in face
C0150055|Chronic pain
C0150055|chronic pain (diagnosis)
C0150055|rndx chronic pain (diagnosis)
C0150055|rndx chronic pain
C0150055|Pain;chronic
C0150055|Chronic Pains
C0150055|Pains, Chronic
C0150055|Chronic Pain [Disease/Finding]
C0150055|Pain, Chronic
C0150055|Chronic pain (finding)
C0150055|chronic; pain
C0150055|pain; chronic
C1719393|Chronic pain due to trauma
C1719393|chronic pain due to trauma (diagnosis)
C1719393|Chronc pain d/t trauma
C0404484|Chronic pain in female pelvis
C0404484|Chronic pelvic pain of female (disorder)
C0404484|Chronic pain in female pelvis (finding)
C0404484|Chronic pelvic pain
C0404484|Chronic pelvic pain of female
C3178789|Pains, Widespread Chronic
C3178789|Chronic Pain, Widespread
C3178789|Widespread Chronic Pains
C3178789|Pain, Widespread Chronic
C3178789|Chronic Pains, Widespread
C3178789|Pain Amplification Syndrome
C3178789|Amplified Musculoskeletal Pain Syndrome
C3178789|Chronic Widespread Pain
C3178789|Widespread Chronic Pain
C3714625|Neuropathic Pain
C3714625|Neuropathic pain (finding)
C0478148|Other chronic pain
C0478148|Chronic pain NEC
C0478148|[X]Other chronic pain
C0478148|Other chronic pain (finding)
C0478148|[X]Other chronic pain (finding)
C0478148|[X]Other chronic pain (context-dependent category)
C1740831|Chronic chest pain
C1740831|Chronic chest pain (finding)
C3649719|chronic post-procedural pain
C3649719|chronic post-procedural pain (diagnosis)
C3649719|chronic pain post-proceduraal
C3662083|Chronic pain in male pelvis (finding)
C3662083|Chronic pain in male pelvis
C3662095|Chronic pain in coccyx for more than three months (finding)
C3662095|Chronic pain in coccyx for more than three months
C3662064|Chronic nonmalignant pain
C3662064|Chronic nonmalignant pain (finding)
C3662093|Chronic pain due to malignancy
C3662093|Chronic pain due to malignancy (finding)
C3662084|Chronic thoracic back pain (finding)
C3662084|Chronic thoracic back pain
C1282310|Intermittent pain (finding)
C1282310|Intermittent pain
C2074900|chronic postoperative pain (diagnosis)
C2074900|chronic postoperative pain
C2074900|Chronic postoperative pain (finding)
C0746815|Chronic neck pain (finding)
C0746815|Chronic neck pain
C0231385|Alteration in comfort: chronic pain
C0231385|Alteration in comfort: chronic pain (finding)
C0232491|abdominal pain chronic / constant
C0232491|chronic abdominal pain
C0232491|chronic abdominal pain (symptom)
C0232491|chronic/constant abdominal pain
C0232491|Chronic abdominal pain (finding)
C0686729|Generalized chronic body aches
C0686729|Generalized chronic body pains
C0686729|Generalised chronic body aches
C0686729|Generalised chronic body pains
C0686729|Generalized chronic body pains (finding)
C1333034|Chronic Cancer Pain
C1719710|Chronic post-thoracotomy pain
C1719710|chronic post-thoracotomy pain (diagnosis)
C1719710|Chron post-thoracot pain
C1719394|Other chronic postoperative pain
C1719394|Chronic postop pain NEC
C1960183|Chronic vaginal pain
C1960183|Chronic vaginal pain (finding)
C1960183|Chronic pain in vagina
C0476481|Chronic intractable pain
C0476481|[D]Chronic intractable pain (context-dependent category)
C0476481|[D]Chronic intractable pain (situation)
C0476481|[D]Chronic intractable pain
C0476481|Chronic intractable pain (finding)
C0476481|pain; chronic, intractable
C2919655|Acute exacerbation of chronic abdominal pain (finding)
C2919655|Acute exacerbation of chronic abdominal pain
C2074609|chronic abdominal pain for more than three months (symptom)
C2074609|chronic / constant abdominal pain for more than 3 months
C2074609|chronic abdominal pain for more than three months
C2074609|chronic/constant abdominal pain for more than three months
C0400882|Chronic nonspecific abdominal pain
C0400882|Chronic nonspecific abdominal pain (finding)
C0457949|lower back pain chronic
C0457949|chronic lower back pain (symptom)
C0457949|chronic lower back pain
C0457949|Pain;back low;chronic
C0457949|Chronic low back pain (finding)
C0457949|Chronic low back pain
C0457949|CLBP - Chronic low back pain
C0457949|Chronic low back pain (disorder)
C0233180|Chaussier sign
C0233180|Chaussier's sign
C0233180|Chaussier's sign (finding)
C0232493|[D]Epigastric pain (context-dependent category)
C0232493|Epigastric pain
C0232493|abdominal pain in the central upper belly
C0232493|abdominal pain epigastric
C0232493|abdominal pain in the central upper belly (epigastric)
C0232493|epigastric pain (symptom)
C0232493|epigastric abdominal pain
C0232493|Epigastric pain epigastralgia
C0232493|Abdmnal pain epigastric
C0232493|Epigastralgia
C0232493|Pain;epigastric
C0232493|[D]Epigastric pain
C0232493|[D]Epigastric pain (situation)
C0232493|Epigastric pain (finding)
C0232493|Epigastric ache
C0232493|Pain epigastric
C0232493|epigastric; pain
C0232493|pain; epigastric
C0232493|abdomen; pain, epigastric
C0232493|Abdominal pain, epigastric
C0555727|On examination - epigastric pain on palpation (finding)
C0555727|On examination - epigastric pain on palp. (finding)
C0555727|O/E - epigastric pain on palp.
C0555727|On examination - epigastric pain on palpation
C0555727|On examination - epigastric pain on palp.
C0555727|On examination - epigastric pain on palp. (context-dependent category)
C0232494|Burning epigastric pain
C0232494|Burning epigastric pain (finding)
C0018834|Heartburn
C0018834|Pyroses
C0018834|[D]Heartburn (context-dependent category)
C0018834|[D]Heartburn NOS (context-dependent category)
C0018834|[D]Pyrosis (context-dependent category)
C0018834|Heart burn
C0018834|heartburn (symptom)
C0018834|Heartburn [Disease/Finding]
C0018834|Pyrosis
C0018834|[D]Heartburn (situation)
C0018834|Heartburn (finding)
C0018834|[D]Heartburn NOS
C0018834|[D]Pyrosis
C0018834|[D]Pyrosis (situation)
C0018834|[D]Heartburn NOS (situation)
C0018834|[D]Heartburn
C0018834|Burning reflux
C0018834|Heartburn symptom
C1291078|Epigastric discomfort
C1291078|Discomfort epigastric
C1291078|Epigastric discomfort (finding)
C0578102|Rebound tenderness of epigastrium
C0578102|Rebound tenderness of epigastrium (finding)
C0578093|Tenderness of epigastrium (finding)
C0578093|Tenderness of epigastrium
C0235296|Epigastric pain not food-related
C0743541|Chronic epigastric pain
C1533286|pain; abdomen, epigastric
