C0036916|Hepatitis STD
C0262661|History of exposure to STD
C2169446|Sex with an HCV infected person
C2169446|Sex with an HCV partner
C2169446|Sex with an HCV person
C2169446|Received blood, fluid, or drug during transfusion or infusion contaminated or infected with hepatitis virus
C0019693|HIV infection
C0019693|HIV Infections
C0019693|HTLV III Infections
C0019693|HTLV III LAV Infections
C0019693|Infection, HIV
C0019693|Infection, HTLV-III
C0019693|Infection, HTLV-III-LAV
C0019693|Infections, HIV
C0019693|Infections, HTLV-III
C0019693|Infections, HTLV-III-LAV
C0019693|Human immunodeficiency virus [HIV] disease
C0019693|Unspecified human immunodeficiency virus [HIV] disease
C0019693|LYMPHOTROPIC VIRUS TYPE III INFECTIONS HUMAN T
C0019693|HTLV III INFECT
C0019693|HTLV WIII LAV INFECTIONS
C0019693|HTLV WIII INFECTIONS
C0019693|T LYMPHOTROPIC VIRUS TYPE III INFECT HUMAN
C0019693|HIV INFECT
C0019693|HTLV III LAV INFECT
C0019693|HTLV-III/LAV infection, NOS
C0019693|human immunodeficiency virus (HIV) infection
C0019693|human immunodeficiency virus (HIV) infection (diagnosis)
C0019693|HTLV-III/LAV infection -RETIRED-
C0019693|human T-lymphotropic virus 3 (HTLV-III) infection (diagnosis)
C0019693|lymphadenopathy-associated virus (diagnosis)
C0019693|lymphadenopathy-associated virus
C0019693|human T-lymphotropic virus 3 (HTLV-III) infection
C0019693|Human immunodeficiency virus infection, unspecified
C0019693|Human immuno virus dis
C0019693|T-Lymphotropic Virus Type III Infections, Human
C0019693|HIV Infections [Disease/Finding]
C0019693|HTLV-III-LAV Infections
C0019693|HTLV-III Infections
C0019693|Infection;HIV
C0019693|Human immunodeficiency virus [HIV] disease (B20)
C0019693|HTLV-III Infection
C0019693|HTLV-III-LAV Infection
C0019693|T Lymphotropic Virus Type III Infections, Human
C0019693|[X]Human immunodeficiency virus disease (disorder)
C0019693|HTLV-III/LAV infection
C0019693|[X]Unspecified human immunodeficiency virus [HIV] disease
C0019693|Human immunodeficiency virus infection
C0019693|[X]Unspecified human immunodeficiency virus [HIV] disease (disorder)
C0019693|[X]Human immunodeficiency virus disease
C0019693|HTLV-III/LAV infection (disorder)
C0019693|HIV
C0019693|Human immunodeficiency virus syndrome
C0019693|HIV disease
C0019693|HIV infection NOS
C0019693|HIV - Human immunodeficiency virus infection
C0019693|Human immunodeficiency virus infection (disorder)
C0019693|HIV disease; disease (i.e. caused by HIV disease)
C0019693|HIV disease; infection
C0019693|disease (or disorder); HIV disease (resulting from HIV disease)
C0019693|disease (or disorder); resulting from HIV disease
C0019693|human immunodeficiency virus; disease
C0019693|immunodeficiency virus disease; human
C0019693|infection; HIV disease as cause
C0019693|Human immunodeficiency virus infection, NOS
C0019693|Human Immunodeficiency Virus
C0019693|Human immunodeficiency virus disease
C0019693|HUMAN IMMUNODEFICIENCY VIRUS [HIV] INFECTION
C0006840|Candidiases
C0006840|Candidiasis
C0006840|Moniliases
C0006840|Candidiasis, unspecified
C0006840|moniliasis
C0006840|candidiasis (diagnosis)
C0006840|Candida infections
C0006840|Candidiasis site NOS
C0006840|candidosis
C0006840|Candidiasis [Disease/Finding]
C0006840|Candidiasis (disorder)
C0006840|Candidiasis NOS (disorder)
C0006840|[X]Candidiasis, unspecified (disorder)
C0006840|Candidiasis NOS
C0006840|[X]Candidiasis, unspecified
C0006840|Candida infection
C0006840|Monilia infection
C0006840|Moniliasis monilia
C0006840|Thrush
C0006840|Candidiasis of unspecified site
C0006840|Monilia NOS
C0006840|Moniliasis NOS
C0006840|Candida NOS
C0006840|Monilial infection
C0006840|Candidal infection NOS
C0006840|Infection by Candida species
C0006840|candida; infection
C0006840|Muguet
C0006840|infection; candidal
C0006840|infection; monilia
C0006840|monilia; infection
C0006840|Candidiasis, NOS
C0006840|Candidosis, NOS
C0006840|Moniliasis, NOS
C0009663|CONDYLOMA ACCUMINATA
C0009663|Condylomata Acuminata
C0009663|Genital Wart
C0009663|Venereal Wart
C0009663|Wart, Genital
C0009663|Wart, Venereal
C0009663|condyloma acuminatum
C0009663|Anogenital (venereal) warts
C0009663|Anogenital warts
C0009663|genital warts (diagnosis)
C0009663|condyloma acuminatum (diagnosis)
C0009663|venereal warts
C0009663|genital warts
C0009663|Condyloma acuminatum -RETIRED-
C0009663|Genital warts NOS
C0009663|Condyloma
C0009663|Condylomata Acuminata [Disease/Finding]
C0009663|Warts, Genital
C0009663|Warts, Venereal
C0009663|Condylomata acuminate
C0009663|Genital warts (disorder)
C0009663|Condyloma acuminatum (disorder)
C0009663|Condylomata acuminatum
C0009663|Verruca acuminata
C0009663|Anogenital wart
C0009663|AGW - Anogenital warts
C0009663|Anogenital warts (disorder)
C0009663|condyloma; acuminata
C0009663|acuminata; condyloma
C0009663|acuminata; verruca
C0009663|anogenital; wart
C0009663|venereal; verruca
C0009663|venereal; wart
C0009663|verruca; acuminata
C0009663|verruca; venereal
C0009663|wart; anogenital
C0009663|wart; venereal
C0009663|Condyloma acuminatum (disorder) [Ambiguous]
C0019342|HERPES GENITALIA
C0019342|Genital Herpes Simplex
C0019342|Herpes Genitalis
C0019342|genital herpes
C0019342|HERPES SIMPLEX VIRUS GENITAL INFECT
C0019342|venereal herpes
C0019342|Genital herpes NOS
C0019342|Herpes Simplex, Genital
C0019342|Herpes Genitalis [Disease/Finding]
C0019342|Herpes Simplex Virus Genital Infection
C0019342|Herpes, Genital
C0019342|Genital herpes unspecified
C0019342|Genital herpes simplex NOS
C0019342|Genital herpes (disorder)
C0019342|Genital herpes unspecified (disorder)
C0019342|Genital herpes simplex NOS (disorder)
C0019342|genital herpes simplex (diagnosis)
C0019342|herpes simplex genitalis
C0019342|Genital herpes, unspecified
C0019342|Herpes genital
C0019342|Genital herpes simplex (disorder)
C0019342|genital; herpes
C0019342|herpes; genital
C0019342|Genital herpes simplex, NOS
C0018081|Gonorrhea
C0018081|Gonorrheas
C0018081|Gonococcal infections
C0018081|Gonococcal infection
C0018081|Gonococcal infection, unspecified
C0018081|gonococcal infections (diagnosis)
C0018081|Gonorrhea [Disease/Finding]
C0018081|Infection due to Neisseria gonorrheae
C0018081|The clap
C0018081|Clap
C0018081|Gonorrhoea
C0018081|Gonococcal infections NOS (disorder)
C0018081|Gonococcal infections NOS
C0018081|Gonococcal infection (disorder)
C0018081|[X]Gonococcal infection, unspecified (disorder)
C0018081|[X]Gonococcal infection, unspecified
C0018081|Gonorrhea NOS
C0018081|Gonorrhoea NOS
C0018081|Infection due to Neisseria gonorrhoeae
C0018081|GC - Gonococcus infection
C0018081|GCI - Gonococcal infection
C0018081|Gonorrhea (disorder)
C0018081|gonococcal; infection
C0018081|gonococcal
C0018081|gonorrhea; specified site not listed
C0018081|infection; gonococcal
C0018081|Gonococcal infection, NOS
C0018081|Gonorrhea, NOS
C0019163|Hepatitis B
C0019163|serum hepatitis
C0019163|hepatitis B infection
C0019163|hepatitis B infection (diagnosis)
C0019163|viral hepatitis B infection
C0019163|hepatitis, B virus
C0019163|Hep B
C0019163|Hepatitis B [Disease/Finding]
C0019163|HBV
C0019163|Serum hepatitis (disorder)
C0019163|SH - Serum hepatitis
C0019163|Viral serum hepatitis B
C0019163|Viral serum hepatitis B (disorder)
C0019163|Viral hepatitis type B
C0019163|Type B viral hepatitis (disorder)
C0019163|Viral hepatitis type B (disorder)
C0019163|Viral hepatitis B
C0019163|Type B viral hepatitis
C0019163|hepatitis; serum
C0019163|hepatitis; virus, type, B
C0019163|serum; hepatitis
C0019163|virus; hepatitis, type, B
C0024286|Lymphogranuloma Venereum
C0024286|Chlamydial lymphogranuloma (venereum)
C0024286|LGV
C0024286|Durand-Nicolas-Favre disease
C0024286|Lymphogranuloma Venereum [Disease/Finding]
C0024286|Lymphogranuloma Inguinale
C0024286|Climatic or tropical bubo
C0024286|chlamydial lymphogranuloma venereum
C0024286|chlamydial infections lymphogranuloma venereum
C0024286|chlamydial lymphogranuloma venereum (diagnosis)
C0024286|Lymphogranuloma venereum (disorder)
C0024286|Chlamydia trachomatis lymphadenitis
C0024286|LGV - Lymphogranuloma venereum
C0024286|Nicholas Favre disease
C0024286|Favre-Nicolas
C0024286|Frei
C0024286|bubo; climactic
C0024286|bubo; tropical
C0024286|inguinal; lymphogranuloma
C0024286|lymphogranuloma; chlamydial
C0024286|lymphogranuloma; inguinale
C0024286|lymphogranuloma; venereum
C0024286|lymphopathia venereum
C0024286|nicolas(-Durand)-Favre disease
C0024286|poradenitis; nostras
C0024286|Chlamydia; lymphadenitis
C0024286|Chlamydia; lymphogranuloma
C0024286|tropical; bubo
C0024286|venereum; lymphogranuloma
C0024286|Durand-Nicolas-Favre
C0024286|Nicolas-Favre disease
C0024286|Climatic AND/OR tropical bubo
C0024286|Lymphogranuloma venereum (disorder) [Ambiguous]
C0024286|climatic; bubo
C0242172|Disease, Pelvic Inflammatory
C0242172|Diseases, Pelvic Inflammatory
C0242172|Inflammatory Diseases, Pelvic
C0242172|Pelvic Inflammatory Disease
C0242172|Pelvic Inflammatory Diseases
C0242172|Unspecified inflammatory disease of female pelvic organs and tissues
C0242172|PID
C0242172|Disease, Inflammatory Pelvic
C0242172|Diseases, Inflammatory Pelvic
C0242172|Inflammatory Pelvic Diseases
C0242172|Pelvic Diseases, Inflammatory
C0242172|Inflammatory diseases of female pelvic organs
C0242172|Female pelvic inflammatory disease, unspecified
C0242172|PELVIC INFLAMM DIS
C0242172|INFLAMM PELVIC DIS
C0242172|PELVIC DIS INFLAMM
C0242172|INFLAMM DIS PELVIC
C0242172|pelvic inflammatory disease (diagnosis)
C0242172|Pelvic Infection
C0242172|Fem pelv inflam dis NOS
C0242172|Pelvic inflammatory disease (PID)
C0242172|Pelvic Disease, Inflammatory
C0242172|Inflammatory Disease, Pelvic
C0242172|Inflammatory Pelvic Disease
C0242172|Pelvic Inflammatory Disease [Disease/Finding]
C0242172|Disease;pelvic inflammatory
C0242172|Infection;pelvic inflammatory
C0242172|Inflammatory diseases of female pelvic organs (N70-N77)
C0242172|Female pelvic inflammatory disease NOS (disorder)
C0242172|Pelvic inflam. disease NOS
C0242172|Pelvic inflammatory disease NOS
C0242172|Female pelvic inflammatory disease
C0242172|Female pelvic inflammatory diseases NOS
C0242172|[X]Inflammatory diseases of female pelvic organs (disorder)
C0242172|Female pelvic infection
C0242172|Female pelvic inflammatory disease NOS
C0242172|PID - pelvic inflammatory disease
C0242172|Female pelvic inflammatory disease (disorder)
C0242172|Inflammatory disease of female pelvic organs AND/OR tissues (disorder)
C0242172|Inflam. dis.- pelvic
C0242172|[X]Inflammatory diseases of female pelvic organs
C0242172|Female pelvic inflammatory diseases NOS (disorder)
C0242172|Inflammatory disease of female pelvic organs AND/OR tissues
C0242172|PID, Pelvic Inflammatory Disease
C0242172|Inflammatory Disease (PID), Pelvic
C0242172|Disease (PID), Pelvic Inflammatory
C0242172|Pelvic Inflammatory Disease, (PID)
C0242172|Pelvic inflammation
C0242172|Disease pelvic inflammatory
C0242172|Inflammation pelvic
C0242172|PID Pelvic inflammatory disease
C0242172|Female pelvic inflammation
C0242172|inflammation; pelvic
C0242172|pelvic inflammatory disease; female
C0242172|Inflammatory disease of female pelvic organs and tissues, NOS
C0242172|Inflammatory disease of female pelvic organs AND/OR tissues [Ambiguous]
C0242172|INFLAMMATORY DISEASE OF FEMALE PELVIC ORGANS
C0242172|pelvic inflammatory infection
C0039128|Syphilis
C0039128|Syphilis, unspecified
C0039128|syphilis (diagnosis)
C0039128|Syphilis NOS
C0039128|Syphilis [Disease/Finding]
C0039128|Great Pox
C0039128|Syphilis (disorder)
C0039128|Syphilis NOS (disorder)
C0039128|[X]Syphilis, unspecified
C0039128|[X]Syphilis, unspecified (disorder)
C0039128|Lues
C0039128|Treponema pallidum infection
C0039128|Infection by Treponema pallidum
C0039128|Luetic disease
C0039128|Treponema pallidum; infection
C0039128|Syphilis, NOS
C0039128|Syphilis, stage unspecified
C0039128|Pox, Great
C0040921|Trichomoniasis
C0040921|Trichomonas Infection
C0040921|Trichomonas Infections
C0040921|Infection, Trichomonas
C0040921|Trichomoniasis, unspecified
C0040921|INFECT TRICHOMONAS
C0040921|TRICHOMONAS INFECT
C0040921|trichomoniasis (diagnosis)
C0040921|Trichomoniasis NOS
C0040921|Infections, Trichomonas
C0040921|Trichomonas Infections [Disease/Finding]
C0040921|Trichomonas NOS
C0040921|[X]Trichomoniasis, unspecified
C0040921|Trichomonas NOS (disorder)
C0040921|[X]Trichomoniasis, unspecified (disorder)
C0040921|Trich
C0040921|Infection caused by Trichomonas (disorder)
C0040921|Disease due to Trichomonadidae (disorder)
C0040921|Disease caused by Trichomonadidae
C0040921|Disease caused by Trichomonadidae (disorder)
C0040921|Infection by Trichomonas (disorder)
C0040921|Infection caused by Trichomonas
C0040921|Trichomonosis
C0040921|Disease due to Trichomonadidae
C0040921|Infection by Trichomonas
C0040921|Trichomonas; infection
C0040921|infection; Trichomonas
C0040921|Infection by Trichomonas, NOS
C0007947|Chancroid
C0007947|Chancroids
C0007947|Ulcus molle
C0007947|Chancroid [Disease/Finding]
C0007947|sexually transmitted disease chancroid
C0007947|chancroid (diagnosis)
C0007947|Chancroidal bubo
C0007947|(Chancroid [& bubo]) or (Ducrey's chancre)
C0007947|(Chancroid [& bubo]) or (Ducrey's chancre) (disorder)
C0007947|Ducrey's chancre
C0007947|Chancroid (disorder)
C0007947|Haemophilus ducreyi chancroid
C0007947|Haemophilus ducreyi infection
C0007947|Hemophilus ducreyi infection
C0007947|Hemophilus ducreyi chancroid
C0007947|Soft chancre - chancroid
C0007947|Soft sore - chancroid
C0007947|Haemophilus ducreyi
C0007947|Hemophilus ducreyi
C0007947|bubo; Haemophilus ducreyi
C0007947|bubo; Hemophilus ducreyi
C0007947|bubo; chancroidal
C0007947|bubo; soft chancre
C0007947|bubo; virulent
C0007947|chancroid; bubo
C0007947|Bacillus; Ducrey
C0007947|molle; ulcer
C0007947|ulcer; molle
C0007947|virulent; bubo
C0007947|Soft chancre
C0007947|Ducrey's disease
C0007947|Bubo due to Haemophilus ducreyi
C0007947|Simple chancre
C0007947|Chancroid (disorder) [Ambiguous]
C0007947|chancroidal; bubo
C0007947|Bubo chancroidal
C0007947|Bubo due to Hemophilus ducreyi
C0007947|Ducrey's simple soft chancre
C0007947|Ulcus molle, cutis
C0007947|Ulcus molle, skin
C0558995|Other and unspecified syphilis
C0558995|Other syphilis (disorder)
C0558995|Other and unspecified syphilis (disorder)
C0558995|Other syphilis
C0153188|Late syphilis
C0153188|Late syphilis, unspecified
C0153188|Tertiary syphilis
C0153188|late syphilis (diagnosis)
C0153188|Late syphilis NOS
C0153188|Syphilis (late)
C0153188|Syphilis, tertiary
C0153188|Late syphilis unspecified (disorder)
C0153188|[X]Late syphilis, unspecified
C0153188|Late syphilis (disorder)
C0153188|[X]Late syphilis, unspecified (disorder)
C0153188|Late syphilis unspecified
C0153188|Tertiary Treponema pallidum infection
C0153188|Late tertiary syphilis
C0153188|late; syphilitic
C0153188|syphilis; late
C0153188|syphilis; tertiary
C0153188|tertiary; syphilitic
C0153188|Late syphilis, NOS
C0039131|Syphilis, Congenital
C0039131|Congenital syphilis
C0039131|Congenital syphilis, unspecified
C0039131|SYPHILIS CONGEN
C0039131|CONGEN SYPHILIS
C0039131|congenital syphilis (diagnosis)
C0039131|Congenital syphilis NOS
C0039131|Syphilis, Congenital [Disease/Finding]
C0039131|Syphilis;congenital
C0039131|[X]Congenital syphilis, unspecified (disorder)
C0039131|Congenital syphilis NOS (disorder)
C0039131|Congenital syphilis (disorder)
C0039131|[X]Congenital syphilis, unspecified
C0039131|Unspecified congenital syphilis
C0039131|Congenital Treponema pallidum infection
C0039131|congenital; syphilitic
C0039131|hereditary; syphilitic
C0039131|syphilis; congenital
C0039131|Congenital syphilis, NOS
C0018190|Granuloma Inguinale
C0018190|granuloma inguinale (diagnosis)
C0018190|Donovanosis
C0018190|Granuloma Venereum
C0018190|Granuloma Inguinale [Disease/Finding]
C0018190|(Granuloma inguinale) or (donovanosis) or (pudendal ulcer) (disorder)
C0018190|(Granuloma inguinale) or (donovanosis) or (pudendal ulcer)
C0018190|Pudendal ulcer
C0018190|Calymmatobacterium granulomatis infection
C0018190|Infection due to Calymmatobacterium granulomatis
C0018190|Infection due to Donovania granulomatis
C0018190|Ulcerating granuloma pudendi
C0018190|Granuloma Donovani
C0018190|GI - Granuloma inguinale
C0018190|Granuloma inguinale (disorder)
C0018190|granuloma; inguinale
C0018190|granuloma; pudendi
C0018190|granuloma; venereum
C0018190|infection; Calymmatobacterium granulomatis
C0018190|inguinal; granuloma
C0018190|Calymmatobacterium granulomatis; infection
C0018190|pudendi; granuloma
C0018190|venereum; granuloma
C0018190|Granuloma pudendi
C0018190|Donovanosis;F
C0018190|Donovanosis;M
C0036916|Disease, Sexually Transmitted
C0036916|Diseases, Sexually Transmitted
C0036916|Diseases, Venereal
C0036916|Sexually Transmitted Disease
C0036916|Sexually Transmitted Diseases
C0036916|Venereal Diseases
C0036916|Disease, Venereal
C0036916|Venereal Disease
C0036916|Infections with a predominantly sexual mode of transmission
C0036916|Unspecified sexually transmitted disease
C0036916|SEX TRANSM DIS
C0036916|VENEREAL DIS
C0036916|STD
C0036916|Sexually transmitted disease, NOS
C0036916|sexually transmitted disease (diagnosis)
C0036916|VD (venereal disease)
C0036916|Venereal disease NOS
C0036916|STDs
C0036916|Sexually Transmitted Diseases [Disease/Finding]
C0036916|Disease;sexually transmitted
C0036916|Infections with a predominantly sexual mode of transmission (A50-A64)
C0036916|Sexually Transmitted Infection
C0036916|Sexually transmitted infections
C0036916|Venereal disease NOS (disorder)
C0036916|[X]Unspecified sexually transmitted disease
C0036916|[X]Infections with a predominantly sexual mode of transmission (disorder)
C0036916|[X]Infections with a predominantly sexual mode of transmission
C0036916|[X]Unspecified sexually transmitted disease (disorder)
C0036916|Statutory venereal disease
C0036916|VD - Venereal disease
C0036916|Venereal disease (disorder)
C0036916|Disease (VD), Venereal
C0036916|Venereal Disease (VD)
C0036916|VD, Venereal Disease
C0036916|STI
C0036916|Transmitted Infections, Sexually
C0036916|Infections, Sexually Transmitted
C0036916|Transmitted Infection, Sexually
C0036916|Infection, Sexually Transmitted
C0036916|Sexually transmitted disease NOS
C0036916|VD
C0036916|Venereal disease, unspecified
C0036916|STIs
C0036916|Disease with a predominantly sexual mode of transmission
C0036916|STD - Sexually transmitted disease
C0036916|Sexually transmissible disease
C0036916|Sexually transmitted infectious disease (disorder)
C0036916|Sexually transmitted infectious disease
C0036916|disease (or disorder); infectious, sexually transmitted
C0036916|disease (or disorder); sexually transmitted
C0036916|disease (or disorder); venereal
C0036916|infectious; disease, sexually transmitted
C0036916|sexual; transmitted disease
C0036916|venereal; disease
C0036916|Venereal disease, NOS
C0036916|Sexually transmitted infectious disease, NOS
C0036916|Diseases (Venereal)
C0036916|Sexually Transmitted Disorder
C0036916|Disease;venereal
C0494060|Anogenital herpesviral [herpes simplex] infection
C0494060|Anogenital herpesviral infection, unspecified
C0494060|Anogenital herpesviral [herpes simplex] infections
C0494060|Anogenital herpes
C0494060|Anogenital herpes simplex virus infection
C0494060|Anogenital herpesviral infection
C0494060|HSV - Anogenital herpes simplex virus infection
C0494060|Anogenital herpesviral infection (disorder)
C0494060|herpes; anogenital
C0494060|infection; viral, herpesvirus, anogenital
C0494060|anogenital; herpes
C0494060|viral; infection, herpesvirus, anogenital
C0348148|Early syphilis, unspecified
C0348148|Early syphilis
C0348148|early syphilis (diagnosis)
C0348148|syphilis early
C0348148|[X]Early syphilis, unspecified
C0348148|[X]Early syphilis, unspecified (disorder)
C0348148|early; syphilitic
C0348148|syphilis; early
C0494062|Other predominantly sexually transmitted diseases, not elsewhere classified
C0494059|Other sexually transmitted chlamydial diseases
C0036918|Disease, Viral Venereal
C0036918|Diseases, Viral Venereal
C0036918|Sexually Transmitted Diseases, Viral
C0036918|Venereal Disease, Viral
C0036918|Viral Venereal Disease
C0036918|SEX TRANSM DIS VIRAL
C0036918|VENEREAL DIS VIRAL
C0036918|VIRAL VENEREAL DIS
C0036918|VIRAL SEX TRANSM DIS
C0036918|Viral Sexually Transmitted Disease
C0036918|Sexually Transmitted Disease, Viral
C0036918|Sexually Transmitted Diseases, Viral [Disease/Finding]
C0036918|Venereal Diseases, Viral
C0036918|Viral Sexually Transmitted Diseases
C0036918|Viral Venereal Diseases
C0036917|Bacterial Venereal Disease
C0036917|Disease, Bacterial Venereal
C0036917|Diseases, Bacterial Venereal
C0036917|Sexually Transmitted Diseases, Bacterial
C0036917|Venereal Disease, Bacterial
C0036917|BACT VENEREAL DIS
C0036917|SEX TRANSM DIS BACT
C0036917|BACT SEX TRANSM DIS
C0036917|VENEREAL DIS BACT
C0036917|Bacterial Sexually Transmitted Disease
C0036917|Bacterial Venereal Diseases
C0036917|Sexually Transmitted Diseases, Bacterial [Disease/Finding]
C0036917|Bacterial Sexually Transmitted Diseases
C0036917|Venereal Diseases, Bacterial
C0036917|Sexually Transmitted Disease, Bacterial
C0040843|Infection, Treponemal
C0040843|Treponemal Infection
C0040843|Treponemal Infections
C0040843|TREPONEMAL INFECT
C0040843|INFECT TREPONEMAL
C0040843|Treponema infection
C0040843|Treponema infections
C0040843|Infections, Treponemal
C0040843|Treponemal Infections [Disease/Finding]
C0040843|Treponemal disease
C3853851|sexually transmitted disease due to Chlamydia trachomatis
C3853851|venereal disease due to Chlamydia trachomatis
C3853851|sexually transmitted disease due to Chlamydia trachomatis (diagnosis)
C3853851|genitourinary venereal disease due to Chlamydia trachomatis
C3853851|sexually transmitted disease of genitourinary tract due to Chlamydia trachomatis (diagnosis)
C3853851|sexually transmitted disease of genitourinary tract due to Chlamydia trachomatis
C3853851|Venereal disease caused by Chlamydia trachomatis (disorder)
C3853851|Venereal disease due to Chlamydia trachomatis (disorder)
C3853851|Venereal disease caused by Chlamydia trachomatis
C0343727|Pathogen-negative nonspecific genital infection
C0343727|Pathogen-negative nonspecific genital infection (disorder)
C0343745|Gay bowel syndrome
C0343745|Gay bowel syndrome (disorder)
C0564699|Syphilitic/venereal/spirochaetal disease
C0564699|Syphilis/venereal/spiroch.dis.
C0564699|Syphilitic/venereal/spirochetal disease
C0564699|syphilitic/venereal/spirochetal disease (diagnosis)
C0564699|Syphilitic/venereal/spirochetal disease (disorder)
C0085166|Bacterial Vaginosis
C0085166|Nonspecific Vaginitis
C0085166|Vaginosis, Bacterial
C0085166|VAGINOSES BACT
C0085166|BACT VAGINOSES
C0085166|VAGINOSIS BACT
C0085166|VAGINITIDES BACT
C0085166|BACT VAGINITIS
C0085166|BACT VAGINOSIS
C0085166|BACT VAGINITIDES
C0085166|VAGINITIS BACT
C0085166|bacterial vaginitis (diagnosis)
C0085166|nonspecific vaginitis (diagnosis)
C0085166|vaginitis bacterial
C0085166|bacterial vaginitis
C0085166|Vaginitis, Bacterial
C0085166|Vaginitis, Nonspecific
C0085166|Bacterial Vaginoses
C0085166|Vaginoses, Bacterial
C0085166|Bacterial Vaginitides
C0085166|Vaginitides, Bacterial
C0085166|Vaginosis, Bacterial [Disease/Finding]
C0085166|Bacterial vaginosis (disorder)
C0085166|BV - Bacterial vaginosis
C0085166|NSV - Nonspecific vaginitis
C0085166|AV - Anaerobic vaginosis
C0085166|BV
C0085166|Vaginosis bacterial
C0085166|Non-specific vaginitis
C0085166|Vaginitis bacterial NOS
C0085166|Vaginosis bacterial NOS
C0558371|Venereal disease in pregnancy
C0558371|Venereal dis+ pregnancy
C0558371|Preg.+ venereal disease
C0558371|Venereal disease in pregnancy (disorder)
C0558371|pregnancy; venereal disease
C1112709|Nonspecific urethritis
C1112709|NGU (nongonococcal urethritis)
C1112709|nongonococcal urethritis
C1112709|nongonococcal urethritis (diagnosis)
C1112709|NGU
C1112709|Unspecified nongonococcal urethritis (NGU)
C1112709|Non-gonococcal urethritis
C1112709|Unspecified non-gonococcal urethritis (NGU)
C1112709|NGU - Non-gonococcal urethritis
C1112709|Nonspecific genital infection
C1112709|NSGI - Nonspecific genital infection
C1112709|Urethritis-non-specific
C1112709|NSU - Nonspecific urethritis
C1112709|Nongonococcal urethritis (disorder)
C1112709|urethritis; nongonococcal
C1112709|NGU, NOS
C1112709|Nongonococcal urethritis, NOS
C1112709|Nonspecific urethritis, NOS
C1112709|non-gonococcal urethritis (NGU)
C0029840|Other specified venereal diseases
C0029840|Venereal disease NEC
C0029840|Other specified venereal diseases (disorder)
C0343665|Syphilis or venereal disease NOS
C0343665|Syphilis or venereal disease NOS (disorder)
C0178243|Syphilis and other venereal diseases (disorder)
C0178243|Syphilis and other venereal diseases
C0343664|Other specified syphilis or other venereal diseases (disorder)
C0343664|Other specified syphilis or other venereal diseases
C0153229|Other venereal diseases
C0153229|Other venereal diseases (disorder)
C3648766|infections with predominantly sexual mode of transmission complicating pregnancy, childbirth, and puerperium
C3648766|infections with predominantly sexual mode of transmission complicating pregnancy, childbirth, and puerperium (diagnosis)
C3648766|infect w/ predominant sexual mode transmission comp preg/childbirth/puerperium
C3648768|infections with predominantly sexual mode of transmission complicating childbirth
C3648768|infections with predominantly sexual mode transmission complicating childbirth
C3648768|infections with predominantly sexual mode of transmission complicating childbirth (diagnosis)
C3648765|infections with predominantly sexual mode of transmission complicating puerperium
C3648765|infections with predominantly sexual mode transmission complicating puerperium
C3648765|infections with predominantly sexual mode of transmission complicating puerperium (diagnosis)
C3648767|infections with predominantly sexual mode of transmission complicating pregnancy
C3648767|infections with predominantly sexual mode of transmission complicating pregnancy (diagnosis)
C0275533|venereal disease in mother complicating pregnancy, childbirth, and puerperium
C0275533|infectious disease in pregnancy, childbirth, and puerperium venereal
C0275533|venereal disease in mother complicating pregnancy, childbirth, and puerperium (diagnosis)
C0275533|Venereal disease in mother complicating pregnancy, childbirth AND/OR puerperium (disorder)
C0275533|Venereal disease in mother complicating pregnancy, childbirth AND/OR puerperium
C0275533|Venereal disease in mother complicating pregnancy, childbirth or puerperium, NOS
C3839894|Sexually transmitted infectious disease in mother complicating childbirth (disorder)
C3839894|Sexually transmitted disease in childbirth
C3839894|Sexually transmitted infectious disease in mother complicating childbirth
C3839894|STD (sexually transmitted disease) in childbirth
C0343740|Donovanosis - anogenital ulcer
C0343740|Donovanosis - anogenital ulcer (disorder)
C0343742|Donovanosis - non-genital lesion
C0343742|Donovanosis - non-genital lesion (disorder)
C0030759|Infestation by Phthirus pubis
C0030759|pediculosis pubis (diagnosis)
C0030759|pediculosis pubis
C0030759|pubic lice
C0030759|pubic lice (physical finding)
C0030759|Phthirus pubis
C0030759|Infestation by crab-louse
C0030759|Infestation (by);lice;pubic
C0030759|Phthirus/pediculus pubis - pubic lice - crabs (& infestation)
C0030759|Crabs - pubic lice
C0030759|Phthiriasis pubis (organism)
C0030759|Pediculus pubis - pubic lice
C0030759|Phthirus pubis (organism)
C0030759|Phthiriasis pubis
C0030759|Phthirus pubis - pubic lice
C0030759|Phthirus/pediculus pubis - pubic lice - crabs (& infestation) (disorder)
C0030759|Pubis pediculosis
C0030759|Infestation caused by crab lice
C0030759|Infestation by Phthirus pubis (disorder)
C0030759|Infestation caused by Phthirus pubis (disorder)
C0030759|Infestation caused by Phthirus pubis
C0030759|Crabs
C0030759|Infestation by crab lice
C0030759|Crabs infestation
C0030759|Pubic louse infestation
C0030759|Phthirus pubis; pediculosis
C0030759|infestation; pubic lice
C0030759|lice; pubic lice
C0030759|pediculosis; Phthirus pubis
C0030759|pubic lice; infestation
C0030759|Phthirus pubis [pubic louse]
C0030759|Pubic louse
C0030759|Pediculus pubis
C0030759|pubic lice infestation
C0040928|Urogenital trichomoniasis
C0040928|urogenital trichomoniasis (diagnosis)
C0040928|Urogenital trichomon NOS
C0040928|Urogenital trichomoniasis, unspecified
C0040928|Urogenital trichomonas NOS (disorder)
C0040928|Unspecified urogenital trichomonas
C0040928|Urogenital trichomonas NOS
C0040928|Unspecified urogenital trichomonas (disorder)
C0040928|Urogenital infection by Trichomonas vaginalis (disorder)
C0040928|Urogenital infection caused by Trichomonas vaginalis (disorder)
C0040928|Urogenital infection caused by Trichomonas vaginalis
C0040928|Urogenital infection by Trichomonas vaginalis
C0040928|TV - Trichomonas vaginalis infection
C0040928|Trichs - Trichomonas vaginalis infection
C0040928|Urogenital trichomonas
C0348156|Other specified predominantly sexually transmitted diseases
C0348156|[X]Other specified predominantly sexually transmitted diseases (disorder)
C0348156|[X]Other specified predominantly sexually transmitted diseases
C0554632|Anogenital Human Papilloma Virus Infection
C0554632|Anogenital Human Papillomavirus Infection
C0554632|Genital wart virus infection
C0554632|HPV - Anogenital human papilloma virus infection
C0554632|WVI - Genital wart virus infection
C0554632|Anogenital human papilloma virus infection (disorder)
C0589616|Genitourinary chlamydia infection
C0589616|Genitourinary chlamydia infection (disorder)
C1304005|Sexually transmitted bacterial disease affecting skin (disorder)
C1304005|Sexually transmitted bacterial disease affecting skin
C0001175|Acquired Immuno Deficiency Syndrome
C0001175|Acquired Immuno-Deficiency Syndromes
C0001175|Acquired Immunodeficiency Syndrome
C0001175|Acquired Immunodeficiency Syndromes
C0001175|AIDS
C0001175|Immuno-Deficiency Syndrome, Acquired
C0001175|Immuno-Deficiency Syndromes, Acquired
C0001175|Immunodeficiency Syndromes, Acquired
C0001175|Syndrome, Acquired Immuno-Deficiency
C0001175|Syndrome, Acquired Immunodeficiency
C0001175|Syndromes, Acquired Immuno-Deficiency
C0001175|Syndromes, Acquired Immunodeficiency
C0001175|AIDS (disorder)
C0001175|Acquired immune deficiency syndrome (AIDS)
C0001175|IMMUNODEFIC SYNDROME ACQUIRED
C0001175|ACQUIRED IMMUNO DEFIC SYNDROME
C0001175|ACQUIRED IMMUNE DEFIC SYNDROME
C0001175|IMMUNOL DEFIC SYNDROME ACQUIRED
C0001175|ACQUIRED IMMUNODEFIC SYNDROME
C0001175|acquired immunodeficiency syndrome (HIV-1 stage 6)
C0001175|acquired immunodeficiency syndrome (AIDS) (diagnosis)
C0001175|acquired immunodeficiency syndrome (AIDS)
C0001175|Acquired immune deficiency syndr
C0001175|acquired immune deficiency syndrome [AIDS]
C0001175|Acquired Immune Deficiency Syndrome
C0001175|Acquired Immunodeficiency Syndrome [Disease/Finding]
C0001175|Immunodeficiency Syndrome, Acquired
C0001175|Acquired Immuno-Deficiency Syndrome
C0001175|Immunologic Deficiency Syndrome, Acquired
C0001175|Acquired immune deficiency syndrome (disorder)
C0001175|Acquired immune defic. synd.
C0001175|Acquired human immunodeficiency virus infection syndrome NOS
C0001175|Acquired human immunodeficiency virus infection syndrome NOS (disorder)
C0001175|Acquired immune defic. syndr.
C0001175|Acquired immune deficiency syndrome (AIDS) (disorder)
C0001175|Acquired Immunodeficiency Disease
C0001175|AIDS, Acquired Immunodeficiency Syndrome
C0001175|Acquired Immunodeficiency Syndrome, AIDS
C0001175|Acquired immunodeficiency syndrome NOS
C0001175|Acquired immunodeficiency syndrome, unspecified
C0001175|Autoimmune deficiency syndrome
C0001175|AIDS - Acquired immunodeficiency syndrome
C0001175|Immunodeficiency due to human immunodeficiency virus infection
C0001175|acquired; immunodeficiency syndrome
C0001175|AIDS, NOS
C0001175|Acquired immune deficiency syndrome, NOS
C0001175|Acquired immunodeficiency syndrome, NOS
C0001175|Acquired Immune Deficiency
C0001175|Acquired Immun-Deficiency Synd
C1389248|balanitis; venereal (etiology)
C1389248|balanitis; venereal (manifestation)
C1389248|venereal; balanitis (etiology)
C1389248|venereal; balanitis (manifestation)
C1390858|bubo; inguinal, venereal
C1390858|inguinal; bubo, venereal
C1390862|bubo; venereal
C1390862|venereal; bubo
C1408024|urethritis; venereal (etiology)
C1408024|urethritis; venereal (manifestation)
C1408024|venereal; urethritis (etiology)
C1408024|venereal; urethritis (manifestation)
C1410755|vaginitis; venereal (etiology)
C1410755|vaginitis; venereal (manifestation)
C1410755|venereal; vaginitis (etiology)
C1410755|venereal; vaginitis (manifestation)
C1410801|venereal; vulvitis (etiology)
C1410801|venereal; vulvitis (manifestation)
C1410801|vulvitis; venereal (etiology)
C1410801|vulvitis; venereal (manifestation)
C1410802|venereal; vulvovaginitis (etiology)
C1410802|venereal; vulvovaginitis (manifestation)
C1410802|vulvovaginitis; venereal (etiology)
C1410802|vulvovaginitis; venereal (manifestation)
C0221385|Syphilitic gumma
C0221385|Syphiloma
C0221385|Gumma (syphilitic)
C0221385|Syphilitic gumma (disorder)
C0221385|syphilitic gumma (diagnosis)
C0221385|syphilis gummatous
C0221385|gumma; syphilitic
C0221385|syphilis; gumma
C0221385|Syphilitic gumma, NOS
C0275865|Congenital syphilitic osteochondritis
C0275865|congenital syphilitic osteochondritis (diagnosis)
C0275865|Congenital syphilitic osteochondritis (disorder)
C0275865|Congenital syphilitic epiphysitis
C0275865|Congenital syphilitic osteochondropathy
C0275865|Wegner's disease
C0275865|Syphilitic osteochondritis
C0153149|Hepatitis in secondary syphilis
C0153149|secondary syphilis with hepatitis
C0153149|secondary syphilis with hepatitis (diagnosis)
C0153149|Syphilitic hepatitis
C0153149|Secondary syphilitic hepatitis
C0153149|Secondary syphilis of liver
C0153149|syphilis secondary of liver
C0153149|Secondary syphilis of liver (diagnosis)
C0153149|Hepatitis in secondary syphilis (disorder)
C0153149|Secondary syphilis of liver (disorder)
C0039130|Syphilis, Cardiovascular
C0039130|Cardiovascular syphilis
C0039130|CV syphilis
C0039130|cardiovascular syphilis (diagnosis)
C0039130|Cardiovascular syph NOS
C0039130|Cardiovascular syphilis, unspecified
C0039130|Syphilis, Cardiovascular [Disease/Finding]
C0039130|Cardiovascular syphilis NOS (disorder)
C0039130|Cardiovascular syphilis (disorder)
C0039130|Cardiovascular syphilis NOS
C0039130|cardiovascular; syphilitic (etiology)
C0039130|cardiovascular; syphilitic (manifestation)
C0039130|disease (or disorder); heart, syphilitic (etiology)
C0039130|disease (or disorder); heart, syphilitic (manifestation)
C0039130|syphilis; cardiovascular (etiology)
C0039130|syphilis; cardiovascular (manifestation)
C0039130|Cardiovascular syphilis, NOS
C0039223|Tabes Dorsalis
C0039223|Neurosyphilis, Tabetic
C0039223|Spinalis, Tabes
C0039223|Tabetic neurosyphilis
C0039223|Tabes Spinalis
C0039223|Tabes Dorsalis [Disease/Finding]
C0039223|Tabes dorsalis - neurosyphilis
C0039223|Tabes dorsalis (disorder)
C0039223|Syphilitic posterior spinal sclerosis
C0039223|Duchenne's disease
C0039223|Tabetic neurosyphilis (disorder)
C0039223|dorsalis; tabes
C0039223|tabes; dorsalis
C0039223|Tabes dorsalis (disorder) [Ambiguous]
C0039223|Duchennes Disease
C0039223|Posterior spinal sclerosis
C0029076|Ophthalmia Neonatorum
C0029076|Ophthalmia neonatorum -RETIRED-
C0029076|neonatal conjunctivitis (diagnosis)
C0029076|neonatal conjunctivitis
C0029076|Ophthalmia neonatorum (gonococcal)
C0029076|Ophthalmia neonatorum NOS
C0029076|Ophthalmia Neonatorum [Disease/Finding]
C0029076|Neonatal conjunctivitis (disorder)
C0029076|Ophthalmia neonatorum (disorder)
C0029076|Conjunctivitis, Infantile
C0029076|Neonatal conjunctivitis NOS
C0029076|conjunctivitis; neonatal
C0029076|neonatal; conjunctivitis
C0029076|neonatorum; ophthalmia
C0029076|ophthalmia; neonatorum
C0029076|Neonatal conjunctivitis, NOS
C0029076|Ophthalmia neonatorum, NOS
C0343714|Gonococcal synovitis and tenosynovitis
C0343714|Gonococcal synovitis or tenosynovitis
C0343714|Gonococcal synovitis
C0343714|gonococcal infections synovitis or tenosynovitis
C0343714|Gonococcal synovitis or tenosynovitis (diagnosis)
C0343714|Gonococcal synovitis or tenosynovitis (disorder)
C1260915|Late syphilis, latent
C1260915|latent late syphilis
C1260915|latent late syphilis (diagnosis)
C1260915|Late syphilis latent
C1260915|Late latent syphilis
C1260915|Late latent syphilis (disorder)
C1260915|syphilis; late, latent
C1278807|urethritis due to Chlamydia trachomatis
C1278807|urethritis due to Chlamydia trachomatis (diagnosis)
C1278807|Chlamydia trachomatis urethritis
C1278807|Venereal urethritis due to chlamydia trachomatis
C1278807|Chlamydial NSU
C1278807|Urethritis chlamydial
C1278807|Chlmyd trachomatis ureth
C1278807|Urethritis;chlamydial
C1278807|Nongonococcal urethritis [NGU] due to Chlamydia trachomatis
C1278807|Other nongonococcal urethritis, chlamydia trachomatis
C1278807|Nongonococcal urethritis due to Chlamydia trachomatis
C1278807|Nongonococcal urethritis due to Chlamydia trachomatis (disorder)
C1278807|NGU due to Chlamydia trachomatis
C1278807|Chlamydia trachomatis urethritis reaction
C1278807|Chlamydial urethritis
C1278807|Chlamydia urethritis
C1278807|Urethritis caused by Chlamydia trachomatis
C1278807|Urethritis due to Chlamydia trachomatis (disorder)
C1278807|Urethritis caused by Chlamydia trachomatis (disorder)
C1278807|Chlamydial urethritis (disorder)
C1278807|Nongonococcal urethritis due to Chlamydia trachomatis (disorder) [Ambiguous]
C0343042|Taches bleuOtres
C0343042|Maculae ceruleae
C0343042|Macula cerulea (morphologic abnormality)
C0343042|Macula cerulea
C0343042|Maculae ceruleae (disorder)
C0343042|Maculae ceruleae - disorder
C0343042|Taches bleuâtres
C0851315|Acute syphil meningitis
C0851315|syphilis secondary with meningitis acute
C0851315|acute secondary syphilis with meningitis
C0851315|acute secondary syphilis with meningitis (diagnosis)
C0851315|Acute syphilitic meningitis (secondary)
C0851315|Acute secondary syphilitic meningitis
C0851315|Acute secondary syphilitic meningitis (disorder)
C0851315|Secondary acute syphilitic meningitis
C0018074|acute gonococcal infections of lower genitourinary tract
C0018074|acute gonococcal infections of lower genitourinary tract (diagnosis)
C0018074|gonococcal infections of lower genitourinary tract (diagnosis)
C0018074|gonococcal infections of lower genitourinary tract
C0018074|Acute gc infect lower gu
C0018074|Acute gonococcal infection of lower genitourinary tract
C0018074|Gonococcal infection (acute) of lower genitourinary tract
C0018074|Gonococcal infection of lower genitourinary tract
C0275654|Gonococcal salpingitis, specified as acute
C0275654|acute gonococcal salpingitis (diagnosis)
C0275654|acute gonococcal salpingitis
C0275654|Acute gc salpingitis
C0275654|Salpingitis gonococcal acute
C0275654|Gonococcal salpingitis acute
C0275654|Acute gonococcal salpingitis (disorder)
C0153199|chronic GC infections of lower GU tract
C0153199|chronic gonococcal infection of lower genitourinary tract (diagnosis)
C0153199|chronic gonorrhea of lower GU tract
C0153199|chronic gonococcal infection of lower genitourinary tract
C0153199|Chr gc infect lower gu
C0153199|Gonococcal infection, chronic, of lower genitourinary tract
C0153215|Other gonococcal infection of eye
C0153215|Gonococcal eye NEC
C0153215|Other gonococcal eye infection
C0153220|Other gonococcal infection of joint
C0153220|Gc infect joint NEC
C0153222|Gonococcal infection of anus and rectum
C0153222|Gc infect anus & rectum
C0153166|meningeal neurosyphilis (diagnosis)
C0153166|meningeal neurosyphilis
C0153166|Syphilitic meningitis
C0153166|Syphilitic aseptic meningitis
C0153166|Meningitis, syphilitic
C0153166|Meningeal syphilis
C0153166|Syphilitic meningitis (disorder)
C0153166|Syphilitic meningitis (disorder) [Ambiguous]
C0153173|syphilitic acoustic neuritis
C0153173|syphilitic acoustic neuritis (diagnosis)
C0153173|neuritis acoustic syphilitic
C0153173|acoustic neuritis due to syphilis
C0153173|Syphil acoustic neuritis
C0153173|Syphilitic acoustic neuritis (disorder)
C0153170|Syph dissem retinitis
C0153170|Syphilitic disseminated retinochoroiditis
C0153170|Syphilitic disseminated retinochoroiditis (disorder)
C0153170|syphilitic disseminated retinochoroiditis (diagnosis)
C0153168|syphilitic encephalitis
C0153168|syphilitic encephalitis (diagnosis)
C0153168|neurosyphilitic encephalitis
C0153168|neurosyphilitic encephalitis (diagnosis)
C0153168|Encephalitis due to syphilis unspecified
C0153168|Encephalitis due to syphilis unspecified (disorder)
C0153168|Syphilis encephalitis
C0153168|Syphilitic encephalitis (disorder)
C0153171|neurosyphilitic optic atrophy
C0153171|neurosyphilitic optic atrophy (diagnosis)
C0153171|Syphilitic optic atrophy
C0153171|Syphilitic optic atrophy (disorder)
C0153169|Parkinson's disease due to syphilis
C0153169|Parkinson's disease due to syphilis (diagnosis)
C0153169|Syphilitic parkinsonism
C0153169|Syphilitic parkinsonism (disorder)
C0153172|retrobulbar neuritis due to syphilis
C0153172|retrobulbar neuritis due to syphilis (diagnosis)
C0153172|Syph retrobulb neuritis
C0153172|Syphilitic retrobulbar neuritis
C0153172|Syphilitic retrobulbar neuritis (disorder)
C0153174|ruptured cerebral aneurysm due to syphilis (diagnosis)
C0153174|ruptured cerebral aneurysm due to syphilis
C0153174|Syph rupt cereb aneurysm
C0153174|Cerebral aneurysm ruptured syphilitic
C0153174|Syphilitic ruptured cerebral aneurysm (disorder)
C0153174|Syphilitic ruptured cerebral aneurysm
C0153174|Rupture of syphilitic cerebral aneurysm
C0153174|Rupture of syphilitic cerebral aneurysm (disorder)
C0153174|cerebral; aneurysm, ruptured, syphilitic (etiology)
C0153174|cerebral; aneurysm, ruptured, syphilitic (manifestation)
C0153174|rupture; cerebral aneurysm, syphilitic (etiology)
C0153174|rupture; cerebral aneurysm, syphilitic (manifestation)
C0153167|Asymptomatic neurosyphilis
C0153167|asymptomatic neurosyphilis (diagnosis)
C0153167|Asymptomat neurosyphilis
C0153167|Neurosyphilis, Asymptomatic
C0153167|Asymptomatic neurosyphilis (disorder)
C0153167|asymptomatic; neurosyphilis
C0153167|neurosyphilis; asymptomatic
C0275859|Early congenital syphilis, unspecified
C0275859|early congenital syphilis (diagnosis)
C0275859|early congenital syphilis
C0275859|Early congen syph NOS
C0275859|Congenital syphilis NOS less than two years after birth.
C0275859|Early congenital syphilis NOS (disorder)
C0275859|[X]Early congenital syphilis, unspecified (disorder)
C0275859|Early congenital syphilis NOS
C0275859|[X]Early congenital syphilis, unspecified
C0275859|Early congenital syphilis (less than 2 years)
C0275859|Early congenital syphilis (less than 2 years) (disorder)
C0275859|Early congenital syphilis, NOS (less than 2 years)
C0275859|Congenital syphilis NOS, less than two years after birth
C0153131|Syphilitic interstitial keratitis
C0153131|Syphilitic interstitial keratitis (disorder)
C0153133|Congenital syphilitic encephalitis
C0153133|congenital syphilitic encephalitis (diagnosis)
C0153133|Congen syph encephalitis
C0153133|Encephalitis due to congenital syphilis
C0153133|Congenital syphilitic encephalitis (disorder)
C0153223|Gonococcal infection of other specified sites
C0153223|Gonococcal infection of other specified site
C0153223|Gonococcal inf site NEC
C0153223|Gonococcal infection of other specified sites (disorder)
C0153228|Other gonococcal heart disease
C0153228|Gonococcal heart dis NEC
C0153228|Other gonococcal heart disease (disorder)
C3665385|congenital syphilitic gumma (diagnosis)
C3665385|Congenital syphilitic gumma
C3665385|syphilis congenital with gumma
C3665385|Congenital syphilis with gumma (diagnosis)
C3665385|Congenital syphilis with gumma
C3665385|Congenital syphilitic gumma (disorder)
C3665385|Congenital syphilis with gumma (disorder)
C3665385|gumma; syphilitic, congenital
C3665385|syphilis; gumma, congenital
C3665385|Gumma due to congenital syphilis
C0275877|neurosyphilis late congenital juvenile taboparesis
C0275877|Juvenile taboparesis
C0275877|Juvenile taboparesis (diagnosis)
C0275877|Juvenile taboparesis (disorder)
C0275877|juvenile; taboparesis
C0275877|taboparesis; juvenile
C0029751|Other specified cardiovascular syphilis
C0029751|Other specified cardiovascular syphilis -RETIRED-
C0029751|Cardiovascular syph NEC
C0029751|Other specified cardiovascular system syphilis
C0029751|Other specified cardiovascular system syphilis NOS (disorder)
C0029751|Other specified cardiovascular system syphilis NOS
C0029751|Other specified cardiovascular syphilis (disorder)
C0029751|Other specified cardiovascular system syphilis (disorder)
C0275849|Taboparesis
C0275849|Tabo paresis
C0275849|taboparesis (diagnosis)
C0275849|Taboparesis (disorder)
C0700641|Syphilitic acoustic neuritis - quaternary stage (diagnosis)
C0700641|neuritis acoustic syphilitic - quaternary stage
C0700641|Syphilitic acoustic neuritis - quaternary stage
C0700641|Syphilitic acoustic neuritis - quaternary stage (disorder)
C0275821|Primary symptomatic early syphilis
C0275821|primary early symptomatic syphilis
C0275821|Primary symptomatic early syphilis (diagnosis)
C0275821|Primary symptomatic early syphilis (disorder)
C0275822|primary syphilis of fingers (diagnosis)
C0275822|primary syphilis of fingers
C0275822|Primary finger syphilis
C0275822|Primary syphilis of fingers (disorder)
C0275822|primary; syphilitic, fingers
C0275822|syphilis; primary, fingers
C0275823|primary syphilis of lip (diagnosis)
C0275823|primary syphilis of lip
C0275823|Primary lip syphilis
C0275823|Primary syphilis of lip (disorder)
C0275823|primary; syphilitic, lip
C0275823|syphilis; lip, primary
C0275823|syphilis; primary, lip
C0275824|primary syphilis of tonsils
C0275824|primary syphilis of tonsils (diagnosis)
C0275824|Primary tonsil syphilis
C0275824|Primary syphilis of tonsils (disorder)
C0275824|primary; syphilitic, tonsils
C0275824|syphilis; primary, tonsils
C0275825|primary syphilis of breast
C0275825|primary syphilis of breast (diagnosis)
C0275825|Primary breast syphilis
C0275825|Primary syphilis of breast (disorder)
C0275826|secondary early symptomatic syphilis
C0275826|secondary early symptomatic syphilis (diagnosis)
C0275826|Secondary symptomatic early syphilis
C0275826|Secondary symptomatic early syphilis (disorder)
C0275826|early; syphilitic, symptomatic, secondary
C0275826|syphilis; early, symptomatic, secondary
C0275827|Secondary syphilis of mucous membrane (diagnosis)
C0275827|Secondary syphilis of mucous membrane
C0275827|syphilis secondary of mucous membrane
C0275827|Secondary syphilis of mucous membrane (disorder)
C0275827|secondary; syphilitic, mucous membranes
C0275827|syphilis; secondary, mucous membranes
C0275828|Condyloma latum -RETIRED-
C0275828|Condyloma latum
C0275828|Condyloma latum (disorder)
C0275828|condyloma lata
C0275828|Condylomata lata
C0275828|Flat condyloma
C0275828|CL - Condylomata lata
C0275828|condyloma; latum
C0275828|latum; condyloma
C0275829|secondary syphilis of anus (diagnosis)
C0275829|secondary syphilis of anus
C0275829|Secondary syphilis of anus (disorder)
C0275829|secondary; syphilitic, anus
C0275829|syphilis; anus, secondary
C0275829|syphilis; secondary, anus
C0275829|anus; syphilitic, secondary
C0275830|secondary syphilis of mouth (diagnosis)
C0275830|secondary syphilis of mouth
C0275830|Secondary syphilis of mouth (disorder)
C0275830|secondary; syphilitic, mouth
C0275830|syphilis; secondary, mouth
C0275831|secondary syphilis of pharynx (diagnosis)
C0275831|secondary syphilis of pharynx
C0275831|Secondary syphilis of pharynx (disorder)
C0275831|pharynx; syphilitic, secondary
C0275831|secondary; syphilitic, pharynx
C0275831|syphilis; pharynx, secondary
C0275831|syphilis; secondary, pharynx
C0275832|secondary syphilis of tonsils (diagnosis)
C0275832|secondary syphilis of tonsils
C0275832|Secondary syphilis of tonsil
C0275832|Secondary syphilis of tonsil (disorder)
C0275832|secondary; syphilitic, tonsil
C0275832|syphilis; secondary, tonsil
C0275833|secondary syphilis of vulva (diagnosis)
C0275833|secondary syphilis of vulva
C0275833|Secondary syphilis of vulva (disorder)
C0275833|secondary; syphilitic, vulva
C0275833|syphilis; secondary, vulva
C0275833|syphilis; vulva, secondary
C0275833|vulva; syphilitic, secondary
C0275837|secondary syphilis of viscera (diagnosis)
C0275837|secondary syphilis of viscera
C0275837|Secondary syphilis of viscera (disorder)
C0275837|secondary; syphilitic, viscera
C0275837|syphilis; secondary, viscera
C0275837|syphilis; visceral, secondary
C0275837|visceral; syphilitic, secondary
C0275838|Secondary syphilis of bone (disorder)
C0275838|Secondary syphilis of bone
C0275840|relapse of secondary syphilis - treated
C0275840|relapse of secondary syphilis - treated (diagnosis)
C0275840|syphilis secondary relapse - treated
C0275840|relapse secondary syphilis - treated
C0275840|Secondary syphilis, relapse (treated)
C0275840|Secondary syphilis, relapse (treated) (disorder)
C0275840|Secondary syphilis relapse, treated
C0275841|relapse of secondary syphilis - untreated (diagnosis)
C0275841|syphilis secondary relapse - untreated
C0275841|relapse secondary syphilis - untreated
C0275841|relapse of secondary syphilis - untreated
C0275841|Secondary syphilis, relapse (untreated)
C0275841|Secondary syphilis, relapse (untreated) (disorder)
C0275841|Secondary syphilis relapse, untreated
C0340379|syphilitic aortic incompetence (diagnosis)
C0340379|Syphilitic aortic incompetence
C0340379|Late quaternary syphilitic aortic regurgitation
C0340379|Syphilitic aortic regurgitation
C0340379|Syphilitic aortic incompetence (disorder)
C0275846|aortic stenosis syphilitic
C0275846|Syphilitic aortic stenosis
C0275846|Syphilitic aortic stenosis (diagnosis)
C0275846|Syphilitic aortic stenosis (disorder)
C0275847|syphilitic ostial coronary artery disease
C0275847|syphilis cardiovascular coronary artery ostial
C0275847|syphilitic ostial coronary artery disease (diagnosis)
C0275847|Syphilitic ostial coronary disease
C0275847|Syphilitic ostial coronary disease (disorder)
C0275852|gummatous neurosyphilis of central nervous system
C0275852|syphilitic gumma of central nervous system
C0275852|syphilitic gumma of central nervous system (diagnosis)
C0275852|Syphilitic gumma of central nervous system (disorder)
C0275852|central nervous system; gumma
C0275852|gumma; central nervous system
C0275852|gumma; syphilitic, central nervous system
C0275852|syphilis; gumma, central nervous system
C0275852|Syphilitic Gumma of central nervous system NOS
C0275852|Gumma of central nervous system NOS
C0275858|Latent syphilis (+ sero.) (disorder)
C0275858|Latent syphilis (+ sero.)
C0275858|Latent syphilis with positive serology (disorder)
C0275858|Latent syphilis with positive serology
C0275858|Latent syphilis with positive serology (diagnosis)
C0275858|syphilis latent with positive serology
C0275858|latent; syphilitic, positive serology
C0275858|syphilis; latent, positive serology
C0275858|Latent syphilis, NOS (+ sero.)
C0730326|congenital syphilitic choroiditis (diagnosis)
C0730326|congenital syphilitic choroiditis
C0730326|Congenital syphilitic chorioretinitis
C0730326|Congenital syphilitic choroiditis (disorder)
C0275861|Congenital syphilitic coryza
C0275861|syphilis congenital early coryza
C0275861|Congenital syphilitic coryza (diagnosis)
C0275861|Congenital syphilitic coryza (disorder)
C0275862|Congenital syphilitic hepatomegaly
C0275862|Congenital syphilitic hepatomegaly (disorder)
C0275862|Congenital syphilitic hepatomegaly (diagnosis)
C0275862|syphilis of liver congenital hepatomegaly
C0275863|Congenital syphilitic mucous patches
C0275863|syphilis congenital early mucous patches
C0275863|Congenital syphilitic mucous patches (diagnosis)
C0275863|Congenital syphilitic mucous patches (disorder)
C0275863|syphilis; mucous patches, congenital
C0275864|congenital syphilitic periostitis
C0275864|congenital syphilitic periostitis (diagnosis)
C0275864|Congenital syphilitic periostitis (disorder)
C0275866|Congenital syphilitic splenomegaly (disorder)
C0275866|Congenital syphilitic splenomegaly
C0275866|congenital syphilitic splenomegaly (diagnosis)
C0275867|congenital syphilitic pemphigus
C0275867|congenital syphilitic pemphigus (diagnosis)
C0275867|Congenital syphilitic pemphigus (disorder)
C0275867|Pemphigus syphiliticus
C0275867|pemphigus; syphilitic
C0275867|syphilis; pemphigus
C0275867|Syphilitic pemphigus
C0275868|Early latent congenital syphilis, positive serology, negative spinal fluid (disorder)
C0275868|Early latent congenital syphilis, positive serology, negative spinal fluid
C0275868|Early congenital syphilis, latent (+ serology. - C.S.F.) (disorder)
C0275868|Early latent congenital syphilis, positive serology, negative spinal fluid (diagnosis)
C0275868|Early congenital syphilis, latent (+ sero. - C.S.F.)
C0554634|Late congenital syphilis, unspecified
C0554634|late congenital syphilis (diagnosis)
C0554634|late symptomatic congenital syphilis
C0554634|late symptomatic congenital syphilis (diagnosis)
C0554634|late congenital syphilis
C0554634|Late congen syph NOS
C0554634|Congenital syphilis NOS two years or more after birth.
C0554634|Unspecified late congenital syphilis
C0554634|[X]Late congenital syphilis, unspecified
C0554634|Unspecified late congenital syphilis (disorder)
C0554634|[X]Late congenital syphilis, unspecified (disorder)
C0554634|Late congenital neurosyphilis
C0554634|Late congenital neurosyphilis (disorder)
C0554634|Late congenital syphilis (2 years OR more) (disorder)
C0554634|Late congenital syphilis (2 years OR more)
C0554634|Late congenital syphilis, symptomatic (2 years OR more)
C0554634|Late congenital syphilis, NOS (2 years or more)
C0554634|Congenital syphilis NOS, two years or more after birth
C0275873|Syphilitic saddle nose
C0275873|Syphilitic saddle nose (disorder)
C0275873|deformity; saddle nose, syphilitic
C0275873|saddle nose; due to syphilis
C0275873|saddle nose; syphilitic
C0275873|syphilis; saddle nose
C0275875|Juvenile general paresis
C0275875|Dementia paralytica juvenilis
C0275875|Dementia paralytica juvenilis (disorder)
C0275875|dementia paralytica; syphilitic, juvenilis
C0275875|dementia; paralytica, paralytic, juvenilis
C0275875|general; paresis, juvenile
C0275875|paralytic; dementia, juvenilis
C0275875|paresis; general, juvenile
C0275875|syphilis; dementia paralytica, juvenilis
C0275876|Juvenile tabes
C0275876|neurosyphilis tabes juvenile
C0275876|Juvenile tabes (diagnosis)
C0275876|Juvenile tabes (disorder)
C0275876|juvenile; tabes
C0275876|tabes; juvenile
C0275876|tabes; neurosyphilis, juvenile
C0019682|HIV
C0019682|Lymphadenopathy Associated Virus
C0019682|Lymphadenopathy-Associated Viruses
C0019682|Virus, Lymphadenopathy-Associated
C0019682|Viruses, Lymphadenopathy-Associated
C0019682|human immunodeficiency virus
C0019682|HUMAN IMMUNODEFIC VIRUSES
C0019682|IMMUNODEFIC VIRUSES HUMAN
C0019682|VIRUS HUMAN IMMUNODEFIC
C0019682|HTLV WIII
C0019682|HUMAN LYMPHOTROPIC VIRUS TYPE III A T
C0019682|HUMAN IMMUNODEFIC VIRUS
C0019682|VIRUSES HUMAN IMMUNODEFIC
C0019682|IMMUNODEFIC VIRUS HUMAN
C0019682|HTLV III
C0019682|LAV
C0019682|Human immunodeficiency virus, NOS
C0019682|Human T Cell Leukemia Virus Type III
C0019682|Virus (HIV), Human Immunodeficiency
C0019682|Human Immunodeficiency Virus (HIV)
C0019682|HIV, Human Immunodeficiency Virus
C0019682|Immunodeficiency Viruses, Human
C0019682|Acquired Immune Deficiency Syndrome Virus
C0019682|Human T Cell Lymphotropic Virus Type III
C0019682|Human T-Cell Lymphotropic Virus Type III
C0019682|LAV-HTLV-III
C0019682|Human T-Cell Leukemia Virus Type III
C0019682|Acquired Immunodeficiency Syndrome Virus
C0019682|Human T Lymphotropic Virus Type III
C0019682|Human T-Lymphotropic Virus Type III
C0019682|Immunodeficiency Virus, Human
C0019682|AIDS Virus
C0019682|Human Immunodeficiency Viruses
C0019682|Lymphadenopathy-Associated Virus
C0019682|Virus, Human Immunodeficiency
C0019682|Viruses, Human Immunodeficiency
C0019682|HTLV-III
C0019682|HIV - Human immunodeficiency virus
C0019682|Human immunodeficiency virus (organism)
C0019682|Human T-lymphotropic virus, type III (HTLV-III)
C0019682|Lymphadenopathy-associated virus (LAV)
C0019682|Lymphadenopathy-associated virus, type I (LAV-I)
C0019682|AIDS Viruses
C0019682|Virus, AIDS
C0019682|Viruses, AIDS
C0019682|Virus-HIV
C0153151|Second syphilis relapse
C0153151|secondary syphilis relapse (diagnosis)
C0153151|secondary syphilis relapse
C0153151|relapse secondary syphilis
C0153151|Secondary syphilis, relapse (disorder)
C0153151|Secondary syphilis, relapse
C0153151|Secondary syphilis relapse (disorder)
C0153158|Endocarditis syphilitic
C0153158|Syphilitic endocarditis
C0153158|syphilitic endocarditis (diagnosis)
C0153158|Syphilitic endocarditis (disorder)
C0153227|gonococcal endocarditis (diagnosis)
C0153227|gonococcal endocarditis
C0153227|Endocarditis gonococcal
C0153227|Gonococcal endocarditis (disorder)
C0153227|Endocarditis - gonococcal
C0205858|General Paralyses
C0205858|Paralyses, General
C0205858|General Paresis
C0205858|General Pareses
C0205858|Pareses, General
C0205858|Neurosyphilis, Paretic
C0205858|Paresis, General
C0205858|paretic neurosyphilis (diagnosis)
C0205858|neurosyphilis paresis (GPI)
C0205858|paretic neurosyphilis
C0205858|Dementia paralytica
C0205858|General paralysis of insane
C0205858|General paresis - neurosyphilis
C0205858|GPI - General paresis of the insane
C0205858|GPI-general paralysis insane
C0205858|Progressive paralysis (finding)
C0205858|Progressive paralysis
C0205858|Paralysis, General
C0205858|General Paralysis
C0205858|General Paresis of the Insane
C0205858|Progressive general paresis
C0205858|General paresis - neurosyphilis (disorder)
C0205858|Paralytic dementia
C0205858|general paresis; neurosyphilis
C0205858|general; paralysis
C0205858|general; paresis
C0205858|neurosyphilis; general paresis
C0205858|paralysis; general
C0205858|paralysis; progressive, general
C0205858|paralysis; progressive
C0205858|paresis; general
C0205858|paresis; syphilitic
C0205858|progressive; paralysis, general
C0205858|progressive; paralysis
C0205858|syphilis; paresis
C0205858|General paresis (disorder)
C0205858|Paresis (General)
C0205858|General paralysis of the insane
C0205858|Progressive general paralysis
C0153132|Late congenital neurosyphilis [juvenile neurosyphilis]
C0153132|Juvenile Neurosyphilis
C0153132|Juvenile neurosyph NOS
C0153132|Juvenile neurosyphilis NOS
C0153132|Juvenile neurosyphilis (disorder)
C0153132|Juvenile neurosyphilis NOS (disorder)
C0153132|Unspecified juvenile neurosyphilis
C0153132|Unspecified juvenile neurosyphilis (disorder)
C0153132|Juvenile neurosyphilis, unspecified
C0153132|Neurosyphilis, Juvenile
C0153132|Juvenile syphilis
C0153132|juvenile; neurosyphilis
C0153132|neurosyphilis; juvenile
C0275647|Acute gonorrhea of genitourinary tract (disorder)
C0275647|Acute gonorrhea of genitourinary tract
C0275647|Acute gonorrhoea of genitourinary tract
C0275647|Acute gonorrhea of genitourinary tract, NOS
C0275647|Acute gonorrhea genitourinary NOS
C0275647|Acute gonorrhea genitourinary tract NOS
C0275648|Acute gonorrhoea of lower genitourinary tract NOS
C0275648|Acute gonorrhoea of lower genitourinary tract
C0275648|Acute gonorrhea of lower genitourinary tract NOS
C0275648|Acute gonorrhea of lower genitourinary tract NOS (disorder)
C0275648|Acute gonorrhea of lower genitourinary tract (disorder)
C0275648|Acute gonorrhea of lower genitourinary tract
C0275648|Acute gonorrhea of lower genitourinary tract, NOS
C0275648|Acute gonorrhea of lower genitourinary tract [dup] (disorder)
C0343699|Acute gonorrhea of upper genitourinary tract (disorder)
C0343699|Acute gonorrhoea upper genitourinary tract NOS
C0343699|Acute unspecified gonorrhoea of upper genitourinary tract
C0343699|Acute unspecified gonorrhea of upper genitourinary tract
C0343699|Acute gonorrhoea of upper genitourinary tract
C0343699|Acute gonorrhea of upper genitourinary tract
C0343699|Acute gonorrhea upper genitourinary tract NOS (disorder)
C0343699|Acute unspecified gonorrhea of upper genitourinary tract (disorder)
C0343699|Acute gonorrhea upper genitourinary tract NOS
C0343699|Acute gonorrhea of upper genitourinary tract, NOS
C0343699|Acute gonorrhea of upper genitourinary tract [dup] (disorder)
C0275651|Acute gonococcal bartholinitis (diagnosis)
C0275651|Acute gonococcal bartholinitis
C0275651|vulvovaginitis gonococcus bartholinitis acute
C0275651|Acute gonococcal bartholinitis (disorder)
C0275652|Acute gonococcal urethritis (diagnosis)
C0275652|urethritis gonococcus, acute
C0275652|Acute gonococcal urethritis
C0275652|Urethritis gonococcal acute
C0275652|Gonococcal urethritis acute
C0275652|Neisseria gonorrheae urethritis acute
C0275652|Neisseria gonorrhoeae urethritis acute
C0275652|Acute gonococcal urethritis (disorder)
C0275653|acute gonococcal vulvovaginitis (diagnosis)
C0275653|acute gonococcal vulvovaginitis
C0275653|acute gonococcus vulvovaginitis
C0275653|Acute gonococcal vulvovaginitis (disorder)
C0275655|Chronic gonorrhea (diagnosis)
C0275655|Chronic gonorrhea
C0275655|gonococcal infections chronic
C0275655|Chronic gonorrhea (disorder)
C0275655|Chronic gonorrhoea
C0275655|Chronic gonorrhea, NOS
C0275656|Chronic gonorrhea of genitourinary tract (diagnosis)
C0275656|Chronic gonorrhea of genitourinary tract
C0275656|gonococcal infections genitourinary tract chronic
C0275656|Chronic gonorrhea of genitourinary tract (disorder)
C0275656|Chronic gonorrhoea of genitourinary tract
C0275656|Chronic gonorrhea of genitourinary tract, NOS
C0275657|Chronic gonorrhea of lower genitourinary tract
C0275657|Chronic gonorrhoea of lower genitourinary tract
C0275657|Chronic gonorrhea of lower genitourinary tract NOS (disorder)
C0275657|Chronic gonorrhoea of lower genitourinary tract NOS
C0275657|Chronic gonorrhea of lower genitourinary tract NOS
C0275657|Chronic gonorrhea of lower genitourinary tract (disorder)
C0275657|Chronic gonorrhea lower genitourinary tract
C0275657|Chronic gonorrhoea lower genitourinary tract
C0275657|Chronic gonorrhea lower genitourinary tract (disorder)
C0275657|Chronic gonorrhea of lower genitourinary tract, NOS
C0343700|Chronic gonorrhea of upper genitourinary tract NOS (disorder)
C0343700|Chronic unspecified gonorrhea of upper genitourinary tract
C0343700|Chronic gonorrhea of upper genitourinary tract
C0343700|Chronic gonorrhea of upper genitourinary tract (disorder)
C0343700|Chronic gonorrhoea of upper genitourinary tract
C0343700|Chronic gonorrhea of upper genitourinary tract NOS
C0343700|Chronic unspecified gonorrhea of upper genitourinary tract (disorder)
C0343700|Chronic unspecified gonorrhoea of upper genitourinary tract
C0343700|Chronic gonorrhoea of upper genitourinary tract NOS
C0343700|Chronic gonorrhea of upper genitourinary tract, NOS
C0343700|Chronic gonorrhea of upper genitourinary tract [dup] (disorder)
C0275659|Chronic gonococcal bartholinitis
C0275659|vulvovaginitis gonococcus bartholinitis chronic
C0275659|chronic gonococcal bartholinitis (diagnosis)
C0275659|Chronic gonococcal bartholinitis (disorder)
C0275660|chronic gonococcal urethritis (diagnosis)
C0275660|chronic gonococcal urethritis
C0275660|Neisseria gonorrheae urethritis chronic
C0275660|Neisseria gonorrhoeae urethritis chronic
C0275660|Urethritis gonococcal chronic
C0275660|Gonococcal urethritis chronic
C0275660|Chronic gonococcal urethritis (disorder)
C0275661|chronic gonococcal vulvovaginitis
C0275661|chronic gonococcal vulvovaginitis (diagnosis)
C0275661|chronic gonococcus vulvovaginitis
C0275661|Chronic gonococcal vulvovaginitis (disorder)
C0275662|Gonococcal synovitis
C0275662|gonococcal synovitis (diagnosis)
C0275662|Gonococcal synovitis (disorder)
C0275662|Gonococcal synovitis (disorder) [Ambiguous]
C0149966|Gonococcal pharyngitis
C0149966|gonococcal pharyngitis (diagnosis)
C0149966|Gonococcal infec pharynx
C0149966|Gonococcal infection of pharynx
C0149966|Pharyngeal gonococcal infection
C0149966|Gonorrhea of pharynx
C0149966|Gonorrhea of pharynx (disorder)
C0149966|Gonorrhoea of pharynx
C0149966|gonococcal; pharyngitis
C0149966|gonococcal; pharynx
C0149966|pharyngitis; gonococcal
C0149966|pharynx; gonococcal
C0275665|gonococcal proctitis (diagnosis)
C0275665|gonococcal proctitis
C0275665|Proctitis gonococcal
C0275665|Gonococcal proctitis NOS
C0275665|Gonococcal proctitis NOS (disorder)
C0275665|Gonorrhea of rectum
C0275665|Rectal gonorrhea
C0275665|Rectal gonorrhoea
C0275665|Gonorrhea of rectum (disorder)
C0275665|Gonorrhoea of rectum
C0275665|gonococcal; proctitis
C0275665|gonococcal; rectum
C0275665|proctitis; gonococcal
C0275665|rectum; gonococcal
C0546991|gonococcal tenosynovitis
C0546991|gonococcal tenosynovitis (diagnosis)
C0546991|Gonococcal teno-synovitis
C0546991|Gonococcal tenosynovitis (disorder)
C0375028|Gonococcal infection (acute) of upper genitourinary tract, site unspecified
C0375028|acute gonococcal infections of upper genitourinary tract (diagnosis)
C0375028|acute gonococcal infections of upper genitourinary tract
C0375028|Gc (acute) upper gu NOS
C0375028|Acute gonococcal infection, of upper genitourinary tract
C0375028|Gonococcal infection (acute) of upper genitourinary tract
C0375028|Acute Gonococcal Infection of Upper Genitourinary Tract
C0375028|Acute gonococcal infection of upper genitourinary tract, site unspecified
C0375029|chronic gonococcal infections of upper genitourinary tract
C0375029|chronic gonococcal infections of upper genitourinary tract (diagnosis)
C0375029|Chr gc upper gu NOS
C0375029|Chronic gonococcal infection of upper genitourinary tract, site unspecified
C0375029|Gonococcal infection, chronic, of upper genitourinary tract
C0375029|Chronic gonococcal infection of upper genitourinary tract
C0014903|Esthiomene
C0014903|esthiomene (diagnosis)
C0014903|Esthiomene (disorder)
C0275874|Late congenital syphilis, latent
C0275874|Late congenital syphilis, latent (+ sero., - C.S.F., 2 years or more)
C0275874|late latent congenital syphilis
C0275874|late latent congenital syphilis (diagnosis)
C0275874|Late congen syph latent
C0275874|Late congenital syphilis, latent (positive serology - cerebrospinal fluid, 2 years OR more) (disorder)
C0275874|Late congenital syphilis, latent (positive serology - cerebrospinal fluid, 2 years OR more)
C0275874|Late congenital syphilis, latent (+ sero., - C.S.F., 2 years OR more) (disorder)
C0275874|Late congenital syphilis - latent
C0275842|Early syphilis, latent
C0275842|Early latent syphilis, positive serology, negative cerebrospinal fluid, less than 2 years after infection (disorder)
C0275842|Early syphilis, latent (+ serology, - C.S.F., less than 2 years after) (disorder)
C0275842|Early latent syphilis, positive serology, negative cerebrospinal fluid, less than 2 years after infection
C0275842|Early syphilis, latent (+ sero., - C.S.F., less than 2 years after)
C0275842|latent early syphilis (diagnosis)
C0275842|latent early syphilis
C0275842|Early syphil latent NOS
C0275842|Latent early syphilis NOS
C0275842|Latent early syphilis NOS (disorder)
C0275842|Early latent syphilis, positive serology, negative cerebrospinal fluid, less than 2 years after infection (diagnosis)
C0275842|early latent syphilis, pos serology neg cerebrospinal fluid less 2 yrs after infection
C0275842|early latent syphilis, pos serology neg cerebrospinal fluid less 2 yrs after inf
C0275842|Early syphilis, latent, unspecified
C0275842|Latent early syphilis (disorder)
C0275842|syphilis; early, latent
C0275842|Early syphilis, latent, NOS (+ sero., - C.S.F., less than 2 years after)
C0751543|Ataxias, Locomotor
C0751543|Locomotor Ataxias
C0751543|Ataxia, Locomotor
C0751543|Locomotor Ataxia
C0751543|Meningomyelitides, Syphilitic
C0751543|Meningomyelitis, Syphilitic
C0751543|Syphilitic Meningomyelitides
C0751543|Syphilis, Spinal Cord
C0751543|Syphilitic Meningomyelitis
C0751543|Spinal Cord Syphilis
C0751543|Myelosyphilis
C0751543|ataxia; locomotor
C0751543|locomotor ataxia; syphilitic
C0751543|locomotor; ataxia
C0751543|spinal cord; syphilitic
C0751543|syphilis; locomotor ataxia
C0751543|syphilis; spinal cord
C0035012|Reiter's syndrome
C0035012|Reiter's disease
C0035012|Reiters Disease
C0035012|REITER DIS
C0035012|Disease, Reiter's
C0035012|Syndrome, Reiter
C0035012|Disease, Reiter
C0035012|REITERS DIS
C0035012|Fiessinger Leroy Reiter syndrome
C0035012|Reiter's syndrome with arthropathy
C0035012|Reiter's syndrome with arthropathy (diagnosis)
C0035012|Reiter's syndrome (diagnosis)
C0035012|Reiter Syndrome
C0035012|Reiter disease
C0035012|Reiter's disease, unspecified site
C0035012|Reiters syndrome
C0035012|Reiter's disease (disorder)
C0035012|Fiessinger-Leroy-Reiter syndrome
C0035012|Urethrooculoarticular syndrome
C0035012|arthritis; urethritica
C0035012|Reiter; triad
C0035012|Reiter
C0035012|syndrome; urethro-oculo-articular
C0035012|triad; Reiter
C0035012|urethritica; arthritis
C0035012|urethro-oculo-articular; syndrome
C0035012|uroarthritis; infectious
C0275857|Late syphilis, latent (+ sero., - C.S.F. 2 years after) (disorder)
C0275857|Late syphilis, latent (positive serology, negative cephalospinal fluid 2 years after) (disorder)
C0275857|Late syphilis, latent (positive serology, negative cephalospinal fluid 2 years after)
C0275857|latent late syphilis, positive serology, negative spinal fluid, 2+ years after infection
C0275857|latent late syphilis, positive serology, negative spinal fluid, 2+ years after infection (diagnosis)
C0275857|Late syphilis, latent (+ sero., - C.S.F. 2 years after)
C0276500|HIV I infection
C0276500|HIV I infection (diagnosis)
C0276500|Human immunodeficiency virus I infection
C0276500|Human immunodeficiency virus I infection (disorder)
C0276501|HIV II infection
C0276501|HIV II infection (diagnosis)
C0276501|HIV 2 infection
C0276501|Human immunodeficiency virus II infection
C0276501|Human immunodeficiency virus II infection (disorder)
C0153196|Gc endometritis (acute)
C0153196|Acute gonococcal endometritis
C0153196|Uterus - acute gonorrhea
C0153196|Uterus - acute gonorrhoea
C0153196|Acute gonococcal endometritis (disorder)
C0153196|endometritis gonococcal acute
C0153196|Acute gonococcal endometritis (diagnosis)
C0153196|Gonococcal endometritis (acute)
C0153196|Acute gonorrhea of uterus
C0153191|acute gonococcal cystitis
C0153191|acute gonococcal cystitis (diagnosis)
C0153191|Gc cystitis (acute)
C0153191|Gonococcal cystitis (acute)
C0153191|Bladder gonorrhea - acute
C0153191|Bladder gonorrhoea - acute
C0153191|Acute gonococcal cystitis (disorder)
C0153191|Acute gonorrhea of bladder
C0153195|Gc cervicitis (acute)
C0153195|cervicitis gonococcus acute
C0153195|Acute gonococcal cervicitis (diagnosis)
C0153195|Acute gonococcal cervicitis
C0153195|Gonococcal cervicitis acute
C0153195|Cervicitis gonococcal acute
C0153195|Acute gonococcal cervicitis (disorder)
C0153195|Gonococcal cervicitis (acute)
C0153195|Acute gonorrhea of cervix
C0153193|acute gonococcal epididymo-orchitis
C0153193|acute gonococcal epididymo-orchitis (diagnosis)
C0153193|Gc orchitis (acute)
C0153193|Gonococcal epididymo-orchitis (acute)
C0153193|Acute gonococcal epididymo-orchitis (disorder)
C0153192|Acute gonococcal prostatitis
C0153192|acute gonococcal prostatitis (diagnosis)
C0153192|Gc prostatitis (acute)
C0153192|Gonococcal prostatitis (acute)
C0153192|Acute gonococcal prostatitis (disorder)
C0153192|Gonococcal prostatitis
C0578661|Gonococcal seminal vesiculitis
C0578661|gonococcal seminal vesiculitis (diagnosis)
C0578661|Seminal vesiculitis gonococcal
C0578661|Gonococcal seminal vesiculitis (disorder)
C0153208|Chronic gonococcal salpingitis
C0153208|chronic gonococcal salpingitis (diagnosis)
C0153208|Gc salpingitis (chronic)
C0153208|Salpingitis gonococcal chronic
C0153208|Gonococcal salpingitis chronic
C0153208|Chronic gonococcal salpingitis (disorder)
C0153208|Gonococcal salpingitis (chronic)
C0153208|Gonococcal salpingitis
C0153202|chronic gonococcal cystitis (diagnosis)
C0153202|chronic gonococcal cystitis
C0153202|Gc cystitis, chronic
C0153202|Gonococcal cystitis, chronic
C0153202|Chronic gonococcal cystitis (disorder)
C0153202|Gonorrhea of bladder, chronic
C0153206|chronic gonococcal cervicitis (diagnosis)
C0153206|chronic gonococcal cervicitis
C0153206|Gc cervicitis, chronic
C0153206|Cervicitis gonococcal chronic
C0153206|Gonococcal cervicitis chronic
C0153206|Chronic gonococcal cervicitis (disorder)
C0153206|Gonococcal cervicitis, chronic
C0153206|Gonococcal cervicitis specified as chronic
C0153206|Gonorrhea of cervix, chronic
C0153207|chronic gonococcal endometritis
C0153207|chronic gonococcal endometritis (diagnosis)
C0153207|Gc endometritis, chronic
C0153207|Chronic gonococcal endometritis (disorder)
C0153207|Uterus - chronic gonorrhoea
C0153207|Uterus - chronic gonorrhea
C0153207|Gonococcal endometritis, chronic
C0153207|Gonococcal endometritis specified as chronic
C0153203|chronic gonococcal prostatitis
C0153203|chronic gonococcal prostatitis (diagnosis)
C0153203|Gc prostatitis, chronic
C0153203|Gonococcal prostatitis, chronic
C0153203|Chronic gonococcal prostatitis (disorder)
C0153203|Gonococcal prostatitis specified as chronic
C0153204|chronic gonococcal epididymo-orchitis
C0153204|chronic gonococcal epididymo-orchitis (diagnosis)
C0153204|Gc orchitis, chronic
C0153204|Gonococcal epididymo-orchitis, chronic
C0153204|Chronic gonococcal epididymo-orchitis (disorder)
C0153204|Gonococcal epididymo-orchitis specified as chronic
C0153205|chronic gonococcal seminal vesiculitis (diagnosis)
C0153205|chronic gonococcal seminal vesiculitis
C0153205|Gc sem vesiculitis, chr
C0153205|Gonococcal seminal vesiculitis, chronic
C0153205|Chronic gonococcal seminal vesiculitis (disorder)
C0153205|Gonococcal seminal vesiculitis specified as chronic
C0153205|Gonorrhea of seminal vesicle, chronic
C0153210|Gonococcal infection of eye
C0153210|gonococcal infection of eye (diagnosis)
C0153210|Eye infection gonococcal
C0153210|Gonococcal infection of eye, unspecified
C0153210|Gonococcal eye infection NOS
C0153210|Gonococcal eye infection NOS (disorder)
C0153210|Gonococcal eye infection
C0153210|Gonococcal infection of eye (disorder)
C0153210|eye; gonococcal (etiology)
C0153210|eye; gonococcal (manifestation)
C0153210|gonococcal; eye (etiology)
C0153210|gonococcal; eye (manifestation)
C0153210|Gonococcal infection of eye, NOS
C0153212|Gonococcal iridocyclitis
C0153212|Gonococcal iridocyclitis (disorder)
C0153212|Gonococcal iridocyclitis (diagnosis)
C0153212|iridocyclitis gonococcal
C0153214|gonococcal keratitis (diagnosis)
C0153214|gonococcal keratitis
C0153214|keratitis blennorrhagica
C0153214|Gonococcal keratitis (disorder)
C0153213|gonococcal endophthalmitis (diagnosis)
C0153213|gonococcal endophthalmitis
C0153213|Gonococcal endophthalmia
C0153213|Gonococcal endophthalmia (disorder)
C0153216|gonococcal infection of a joint
C0153216|gonococcal infection of joint (diagnosis)
C0153216|gonococcal infection of joint
C0153216|Gonococcal joint infection
C0153216|Arthritis gonococcal
C0153216|Gonococcal arthritis
C0153216|Gonococcal: [joint infection NOS] or [rheumatism]
C0153216|Gonococcal joint infection NOS
C0153216|Gonococcal: [joint infection NOS] or [rheumatism] (disorder)
C0153216|Rheumatism - gonococcal
C0153216|Gonococcal joint infection NOS (disorder)
C0153216|Gonococcal arthritis (disorder)
C0153216|Gonococcal rheumatism
C0153216|Gonococcal infection of joint (disorder)
C0153216|Gonococcal infection of joint, NOS
C0153216|Gonococcal infection of joint NOS
C0153218|Gonococcal bursitis
C0153218|Gonococcal bursitis (diagnosis)
C0153218|bursitis gonococcal
C0153218|Gonococcal bursitis (disorder)
C0153219|gonococcal spondylitis (diagnosis)
C0153219|gonococcal spondylitis
C0153219|Gonococcal spondylitis (disorder)
C0153225|gonococcal meningitis
C0153225|gonococcal meningitis (diagnosis)
C0153225|Meningitis gonococcal
C0153225|Gonococcal meningitis (disorder)
C0153225|Meningitis due to gonococcus
C0018077|Gonococcal peritonitis
C0018077|Peritonitis gonococcal
C0018077|Gonococcal peritonitis (disorder)
C0018077|gonococcal; peritonitis (etiology)
C0018077|gonococcal; peritonitis (manifestation)
C0018077|peritonitis; gonococcal (etiology)
C0018077|peritonitis; gonococcal (manifestation)
C0018077|Gonococcal peritonitis (disorder) [Ambiguous]
C0018075|Gonococcal keratosis
C0018075|gonococcal keratosis (diagnosis)
C0018075|Keratosis gonococcal
C0018075|Gonococcal keratosis (blennorrhagica)
C0018075|Gonococcal keratosis (disorder)
C0018075|Gonococcal blennorrhagica
C0153226|gonococcal pericarditis
C0153226|gonococcal pericarditis (diagnosis)
C0153226|Pericarditis gonococcal
C0153226|Gonococcal pericarditis (disorder)
C0153180|Renal syphilis
C0153180|Syphilis of kidney
C0153180|syphilis of kidney (diagnosis)
C0153180|Syphilis of kidney (disorder)
C0153179|Syphilis of liver
C0153179|syphilis of liver (diagnosis)
C0153179|Syphilis of liver (disorder)
C0153182|Syphilis of muscle
C0153182|syphilis of muscle (diagnosis)
C0153182|Syphilis of muscle (disorder)
C0153139|Symptomatic early syphilis (disorder)
C0153139|Symptomatic early syphilis
C0153139|early symptomatic syphilis (diagnosis)
C0153139|syphilis early symptomatic
C0153139|early symptomatic syphilis
C0153139|Early syphilis, symptomatic
C0153139|Early symptomatic syphilis (disorder)
C0153139|early; syphilitic, symptomatic
C0153139|syphilis; early, symptomatic
C0153139|Symptomatic early syphilis, NOS
C0017418|Primary genital syphilis
C0017418|Syphilis genital
C0017418|syphilis primary genital
C0017418|primary genital syphilis (diagnosis)
C0017418|Primary genital syphilis (disorder)
C0017418|Genital syphilis (primary)
C0017418|Genital chancre
C0017418|genital; syphilitic
C0017418|primary; syphilitic, genital
C0017418|syphilis; genital
C0017418|syphilis; primary, genital
C0017418|Primary genital syphilis (disorder) [Ambiguous]
C0017418|Genital syphilis
C0153140|Primary anal syphilis
C0153140|primary syphilis of anus
C0153140|primary syphilis of anus (diagnosis)
C0153140|Primary anal syphilis (disorder)
C0153140|syphilis; anus, primary
C0153140|syphilis; primary, anal
C0275834|Secondary syphilitic adenopathy
C0275834|secondary syphilis with adenopathy (diagnosis)
C0275834|secondary syphilis with adenopathy
C0275834|Syphilitic adenopathy
C0275834|Secondary syphilitic lymphadenopathy
C0275834|Adenopathy due to secondary syphilis
C0275834|Secondary syphilitic lymphadenitis
C0275834|Secondary syphilitic adenopathy (disorder)
C0275834|secondary; syphilitic, adenopathy
C0275834|secondary; syphilitic, lymphadenitis
C0275834|syphilis; secondary, adenopathy
C0275834|syphilis; secondary, lymphadenitis
C0153150|Secondary syphilis of other viscera
C0153150|Secondary syphilis of other viscera -RETIRED-
C0153150|Second syph viscera NEC
C0153150|Secondary syphilis of other viscera (disorder)
C0153177|pulmonary syphilis (diagnosis)
C0153177|pulmonary syphilis
C0153177|Syphilis of lung
C0153177|Lung disease with syphilis (disorder)
C0153177|Lung disease with syphilis
C0153177|Syphilis of lung (disorder)
C0153177|disease (or disorder); lung, in syphilis (etiology)
C0153177|disease (or disorder); lung, in syphilis (manifestation)
C0153177|lung; disease, in syphilis (etiology)
C0153177|lung; disease, in syphilis (manifestation)
C0153177|lung; syphilitic (etiology)
C0153177|lung; syphilitic (manifestation)
C0153177|pulmonary; syphilitic (etiology)
C0153177|pulmonary; syphilitic (manifestation)
C0153177|syphilis; lung (etiology)
C0153177|syphilis; lung (manifestation)
C0153177|syphilis; pulmonary (etiology)
C0153177|syphilis; pulmonary (manifestation)
C0275844|syphilis CV of an aortic artery aneurysm
C0275844|syphilis of aortic artery aneurysm
C0275844|syphilis of an aortic artery aneurysm
C0275844|syphilis of aortic artery aneurysm (diagnosis)
C0275844|Aortic aneurysm syphilitic
C0275844|Aortic aneurysm, syphil
C0275844|Syphilitic aneurysm of aorta
C0275844|Syphilitic aortic aneurysm
C0275844|Syphilitic aortic aneurysm (disorder)
C0275844|Aneurysm of aorta, specified as syphilitic
C0275844|Syphilitic dilatation of aorta
C0275844|Late quaternary syphilitic aortic aneurysm
C0275844|Syphilitic aneurysm of aorta (disorder)
C0275844|Dilatation of aorta, specified as syphilitic
C0153165|syphilitic myocarditis (diagnosis)
C0153165|syphilitic myocarditis
C0153165|syphilis CV myocarditis
C0153165|Myocarditis syphilitic
C0153165|Syphilitic myocarditis (disorder)
C0003511|Aortitides, Syphilitic
C0003511|Syphilitic Aortitides
C0003511|syphilitic aortitis (diagnosis)
C0003511|CV syphilis of aortic artery
C0003511|syphilitic aortitis
C0003511|Aortitis syphilitic
C0003511|Syphilitic aortitis (disorder)
C0003511|Late quaternary syphilitic aortitis
C0003511|aortitis; Doehle-Heller (etiology)
C0003511|aortitis; Doehle-Heller (manifestation)
C0003511|Doehle-Heller (etiology)
C0003511|Doehle-Heller (manifestation)
C0003511|Doehle-Heller; aortitis (etiology)
C0003511|Doehle-Heller; aortitis (manifestation)
C0003511|Aortitis, Syphilitic
C0153164|syphilis CV pericarditis
C0153164|syphilitic pericarditis (diagnosis)
C0153164|syphilitic pericarditis
C0153164|Pericarditis syphilitic
C0153164|Syphilitic pericarditis (disorder)
C0275854|syphilis of mitral valve
C0275854|syphilis of mitral valve (diagnosis)
C0275854|Syphilis of mitral valve (disorder)
C0275855|syphilis of tricuspid valve (diagnosis)
C0275855|syphilis of tricuspid valve
C0275855|Syphilis of tricuspid valve (disorder)
C0275856|syphilis of pulmonary valve (diagnosis)
C0275856|syphilis of pulmonary valve
C0275856|Syphilis of pulmonary valve (disorder)
C0275856|pulmonary; syphilitic, valve (etiology)
C0275856|pulmonary; syphilitic, valve (manifestation)
C0275856|syphilis; pulmonary, valve (etiology)
C0275856|syphilis; pulmonary, valve (manifestation)
C0275843|Early latent syphilis, positive serology, negative cerebrospinal fluid, with relapse after treatment (disorder)
C0275843|Early syphilis, latent (+ sero., - C.S.F., relapse after treatment)
C0275843|Early latent syphilis, positive serology, negative cerebrospinal fluid, with relapse after treatment
C0275843|Early syphilis, latent (+ serology, - C.S.F., relapse after treatment) (disorder)
C0275843|syphilis latent w/positive serology, neg cerebrospinal fluid, w/relapse after tx
C0275843|early latent syphilis with positive serology, negative cerebrospinal fluid with relapse after treatment (diagnosis)
C0275843|early latent syphilis with positive serology, negative cerebrospinal fluid with relapse after treatment
C0153146|Secondary syphilitic iridocyclitis
C0153146|secondary syphilis with iridocyclitis
C0153146|secondary syphilis with iridocyclitis (diagnosis)
C0153146|Syphilitic iridocyclitis
C0153146|Secondary syphilitic iridocyclitis (disorder)
C0153146|Syphilitic iridocyclitis (secondary)
C0002181|secondary syphilis with alopecia
C0002181|secondary syphilis with alopecia (diagnosis)
C0002181|Alopecia syphilitic
C0002181|Syphilitic alopecia
C0002181|Syphilitic alopecia (disorder)
C0275836|secondary syphilis with uveitis (diagnosis)
C0275836|secondary syphilis with uveitis
C0275836|Syphilitic uveitis NOS
C0275836|Secondary syphilitic uveitis
C0275836|Syphilitic uveitis unspecified
C0275836|Secondary syphilitic uveitis NOS
C0275836|Syphilitic uveitis unspecified (disorder)
C0275836|Secondary syphilitic uveitis NOS (disorder)
C0275836|uveitis due to secondary syphilis (diagnosis)
C0275836|Uveitis due to secondary syphilis
C0275836|Syphilitic uveitis, unspecified
C0275836|Secondary syphilitic uveitis (disorder)
C0275836|Uveitis due to secondary syphilis (disorder)
C0275836|uveitis; syphilitic (etiology)
C0275836|uveitis; syphilitic (manifestation)
C0153145|secondary syphilis with chorioretinitis (diagnosis)
C0153145|secondary syphilis with chorioretinitis
C0153145|Syphilit chorioretinitis
C0153145|Secondary syphilitic chorioretinitis
C0153145|Syphilitic chorioretinitis (secondary)
C0153145|Secondary syphilitic chorioretinitis (disorder)
C0153148|secondary syphilis with periostitis (diagnosis)
C0153148|secondary syphilis with periostitis
C0153148|Syphilitic periostitis
C0153148|Secondary syphilitic periostitis
C0153148|Secondary syphilitic periostitis (disorder)
C0275817|late syphilis involving synovium (diagnosis)
C0275817|late syphilis involving synovium
C0275817|Syphilis of synovium
C0275817|Syphilis of synovium (disorder)
C0153176|late syphilis with episcleritis
C0153176|late syphilis with episcleritis (diagnosis)
C0153176|Syphilitic episcleritis
C0153176|Syphilitic episcleritis (disorder)
C0275819|late syphilis involving bursa
C0275819|late syphilis involving bursa (diagnosis)
C0275819|Syphilis of bursa
C0275819|Syphilis of bursa (disorder)
C0153181|late syphilis involving bone (diagnosis)
C0153181|late syphilis involving bone
C0153181|Syphilis of bone
C0153181|Syphilis of bone (disorder)
C0275818|late syphilis involving tendon (diagnosis)
C0275818|late syphilis involving tendon
C0275818|Syphilis of tendon
C0275818|Syphilis of tendon (disorder)
C0275818|syphilis; tendon (etiology)
C0275818|syphilis; tendon (manifestation)
C0275818|tendon; syphilitic (etiology)
C0275818|tendon; syphilitic (manifestation)
C0153178|Syphilitic peritonitis
C0153178|late syphilis with peritonitis
C0153178|late syphilis with peritonitis (diagnosis)
C0153178|Peritonitis syphilitic
C0153178|Syphilitic peritonitis (disorder)
C0153178|Peritonitis - syphilitic
C0153134|Congenital syphilitic meningitis
C0153134|congenital syphilitic meningitis (diagnosis)
C0153134|Congen syph meningitis
C0153134|Congenital syphilitic meningitis (disorder)
C0153134|Meningitis due to congenital syphilis
C0411274|gonococcal infection of anus
C0411274|gonococcal infection of anus (diagnosis)
C0411274|Gonorrhoea of anus
C0411274|Gonorrhea of anus (disorder)
C0411274|Gonorrhea of anus
C0411274|Gonococcal anal infection
C0411274|Gonococcal anal infection (disorder)
C0411274|gonococcal; anus
C0411274|anus; gonococcal
C0275666|gonococcal infection of heart (diagnosis)
C0275666|gonococcal infection of heart
C0275666|Gonococcal heart infection
C0275666|Heart disease gonococcal NOS
C0275666|Gonococcal heart disease (disorder)
C0275666|Gonococcal heart disease
C0275666|Gonococcal heart disease, NOS
C0276055|urethritis due to ureaplasma urealyticum (diagnosis)
C0276055|urethritis due to ureaplasma urealyticum
C0276055|ureaplasma urealyticum ('T mycoplasma') urethritis
C0276055|Nongonococcal urethritis caused by Ureaplasma urealyticum
C0276055|Nongonococcal urethritis caused by Ureaplasma urealyticum (disorder)
C0276055|NGU caused by ureaplasma urealyticum
C0276055|Nongonococcal urethritis due to Ureaplasma urealyticum (disorder)
C0276055|NGU due to ureaplasma urealyticum
C0276055|Nongonococcal urethritis due to Ureaplasma urealyticum
C2732455|Exposure to sexually transmissible disorder
C2732455|Exposure to sexually transmissible disorder (event)
C0749210|exposure to syphilis
C0749210|exposure to syphilis (history)
C0749210|exposure; syphilis
C0749210|syphilis; exposure
C0744453|History of exposure to gonorrhea
C0744453|exposure to gonorrhea (history)
C0744453|exposure to gonorrhea
C0744453|exposure; gonorrhea
C0744453|gonorrhea; exposure
