C3494624|Current Heavy tobacco smoker (SNOMED:428071000124103) 
C3494624|Current Light tobacco smoker (SNOMED:428061000124105) 
C1880200|Current some day smoker	 (SNOMED:428041000124106) 
C0337671|Ex-smoker (finding)	Former smoker(SNOMED:8517006) 
C0425293|Never smoked tobacco (finding)	Never smoker (SNOMED:266919005) 
C0337664|Smoker (finding)	Smoker, current status unknown (SNOMED:77176002) 
C3266136|Smokes tobacco daily (finding)	Current every day smoker (SNOMED:449868002) 
C0425306|Tobacco smoking consumption unknown (finding)	Unknown if ever smoked (SNOMED:266927001) 
C3494624|Light tobacco smoker (finding)
C3494624|Light tobacco smoker
C3494624|Current light tobacco smoker
C3494624|current light tobacco smoker (history)
C1880200|Some Day Smoker
C1880200|Non-Daily Smoker
C1880200|Occasional Smoker
C1880200|Current Some Day Smoker
C1880200|current some day smoker (history)
C1880200|Chipper
C1880200|Occasional tobacco smoker
C1880200|Occasional tobacco smoker (finding)
C1880200|Some-day smoker
C3649460|current occasional tobacco smoker
C3649460|current occasional tobacco smoker (history)
C2114448|previous history of smoking
C2114448|previous history of smoking (history)
C3468596|former cigarette chain smoker
C3468596|former cigarette chain smoker (history)
C0337671|Former smoker
C0337671|Prior Smoker
C0337671|Past tobacco smoker
C0337671|Ex-smoker
C0337671|Ex-smoker (finding)
C0337671|Previous Tobacco Use
C0337671|Recovered smoker
C0337671|Cessation of smoking
C0337671|Ex-smoker (life style)
C3494626|Former heavy tobacco smoker (finding)
C3494626|Ex-heavy tobacco smoker
C3494626|Former heavy tobacco smoker
C3494626|former heavy tobacco smoker (history)
C3494627|Ex-light tobacco smoker
C3494627|Former light tobacco smoker
C3494627|Former light tobacco smoker (finding)
C3494627|former light tobacco smoker (history)
C3693442|stopped smoking ___ years ago
C3693442|stopped smoking ___ years ago (history)
C4041321|Ex-smoker for more than 1 year (finding)
C4041321|Ex-smoker for more than 1 year
C0521323|Aggressive ex-smoker (life style)
C0521323|Aggressive ex-smoker
C0521323|Aggressive ex-smoker (finding)
C0521323|Aggressive ex-smoker (life style) [Ambiguous]
C0425314|Ex-cigar smoker
C0425314|Ex-cigar smoker (finding)
C0425314|former cigar smoker (history)
C0425314|former cigar smoker
C0425314|Ex-cigar smoker (life style)
C0459838|Ex-cigarette smoker
C0459838|Ex-cigarette smoker (finding)
C0459838|Ex-cigarette smoker (life style)
C0425313|Ex-pipe smoker
C0425313|Ex-pipe smoker (finding)
C0425313|former pipe smoker
C0425313|former pipe smoker (history)
C0425313|Ex-pipe smoker (life style)
C1261257|Intolerant ex-smoker
C1261257|Intolerant ex-smoker (finding)
C1261257|Intolerant ex-smoker (life style)
C0425310|Stopped smoking
C0425310|Stopped smoking (finding)
C0425310|Stopped smoking (life style)
C0521322|Tolerant ex-smoker
C0521322|Tolerant ex-smoker (finding)
C0521322|Tolerant ex-smoker (life style)
C0558928|Ex-light smoker (1-9/day) (finding)
C0558928|Ex-light smoker (1-9/day)
C0558928|Ex-light smoker (1-9/day) (life style)
C0558927|Ex-trivial smoker (<1/day)
C0558927|Ex-trivial smoker (<1/day) (finding)
C0558927|Ex-trivial smoker (<1/day) (life style)
C0558929|Ex-moderate smoker (10-19/day)
C0558929|Ex-moderate smoker (10-19/day) (finding)
C0558929|Ex-moderate smoker (10-19/day) (life style)
C0558930|Ex-heavy smoker (20-39/day)
C0558930|Ex-heavy smoker (20-39/day) (finding)
C0558930|Ex-heavy smoker (20-39/day) (life style)
C0558931|Ex-very heavy smoker (40+/day) (finding)
C0558931|Ex-very heavy smoker (40+/day)
C0558931|Ex-very heavy smoker (40+/day) (life style)
C0558932|Ex-smoker - amount unknown
C0558932|Ex-smoker - amount unknown (finding)
C0558932|Ex-smoker - amount unknown (life style)
C3469008|never a smoker - tolerant
C3469008|never a smoker - tolerant (history)
C3469007|never a smoker - intolerant
C3469007|never a smoker - intolerant (history)
C3469006|never a smoker - aggressive (history)
C3469006|never a smoker - aggressive
C3472670|Never smoked any substance
C3472670|Never smoked any substance (finding)
C0425293|Never Smoked
C0425293|Never Smoker
C0425293|never smoked (history)
C0425293|Non-Smoker
C0425293|Never smoked tobacco
C0425293|Never smoked tobacco (finding)
C0425293|Never smoked tobacco (life style)
C3241966|Current Smoker
C3241966|current smoker (history)
C0337664|Smoker
C0337664|Smoker, NOS
C0337664|Smoker (finding)
C0337664|Smoker (life style)
C3494625|Current heavy tobacco smoker
C3494625|Heavy tobacco smoker (finding)
C3494625|Heavy tobacco smoker
C3494625|current heavy tobacco smoker (history)
C1883049|Smoker, Current Status Unknown
C1883049|smoker, current status unknown (history)
C3694955|current smoker duration (___ years) (history)
C3694955|current smoker duration (___ years)
C0459847|Heavy cigarette smoker
C0459847|Heavy cigarette smoker (finding)
C0459847|Heavy cigarette smoker (life style)
C0337666|Cigar smoker
C0337666|Smoking, Cigar
C0337666|Cigar smoking
C0337666|Cigar smoker (finding)
C0337666|Cigar smoker (life style)
C0337667|smoking cigarettes
C0337667|cigarette smoker
C0337667|smoking cigarettes (history)
C0337667|smokes cigarettes
C0337667|Cigarette smoker (finding)
C0337667|Cigarette smoker, NOS
C0337667|Cigarette smoker (life style)
C0337669|Heavy smoker (over 20 per day)
C0337669|Heavy smoker (over 20 per day) (finding)
C0337669|Heavy smoker (over 20 per day) (life style)
C0337668|current moderate tobacco smoker (history)
C0337668|current moderate tobacco smoker
C0337668|Moderate smoker (20 or less per day)
C0337668|Moderate smoker (20 or less per day) (finding)
C0337668|Moderate smoker (20 or less per day) (life style)
C0337665|Pipe smoker
C0337665|Pipe smoker (finding)
C0337665|Pipe smoker (life style)
C0425315|Smoking started - finding
C0425315|Smoking started
C0425315|Smoking started (finding)
C0425315|Smoking started (life style)
C3266136|Daily Smoker
C3266136|Current Every Day Smoker
C3266136|Every Day Smoker
C3266136|current every day smoker (history)
C3266136|Smokes tobacco daily
C3266136|Smokes tobacco daily (finding)
C3266136|Daily tobacco smoker
C3266136|Every-day smoker
C1883465|Unknown If Ever Smoked
C1883465|unknown if ever smoked (history)
