C0012634|T047|Diseases|
C0012634|T047|Disease|
C0012634|T047|DIS|
C0012634|T047|Disease or Disorder|
C0012634|T047|Diseases and Disorders|
C0012634|T047|diagnoses, syndromes, and conditions (diagnosis)|
C0012634|T047|diagnoses, syndromes, and conditions|
C0012634|T047|Disease [Disease/Finding]|
C0012634|T047|disease/disorder|
C0012634|T047|condition|
C0012634|T047|disorder|
C0012634|T047|Disorders|
C0012634|T047|Clinical disease AND/OR syndrome present|
C0012634|T047|Clinical disease AND/OR syndrome|
C0012634|T047|Disease (disorder)|
C0012634|T047|Disease AND/OR syndrome present|
C0012634|T047|disease (or disorder)|
C0012634|T047|Clinical disease or syndrome present, NOS|
C0012634|T047|Clinical disease or syndrome, NOS|
C0012634|T047|Disease or syndrome present, NOS|
C0012634|T047|Disease, NOS|
C0012634|T047|Disorder, NOS|
C1627937|T033|Medications on admission|
C1968515|T074|Pack (physical object)|
C1968515|T074|Pack|
C3840745|T033|Hospital emergency department|
C0225326|T121|Fiber|
C0225326|T121|Fiber, NOS|
C0225326|T121|Fiber -RETIRED-|
C0225326|T121|Fibre -RETIRED-|
C0225326|T121|Fibra|
C0225326|T121|Fibre|
C0225326|T121|Fiber (substance)|
C0225326|T121|Fiber (product)|
C1546956|T033|patient expired|
C1546956|T033|patient expired (diagnosis)|
C1546956|T033|overall condition: expired|
C1546956|T033|Dead|
C1546956|T033|Died|
C1546956|T033|Patient Outcome - Died|
C1546956|T033|Has died|
C1546956|T033|Dead (finding)|
C0275723|T047|Ovine interdigital dermatitis|
C0275723|T047|Foot scald|
C0275723|T047|Ovine interdigital dermatitis (disorder)|
C0275723|T047|OID|
C1522704|T061|Exercise|
C1522704|T061|Exercise Pain Management|
C0239966|T033|Hospital patient|
C0239966|T033|Hospital patient (& [inpatient])|
C0239966|T033|Hospital patient (& [inpatient]) (finding)|
C0239966|T033|Hospital inpatient|
C0239966|T033|patient currently in hospital (treatment)|
C0239966|T033|patient currently in hospital|
C0239966|T033|Hospital patient (finding)|
C0425043|T033|Death of relative|
C0425043|T033|Relative dying (context-dependent category)|
C0425043|T033|Relative dying (situation)|
C0425043|T033|Death in family|
C0425043|T033|death in family (history)|
C0425043|T033|Death in family, NOS|
C0425043|T033|Deceased Family Member|
C0425043|T033|Loss (of);relative;death|
C0425043|T033|Loss (of);relative|
C0425043|T033|Family members deceased|
C0425043|T033|Relatives died|
C0425043|T033|Family bereavement (finding)|
C0425043|T033|Family bereavement|
C0425043|T033|Relatives dead|
C0425043|T033|Relatives deceased|
C0425043|T033|Relatives died (finding)|
C0425043|T033|Death of family member|
C0425043|T033|Family members dead|
C0425043|T033|Family members died|
C0425043|T033|Death of relative (event)|
C0425043|T033|Cagemate death|
C0425043|T033|Relative dying|
C0425043|T033|loss of relative from death|
C0425043|T033|loss of relative|
C0425043|T033|Relative died|
C0557086|T033|No family|
C0557086|T033|No relatives|
C0557086|T033|No relatives (finding)|
C0011900|T033|Diagnoses|
C0011900|T033|Diagnosis|
C0011900|T033|Dx|
C0011900|T033|DIAG|
C0011900|T033|Diagnostic|
C0011900|T033|Diagnosed|
C0011900|T033|Diagnosis (observable entity)|
C0011900|T033|{Diagnosis}|
C0007465|T033|Cause of Death|
C0007465|T033|Death Cause|
C0007465|T033|Death Causes|
C0007465|T033|Death diagnosis (contextual qualifier)|
C0007465|T033|COD|
C0007465|T033|Cause of death (observable entity)|
C0007465|T033|Death--Causes|
C0007465|T033|Death Diagnosis|
C0007465|T033|DEATHD|
C0007465|T033|Causes of Death|
C0007465|T033|Condition fatal-cause of death|
C0007465|T033|Major cause of death|
C0007465|T033|DD|
C0007465|T033|Death diagnosis (contextual qualifier) (qualifier value)|
C0007465|T033|Cause of death (finding)|
C0002638|T031|Amniotic Fluid|
C0002638|T031|Amniotic Fluids|
C0002638|T031|Fluid, Amniotic|
C0002638|T031|Fluids, Amniotic|
C0002638|T031|Amniotic fluid (substance)|
C0002638|T031|AF - Amniotic fluid|
C0002638|T031|Liquor|
C0002638|T031|Aqua Amnii|
C0002638|T031|Liquor Amnii|
C0002638|T031|Waters (Amniotic Fluid)|
C0026606|T056|Activities, Motor|
C0026606|T056|Activity, Motor|
C0026606|T056|Motor Activities|
C0026606|T056|Motor Activity|
C0026606|T056|Physical Activities|
C0026606|T056|Physical activity|
C0026606|T056|Activities, Locomotor|
C0026606|T056|Activity, Locomotor|
C0026606|T056|Locomotor Activities|
C0026606|T056|Engaged in physical activity|
C0026606|T056|rndx activity|
C0026606|T056|rndx activity (diagnosis)|
C0026606|T056|Physical activity (observable entity)|
C0026606|T056|Physical activity (qualifier value)|
C0026606|T056|Activities, Physical|
C0026606|T056|Activity, Physical|
C0026606|T056|Locomotor Activity|
C0026606|T056|Motor behavior|
C0026606|T056|Motor behaviour|
C0026606|T056|Physical behavior|
C0026606|T056|Physical behaviour|
C0026606|T056|Motor activity, NOS|
C0026606|T056|Motor behavior, NOS|
C0026606|T056|Physical behavior, NOS|
C0026606|T056|Engaged in physical activity, NOS|
C0026606|T056|Motor behavior (function)|
C0026606|T056|Motor behavior, function (observable entity)|
C0026606|T056|Motor behavior (observable entity)|
C2349001|T016|Study Participant|
C2349001|T016|Human Study Subject|
C2349001|T016|Subject|
C2349001|T016|Human Subject|
C0455458|T033|History of - medical history NOS (context-dependent category)|
C0455458|T033|past medical history|
C0455458|T033|PMH|
C0455458|T033|past medical history (history)|
C0455458|T033|Health History|
C0455458|T033|PH|
C0455458|T033|H/O: medical history NOS (situation)|
C0455458|T033|Past medical history (situation)|
C0455458|T033|H/O: medical history NOS|
C0455458|T033|Past medical history of (contextual qualifier) (context-dependent category)|
C0455458|T033|History of - medical history NOS|
C0455458|T033|History of - medical history NOS (situation)|
C0455458|T033|Past medical history of|
C0455458|T033|PMH - past medical history|
C0455458|T033|Past history of|
C0455458|T033|health Hx|
C0006826|T191|Cancer|
C0006826|T191|Cancers|
C0006826|T191|Malignant neoplasm without specification of site|
C0006826|T191|Malignant Neoplasms|
C0006826|T191|CA|
C0006826|T191|Malignant neoplastic disease|
C0006826|T191|malignant neoplasm|
C0006826|T191|unspecified malignant neoplasm|
C0006826|T191|malignant neoplasm (diagnosis)|
C0006826|T191|cancer, NOS|
C0006826|T191|unspecified malignant neoplasm (diagnosis)|
C0006826|T191|Cancer NOS|
C0006826|T191|Malignancy|
C0006826|T191|neoplasm/cancer|
C0006826|T191|CA - Cancer|
C0006826|T191|Malignant neoplasm of unspecified site NOS (disorder)|
C0006826|T191|Malignant neoplasm of unspecified site|
C0006826|T191|Malignant tumor|
C0006826|T191|Malignant neoplasm of unspecified site (disorder)|
C0006826|T191|Malignant tumour|
C0006826|T191|Ca - unspecified site NOS|
C0006826|T191|Ca - unspecified site|
C0006826|T191|[X]Malignant neoplasm without specification of site|
C0006826|T191|Malignant neoplasm NOS|
C0006826|T191|Ca - unspecified site NOS (disorder)|
C0006826|T191|(Neoplasms) or (cancers) (disorder)|
C0006826|T191|Neoplasms - malignant|
C0006826|T191|[X]Malignant neoplasm without specification of site (disorder)|
C0006826|T191|Malignant tumour (disorder)|
C0006826|T191|(Neoplasms) or (cancers)|
C0006826|T191|Malignant neoplasm of unspecified site NOS|
C0006826|T191|NEOPLASM, MALIGNANT|
C0006826|T191|Malignant Growth|
C0006826|T191|Neoplasm malignant|
C0006826|T191|Cancer (NOS)|
C0006826|T191|Med: Malignant neoplastic disease|
C0006826|T191|Malignant neoplastic disease (disorder)|
C0006826|T191|tumor; malignant, unclassified|
C0006826|T191|tumor; unclassified, malignant|
C0006826|T191|Malignant tumor (disorder)|
C0006826|T191|Cancer, unspecified site|
C0006826|T191|Malignancy, unspecified site|
C0039082|T047|Syndromes|
C0039082|T047|Syndrome|
C0039082|T047|Syndrome [Disease/Finding]|
C0039082|T047|Clusters, Symptom|
C0039082|T047|Symptom Clusters|
C0039082|T047|Cluster, Symptom|
C0039082|T047|Symptom Cluster|
C0039082|T047|Syndrome, NOS|
C1509143|T033|H&P.PX|
C1509143|T033|Physical|
C1509143|T033|Physical assessment findings|
C1305866|T060|Weight|
C1305866|T060|Weighing Patient|
C1305866|T060|Weighing|
C1305866|T060|Weighing patient (procedure)|
C0080103|T099|Relation|
C0080103|T099|Relative (related person)|
C0080103|T099|Relative|
C0080103|T099|Relative (person)|
C0080103|T099|Relatives|
C0040336|T033|TOBACCO ABUSE|
C0040336|T033|Disorder, Tobacco Use|
C0040336|T033|Disorder, Tobacco-Use|
C0040336|T033|Tobacco Use Disorder|
C0040336|T033|Tobacco Use Disorders|
C0040336|T033|TOBACCO USE DIS|
C0040336|T033|Tobacco-Use Disorder|
C0040336|T033|Tobacco Use Disorder [Disease/Finding]|
C0040336|T033|rndx tobacco abuse|
C0040336|T033|rndx tobacco abuse (diagnosis)|
C0040336|T033|Abuse;tobacco|
C0040336|T033|tobacco abuse (diagnosis)|
C0040336|T033|abuse; tobacco|
C0040336|T033|tobacco; abuse|
C1514241|T033|Positive|
C1514241|T033|Positive Finding|
C0007457|T098|Caucasoid Race|
C0007457|T098|white race|
C0007457|T098|racial background Caucasian|
C0007457|T098|racial background Caucasian (history)|
C0007457|T098|Race: Caucasian|
C0007457|T098|Caucasian race|
C0007457|T098|Race: Caucasian (racial group)|
C0007457|T098|Race: Caucasian (finding)|
C0007457|T098|Race: White|
C0007457|T098|Caucasoid|
C0007457|T098|WHITE|
C0007457|T098|Caucasian Races|
C0007457|T098|Caucasoid Races|
C0007457|T098|Race, Caucasian|
C0007457|T098|Race, Caucasoid|
C0007457|T098|Races, Caucasian|
C0007457|T098|Races, Caucasoid|
C0007457|T098|Caucasian|
C0007457|T098|Whites|
C0007457|T098|Caucasians|
C0007457|T098|Occidental|
C0007457|T098|Caucasian (racial group)|
C0043157|T098|Caucasians|
C0043157|T098|caucasian|
C0043157|T098|RaceWhite|
C0043157|T098|Caucasian (living organism) (ethnic group)|
C0043157|T098|White - ethnic group (ethnic group)|
C0043157|T098|White - ethnic group|
C0043157|T098|White|
C0043157|T098|White/Caucasian|
C0043157|T098|Whites|
C0043157|T098|Caucasoid|
C0043157|T098|Caucasian (ethnic group)|
C0043157|T098|Caucasian, NOS|
C0043157|T098|Caucasian (living organism)|
C1261327|T033|Family history: Asthma (context-dependent category)|
C1261327|T033|Family history: Asthma (situation)|
C1261327|T033|Family history: Asthma|
C1261327|T033|FH: Asthma (situation)|
C1261327|T033|FH: Asthma|
C1261327|T033|Family history of asthma|
C1261327|T033|family history; asthma|
C1261327|T033|history; family, with asthma|
C0869014|T054|Relations|
C0262926|T033|Medical History|
C0262926|T033|Personal History|
C0262926|T033|History of (contextual qualifier)|
C0262926|T033|History|
C0262926|T033|Hx|
C0262926|T033|H&P.HX|
C0262926|T033|Past Medical History|
C0262926|T033|PMH|
C0262926|T033|personal medical history|
C0262926|T033|personal health record|
C0262926|T033|History of|
C0262926|T033|History of (contextual qualifier) (qualifier value)|
C0035253|T056|Rest|
C0035253|T056|Rests|
C0035253|T056|resting|
C0035253|T056|Rest (observable entity)|
C0035253|T056|Rest (qualifier value)|
C0489531|T033|History of allergies|
C0489531|T033|allergy (history)|
C0489531|T033|allergy|
C0489531|T033|allergies|
C0489531|T033|History of allergy|
C0424909|T033|Family history: Father (context-dependent category)|
C0424909|T033|Family history: Father NOS (context-dependent category)|
C0424909|T033|Family history: Father|
C0424909|T033|Family history with explicit context pertaining to father (situation)|
C0424909|T033|FH: Father|
C0424909|T033|Family history with explicit context pertaining to father|
C0424909|T033|Family history: Father (situation)|
C0424909|T033|FH: Father (situation)|
C0424909|T033|FH: Father NOS|
C0424909|T033|Family history: Father NOS (situation)|
C0424909|T033|Family history: Father NOS|
C0424909|T033|FH: Father NOS (situation)|
C0424909|T033|Paternal history|
C0042196|T061|Vaccination|
C0042196|T061|Vaccinations|
C0042196|T061|vaccinations (medication)|
C0042196|T061|vaccinations [use for free text]|
C0042196|T061|VACCIN|
C0042196|T061|Vaccine|
C0042196|T061|Inoculations - prophylactic|
C0042196|T061|Prophylactic vaccination|
C0042196|T061|Inoculation|
C0042196|T061|Vaccination, NOS|
C0042196|T061|Inoculation, NOS|
C0042196|T061|Vaccination NOS|
C0337671|T033|Former smoker|
C0337671|T033|Prior Smoker|
C0337671|T033|Past tobacco smoker|
C0337671|T033|Ex-smoker|
C0337671|T033|Ex-smoker (finding)|
C0337671|T033|Previous Tobacco Use|
C0337671|T033|Recovered smoker|
C0337671|T033|Cessation of smoking|
C0337671|T033|Ex-smoker (life style)|
C3668988|T033|Alert status|
C0301611|T168|Liquor|
C0301611|T168|distilled alcoholic beverage|
C0301611|T168|Distilled spirits|
C0301611|T168|Alcoholic spirits|
C0301611|T168|Spirits|
C0301611|T168|Distilled spirits (substance)|
C0559546|T046|Adverse Reaction|
C0559546|T046|ADR|
C0559546|T046|AR|
C0559546|T046|Adverse reactions|
C0559546|T046|Adverse reactions (disorder)|
C0559546|T046|Adverse reaction (disorder)|
C0559546|T046|adverse effect|
C0559546|T046|Adverse reactions (finding)|
C1527075|T061|Revision|
C1527075|T061|Revised|
C1527075|T061|Revise|
C1527075|T061|revision procedure (treatment)|
C1527075|T061|revision procedure|
C1527075|T061|Revision procedure (qualifier value)|
C0032854|T102|Poverty|
C0032854|T102|Poverty status|
C0032854|T102|Low Income|
C0032854|T102|Poor|
C0032854|T102|Financially poor|
C0032854|T102|Financially poor (finding)|
C0032854|T102|Social problem - poverty|
C0032854|T102|Economic deprivation|
C0032854|T102|Pauper|
C0032854|T102|Severe lack of money|
C0032854|T102|Living in poverty|
C0037125|T196|Silver|
C0037125|T196|Ag|
C0037125|T196|Silver [Chemical/Ingredient]|
C0037125|T196|Ag element|
C0037125|T196|Ag - Silver|
C0037125|T196|Silver (substance)|
C0037125|T196|Silver, NOS|
C3841837|T033|Hospitalization 3|
C1628992|T033|Admission diagnosis|

# C0015259|T056|Exercise| # JIRA/BIOMED-379
# C0015259|T056|Exercises|
# C0015259|T056|Exercises, Physical|
# C0015259|T056|Physical Exercise|
# C0015259|T056|Physical Exercises|
# C0015259|T056|Physical exercise NOS (procedure)|
# C0015259|T056|Physical exercises (procedure)|
# C0015259|T056|Physical exercise NOS (regime/therapy)|
# C0015259|T056|Physical exercise NOS|
# C0015259|T056|Exercise Type|
# C0015259|T056|Exercise, Physical|
# C0015259|T056|Physical exercises (regime/therapy)|
# C0015259|T056|Physical exercise, NOS|
# C0015259|T056|Exercise (observable entity)|
# C0015259|T056|Physical exercise (observable entity)|
# C0015259|T056|Exercise (qualifier value)|
# C0015259|T056|Physical exercise (qualifier value)|

C0241889|T033|Family history of (contextual qualifier) (context-dependent category)|
C0241889|T033|Family history: NOS (context-dependent category)|
C0241889|T033|family history|
C0241889|T033|family history (history)|
C0241889|T033|free text for family history (history)|
C0241889|T033|free text for family history|
C0241889|T033|family history free text|
C0241889|T033|Family history with explicit context|
C0241889|T033|Family history with explicit context (situation)|
C0241889|T033|Family history of (contextual qualifier) (situation)|
C0241889|T033|Family history of|
C0241889|T033|Family history of (contextual qualifier)|
C0241889|T033|Family health history (context-dependent category)|
C0241889|T033|Family history (situation)|
C0241889|T033|FH: NOS|
C0241889|T033|Family history: NOS|
C0241889|T033|Family history: NOS (situation)|
C0241889|T033|Family health history|
C0241889|T033|FH: NOS (situation)|
C0241889|T033|Family Medical History|
C0241889|T033|FH|
C0241889|T033|FH - Family history|
C0241889|T033|Family health history (finding)|
C0241889|T033|Epidemiology, Family Medical History|
C0204658|T060|Measuring height of patient|
C0204658|T060|Measuring height of patient (procedure)|
C0332123|T033|No family history: NOS (context-dependent category)|
C0332123|T033|No relevant family history (context-dependent category)|
C0332123|T033|No family history of (contextual qualifier)|
C0332123|T033|No family history of clinical finding (situation)|
C0332123|T033|No family history of clinical finding|
C0332123|T033|No relevant family history (situation)|
C0332123|T033|No family history|
C0332123|T033|No FH: NOS|
C0332123|T033|No FH: NOS (situation)|
C0332123|T033|No family history: NOS (situation)|
C0332123|T033|No family history: NOS|
C0332123|T033|NFH|
C0332123|T033|No family history of|
C0332123|T033|No relevant FH: family history|
C0332123|T033|No significant family history|
C0332123|T033|No family history of (contextual qualifier) (qualifier value)|
C0332123|T033|No relevant family history|
C0442735|T033|Nothing|
C0442735|T033|Nothing (qualifier value)|
C1519384|T033|Smoking History|
C1519384|T033|History of smoking (situation)|
C1519384|T033|History of smoking|
C0421451|T033|Patient date of birth|
C0421451|T033|BD|
C0421451|T033|DOB|
C0421451|T033|Date of Birth|
C0421451|T033|Birth Date|
C0421451|T033|Date of birth (finding)|
C0421451|T033|BRTHDAT|
C0421451|T033|birthDate|
C0421451|T033|DOB - Date of birth|
C0421451|T033|Date of birth (observable entity)|
C0421451|T033|Date of birth of person cared for|
C0421451|T033|Date of birth of recipient of care (observable entity)|
C0421451|T033|Date of birth of recipient of care|