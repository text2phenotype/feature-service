Procedure|surgery||ectomy|hysterectomy|removal, excision, resection
Procedure|surgery||tomy|orchidotomy|incision, cutting
Procedure|surgery||tome|osteotome|instrument to cut
Procedure|surgery||rrhaphy|herniorrhaphy|suture, repair
Procedure|surgery||plasty|rhytidoplasty|surgical repair
Procedure|surgery||desis|arthrodesis|binding
Procedure|surgery||clasis|osteoclasis|intentional breaking
Procedure|surgery||centesis|arthrocentisis|surgical puncture
Procedure|surgery||lithotomy|choledocholithotomy|incision for removal of a stone
Procedure|surgery||pexy|nephropexy|fixation, suspension
Procedure|surgery||stomy|gastrostomy|new opening
Procedure|surgery||pheresis|plasmapheresis|removal
Procedure|device|echo||echocardiography|sound, reverberation
Procedure|device||gram|echocardiogram|record, recording
Procedure|device||graph|echocardiograph|instrument to record
Procedure|device||graphy|echocardiography|process of recording
Procedure|viewing||opsy|biopsy|process of viewing
Procedure|viewing||scopy|bronchoscopy|process of viewing
Procedure|viewing||scope|otoscope|instrument to view
Procedure|measure||meter|tympanometer|instrument to measure
Procedure|measure||metry|spirometry|process of measurement
Procedure|device||trite|lithotrite|instrument to crush
Procedure|treatment||fusion|infusion|process of pouring
Procedure|treatment||therapy|hydrotherapy|treatment
Procedure|treatment||tripsy|lithotripsy|process of crushing
