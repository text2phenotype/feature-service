C0201838|Albumin measurement
C0523464|Albumin renal clearance measurement
C0523464|Albumin renal clearance measurement (procedure)
C0201837|Albumin/Globulin ratio
C0201837|Albumin globulin ratio
C0201837|A/G ratio
C0201837|Albumin/Globulin ratio (procedure)
C0523465|Serum albumin
C0523465|Serum Albumin Measurement
C0523465|ALBUMIN SERUM PLASMA/WHOLE BLOOD
C0523465|Albumin; serum, plasma or whole blood
C0523465|serum albumin measurement (lab test)
C0523465|Measurement of albumin in serum
C0523465|Serum albumin (& level) (procedure)
C0523465|Albumin - serum
C0523465|Serum albumin (& level)
C0523465|Serum Albumin Test
C0523465|Albumin measurement, serum
C0523465|Serum albumin level
C0523465|SA - Serum albumin
C0523465|Albumin measurement, serum (procedure)
C0523465|ASSAY OF SERUM ALBUMIN
C0201838|Albumin measurement
C0201838|Test;albumin
C0201838|Measurement of albumin
C0201838|Albumin
C0201838|ALB
C0201838|Microalbumin
C0201838|Albumin measurement (procedure)
C0201838|albumin test
C1278236|24 hour urine albumin output
C1278236|24 hour urine albumin output (procedure)
C1278236|24 hour urine albumin output measurement (procedure)
C1278236|24 hour urine albumin output measurement
C0523466|Albumin; urine or other source, quantitative, each specimen
C0523466|ALBUMIN URINE/OTHER SOURCE QUAN EACH SPECIMEN
C0523466|Albumin measurement, urine, quantitative
C0523466|Albumin measurement, urine, quantitative (procedure)
C0523466|ASSAY OF URINE ALBUMIN
C0373533|Albumin; urine, microalbumin, semiquantitative (eg, reagent strip assay)
C0373533|MICROALBUMIN SEMIQUANT
C0373533|ALBUMIN URINE MICROALBUMIN SEMIQUANTITATIVE
C0373533|Semiquantitative analysis of microalbumin in urine
C1504155|serum albumin ischemia modified (lab test)
C1504155|serum albumin ischemia modified
C1504155|ischemia-modified serum albumin
C1504155|ALBUMIN ISCHEMIA MODIFIED
C1504155|serum albumin ischemia modified lab procedure
C1504155|Albumin; ischemia modified
C0373532|Albumin; urine, microalbumin, quantitative
C0373532|MICROALBUMIN QUANTITATIVE
C0373532|ALBUMIN URINE MICROALBUMIN QUANTIATIVE
C0523674|ALBGLYCA
C0523674|Glycated Albumin
C0523674|Glycated Albumin Measurement
C0523674|Glycated albumin measurement (procedure)
C1278275|Cerebrospinal fluid albumin level
C1278275|Cerebrospinal fluid albumin level (procedure)
C1278275|Cerebrospinal fluid albumin measurement (procedure)
C1278275|Cerebrospinal fluid albumin measurement
C0428520|Fluid sample albumin level
C0428520|Fluid sample albumin measurement (procedure)
C0428520|Fluid sample albumin measurement
C0428623|Albumin/immunoglobulin G ratio
C0428623|IgG - Albumin/immunoglobulin G ratio
C0428623|Albumin/immunoglobulin G ratio measurement (procedure)
C0428623|Albumin/immunoglobulin G ratio measurement
C1272106|Plasma albumin level (procedure)
C1272106|Plasma albumin level
C1273508|Serum prealbumin level
C1273508|Serum prealbumin level (procedure)
C1318429|Measurement of albumin in urine
C1318429|Urine albumin (& level) (procedure)
C1318429|Urine albumin (& level)
C1318429|Urine albumin level
C1318429|Urine albumin measurement (procedure)
C1318429|Urine albumin measurement
C0523463|CSF albumin/plasma albumin ratio measurement (procedure)
C0523463|Cerebrospinal fluid albumin/plasma albumin ratio measurement (procedure)
C0523463|Cerebrospinal fluid albumin/plasma albumin ratio measurement
C0523463|CSF albumin/plasma albumin ratio measurement
C0025634|Methemalbumin
C0025634|Methemalbumin Assay
C0025634|Methemalbumin (protein) level
C0025634|Measurement of methemalbumin
C0025634|Methemalbumin measurement
C0025634|Methaemalbumin measurement
C0025634|Methemalbumin measurement (procedure)
C0025634|ASSAY OF METHEMALBUMIN
C1293929|Measurement of ratio of analyte to albumin (procedure)
C1293929|Measurement of ratio of analyte to albumin
